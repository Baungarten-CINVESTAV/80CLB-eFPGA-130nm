magic
tech sky130A
magscale 1 2
timestamp 1708041251
<< obsli1 >>
rect 1104 2159 10856 9809
<< obsm1 >>
rect 842 1640 11118 9840
<< metal2 >>
rect 846 0 902 800
rect 1766 0 1822 800
rect 2686 0 2742 800
rect 3606 0 3662 800
rect 4526 0 4582 800
rect 5446 0 5502 800
rect 6366 0 6422 800
rect 7286 0 7342 800
rect 8206 0 8262 800
rect 9126 0 9182 800
rect 10046 0 10102 800
<< obsm2 >>
rect 848 856 11114 11529
rect 958 31 1710 856
rect 1878 31 2630 856
rect 2798 31 3550 856
rect 3718 31 4470 856
rect 4638 31 5390 856
rect 5558 31 6310 856
rect 6478 31 7230 856
rect 7398 31 8150 856
rect 8318 31 9070 856
rect 9238 31 9990 856
rect 10158 31 11114 856
<< metal3 >>
rect 11200 11432 12000 11552
rect 0 11160 800 11280
rect 11200 10888 12000 11008
rect 11200 10344 12000 10464
rect 0 10072 800 10192
rect 11200 9800 12000 9920
rect 11200 9256 12000 9376
rect 0 8984 800 9104
rect 11200 8712 12000 8832
rect 11200 8168 12000 8288
rect 0 7896 800 8016
rect 11200 7624 12000 7744
rect 11200 7080 12000 7200
rect 0 6808 800 6928
rect 11200 6536 12000 6656
rect 11200 5992 12000 6112
rect 0 5720 800 5840
rect 11200 5448 12000 5568
rect 11200 4904 12000 5024
rect 0 4632 800 4752
rect 11200 4360 12000 4480
rect 11200 3816 12000 3936
rect 0 3544 800 3664
rect 11200 3272 12000 3392
rect 11200 2728 12000 2848
rect 0 2456 800 2576
rect 11200 2184 12000 2304
rect 11200 1640 12000 1760
rect 0 1368 800 1488
rect 11200 1096 12000 1216
rect 11200 552 12000 672
rect 11200 8 12000 128
<< obsm3 >>
rect 798 11360 11120 11525
rect 880 11352 11120 11360
rect 880 11088 11530 11352
rect 880 11080 11120 11088
rect 798 10808 11120 11080
rect 798 10544 11530 10808
rect 798 10272 11120 10544
rect 880 10264 11120 10272
rect 880 10000 11530 10264
rect 880 9992 11120 10000
rect 798 9720 11120 9992
rect 798 9456 11530 9720
rect 798 9184 11120 9456
rect 880 9176 11120 9184
rect 880 8912 11530 9176
rect 880 8904 11120 8912
rect 798 8632 11120 8904
rect 798 8368 11530 8632
rect 798 8096 11120 8368
rect 880 8088 11120 8096
rect 880 7824 11530 8088
rect 880 7816 11120 7824
rect 798 7544 11120 7816
rect 798 7280 11530 7544
rect 798 7008 11120 7280
rect 880 7000 11120 7008
rect 880 6736 11530 7000
rect 880 6728 11120 6736
rect 798 6456 11120 6728
rect 798 6192 11530 6456
rect 798 5920 11120 6192
rect 880 5912 11120 5920
rect 880 5648 11530 5912
rect 880 5640 11120 5648
rect 798 5368 11120 5640
rect 798 5104 11530 5368
rect 798 4832 11120 5104
rect 880 4824 11120 4832
rect 880 4560 11530 4824
rect 880 4552 11120 4560
rect 798 4280 11120 4552
rect 798 4016 11530 4280
rect 798 3744 11120 4016
rect 880 3736 11120 3744
rect 880 3472 11530 3736
rect 880 3464 11120 3472
rect 798 3192 11120 3464
rect 798 2928 11530 3192
rect 798 2656 11120 2928
rect 880 2648 11120 2656
rect 880 2384 11530 2648
rect 880 2376 11120 2384
rect 798 2104 11120 2376
rect 798 1840 11530 2104
rect 798 1568 11120 1840
rect 880 1560 11120 1568
rect 880 1296 11530 1560
rect 880 1288 11120 1296
rect 798 1016 11120 1288
rect 798 752 11530 1016
rect 798 472 11120 752
rect 798 208 11530 472
rect 798 35 11120 208
<< metal4 >>
rect 2163 2128 2483 9840
rect 3382 2128 3702 9840
rect 4601 2128 4921 9840
rect 5820 2128 6140 9840
rect 7039 2128 7359 9840
rect 8258 2128 8578 9840
rect 9477 2128 9797 9840
rect 10696 2128 11016 9840
<< labels >>
rlabel metal2 s 846 0 902 800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 2 nsew signal input
rlabel metal3 s 11200 5448 12000 5568 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 11200 5992 12000 6112 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 11200 552 12000 672 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 11200 1096 12000 1216 6 chanx_right_in[1]
port 6 nsew signal input
rlabel metal3 s 11200 1640 12000 1760 6 chanx_right_in[2]
port 7 nsew signal input
rlabel metal3 s 11200 2184 12000 2304 6 chanx_right_in[3]
port 8 nsew signal input
rlabel metal3 s 11200 2728 12000 2848 6 chanx_right_in[4]
port 9 nsew signal input
rlabel metal3 s 11200 3272 12000 3392 6 chanx_right_in[5]
port 10 nsew signal input
rlabel metal3 s 11200 3816 12000 3936 6 chanx_right_in[6]
port 11 nsew signal input
rlabel metal3 s 11200 4360 12000 4480 6 chanx_right_in[7]
port 12 nsew signal input
rlabel metal3 s 11200 4904 12000 5024 6 chanx_right_in[8]
port 13 nsew signal input
rlabel metal3 s 11200 7080 12000 7200 6 chanx_right_out[0]
port 14 nsew signal output
rlabel metal3 s 11200 7624 12000 7744 6 chanx_right_out[1]
port 15 nsew signal output
rlabel metal3 s 11200 8168 12000 8288 6 chanx_right_out[2]
port 16 nsew signal output
rlabel metal3 s 11200 8712 12000 8832 6 chanx_right_out[3]
port 17 nsew signal output
rlabel metal3 s 11200 9256 12000 9376 6 chanx_right_out[4]
port 18 nsew signal output
rlabel metal3 s 11200 9800 12000 9920 6 chanx_right_out[5]
port 19 nsew signal output
rlabel metal3 s 11200 10344 12000 10464 6 chanx_right_out[6]
port 20 nsew signal output
rlabel metal3 s 11200 10888 12000 11008 6 chanx_right_out[7]
port 21 nsew signal output
rlabel metal3 s 11200 11432 12000 11552 6 chanx_right_out[8]
port 22 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[0]
port 23 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_in[1]
port 24 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_in[2]
port 25 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[3]
port 26 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[4]
port 27 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[5]
port 28 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[6]
port 29 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_in[7]
port 30 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[8]
port 31 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 chany_bottom_out[0]
port 32 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 chany_bottom_out[1]
port 33 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 chany_bottom_out[2]
port 34 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 chany_bottom_out[3]
port 35 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 chany_bottom_out[4]
port 36 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 chany_bottom_out[5]
port 37 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 chany_bottom_out[6]
port 38 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 chany_bottom_out[7]
port 39 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 chany_bottom_out[8]
port 40 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 prog_clk
port 41 nsew signal input
rlabel metal3 s 11200 6536 12000 6656 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 42 nsew signal input
rlabel metal3 s 11200 8 12000 128 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 43 nsew signal input
rlabel metal4 s 2163 2128 2483 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 3382 2128 3702 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 5820 2128 6140 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 8258 2128 8578 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 10696 2128 11016 9840 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 364594
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_0__10_/runs/24_02_15_17_53/results/signoff/sb_0__10_.magic.gds
string GDS_START 89996
<< end >>

