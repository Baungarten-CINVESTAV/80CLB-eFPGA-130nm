magic
tech sky130A
magscale 1 2
timestamp 1707852921
<< viali >>
rect 4721 9673 4755 9707
rect 10241 9673 10275 9707
rect 1777 9605 1811 9639
rect 2145 9605 2179 9639
rect 2973 9605 3007 9639
rect 1501 9537 1535 9571
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3617 9537 3651 9571
rect 4353 9537 4387 9571
rect 4445 9537 4479 9571
rect 4905 9537 4939 9571
rect 6193 9537 6227 9571
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 7573 9537 7607 9571
rect 7849 9537 7883 9571
rect 8769 9537 8803 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 7941 9469 7975 9503
rect 7113 9401 7147 9435
rect 9597 9401 9631 9435
rect 1685 9333 1719 9367
rect 2605 9333 2639 9367
rect 3341 9333 3375 9367
rect 3433 9333 3467 9367
rect 4261 9333 4295 9367
rect 4537 9333 4571 9367
rect 4997 9333 5031 9367
rect 6009 9333 6043 9367
rect 6745 9333 6779 9367
rect 7481 9333 7515 9367
rect 7665 9333 7699 9367
rect 8585 9333 8619 9367
rect 1685 9129 1719 9163
rect 4353 9129 4387 9163
rect 5825 9129 5859 9163
rect 7481 9129 7515 9163
rect 8309 9129 8343 9163
rect 10425 9129 10459 9163
rect 3617 9061 3651 9095
rect 3801 9061 3835 9095
rect 7941 9061 7975 9095
rect 2237 8993 2271 9027
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 7757 8993 7791 9027
rect 1961 8925 1995 8959
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 4813 8925 4847 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 7573 8925 7607 8959
rect 8493 8925 8527 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 2513 8857 2547 8891
rect 6368 8857 6402 8891
rect 2697 8789 2731 8823
rect 2973 8789 3007 8823
rect 5457 8789 5491 8823
rect 9689 8789 9723 8823
rect 9965 8789 9999 8823
rect 3249 8585 3283 8619
rect 6377 8585 6411 8619
rect 7113 8585 7147 8619
rect 1777 8517 1811 8551
rect 4988 8517 5022 8551
rect 9260 8517 9294 8551
rect 2965 8449 2999 8483
rect 3065 8449 3099 8483
rect 4362 8449 4396 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 9781 8449 9815 8483
rect 10149 8449 10183 8483
rect 2145 8381 2179 8415
rect 2329 8381 2363 8415
rect 4629 8381 4663 8415
rect 4721 8381 4755 8415
rect 6929 8381 6963 8415
rect 9505 8381 9539 8415
rect 1501 8313 1535 8347
rect 6101 8313 6135 8347
rect 2697 8245 2731 8279
rect 8125 8245 8159 8279
rect 9689 8245 9723 8279
rect 10425 8245 10459 8279
rect 4445 8041 4479 8075
rect 4997 8041 5031 8075
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 3433 7973 3467 8007
rect 3801 7905 3835 7939
rect 6193 7905 6227 7939
rect 7573 7905 7607 7939
rect 9781 7905 9815 7939
rect 2053 7837 2087 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 6101 7837 6135 7871
rect 6377 7837 6411 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 7389 7837 7423 7871
rect 8585 7837 8619 7871
rect 9597 7837 9631 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 1409 7769 1443 7803
rect 1777 7769 1811 7803
rect 2298 7769 2332 7803
rect 6561 7701 6595 7735
rect 8769 7701 8803 7735
rect 9137 7701 9171 7735
rect 10057 7701 10091 7735
rect 10425 7701 10459 7735
rect 2053 7497 2087 7531
rect 3525 7497 3559 7531
rect 4629 7497 4663 7531
rect 5089 7497 5123 7531
rect 5457 7497 5491 7531
rect 9045 7497 9079 7531
rect 9229 7497 9263 7531
rect 1501 7361 1535 7395
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 3893 7361 3927 7395
rect 5181 7361 5215 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6653 7361 6687 7395
rect 8585 7361 8619 7395
rect 8861 7361 8895 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 2605 7293 2639 7327
rect 2789 7293 2823 7327
rect 3985 7293 4019 7327
rect 4169 7293 4203 7327
rect 4721 7293 4755 7327
rect 6101 7293 6135 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 8309 7293 8343 7327
rect 9689 7293 9723 7327
rect 9873 7293 9907 7327
rect 10057 7293 10091 7327
rect 2973 7225 3007 7259
rect 3341 7225 3375 7259
rect 3709 7225 3743 7259
rect 6561 7225 6595 7259
rect 6837 7225 6871 7259
rect 8401 7225 8435 7259
rect 10333 7225 10367 7259
rect 2421 7157 2455 7191
rect 5825 7157 5859 7191
rect 7573 7157 7607 7191
rect 7665 7157 7699 7191
rect 1409 6953 1443 6987
rect 7757 6953 7791 6987
rect 10057 6953 10091 6987
rect 10425 6953 10459 6987
rect 5089 6885 5123 6919
rect 2789 6817 2823 6851
rect 4721 6817 4755 6851
rect 5457 6817 5491 6851
rect 9229 6817 9263 6851
rect 3525 6749 3559 6783
rect 3801 6749 3835 6783
rect 4537 6749 4571 6783
rect 5273 6749 5307 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 8585 6749 8619 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9965 6749 9999 6783
rect 10241 6749 10275 6783
rect 2544 6681 2578 6715
rect 2973 6681 3007 6715
rect 4077 6681 4111 6715
rect 5549 6681 5583 6715
rect 3985 6613 4019 6647
rect 6837 6613 6871 6647
rect 8769 6613 8803 6647
rect 8953 6613 8987 6647
rect 9873 6613 9907 6647
rect 2145 6409 2179 6443
rect 5549 6409 5583 6443
rect 7205 6409 7239 6443
rect 8953 6409 8987 6443
rect 9873 6409 9907 6443
rect 6377 6341 6411 6375
rect 1409 6273 1443 6307
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 3433 6273 3467 6307
rect 4741 6273 4775 6307
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 6193 6273 6227 6307
rect 7113 6273 7147 6307
rect 7573 6273 7607 6307
rect 7849 6273 7883 6307
rect 8769 6273 8803 6307
rect 8861 6273 8895 6307
rect 9229 6273 9263 6307
rect 9965 6273 9999 6307
rect 10241 6273 10275 6307
rect 3249 6205 3283 6239
rect 6009 6205 6043 6239
rect 6837 6205 6871 6239
rect 7021 6205 7055 6239
rect 8033 6205 8067 6239
rect 9413 6205 9447 6239
rect 7757 6137 7791 6171
rect 8585 6137 8619 6171
rect 2329 6069 2363 6103
rect 2697 6069 2731 6103
rect 3065 6069 3099 6103
rect 3617 6069 3651 6103
rect 5457 6069 5491 6103
rect 8493 6069 8527 6103
rect 10425 6069 10459 6103
rect 2145 5865 2179 5899
rect 3617 5865 3651 5899
rect 4905 5865 4939 5899
rect 5917 5865 5951 5899
rect 6837 5865 6871 5899
rect 7849 5865 7883 5899
rect 2513 5797 2547 5831
rect 4721 5797 4755 5831
rect 6101 5797 6135 5831
rect 2605 5729 2639 5763
rect 2789 5729 2823 5763
rect 9045 5729 9079 5763
rect 9689 5729 9723 5763
rect 10149 5729 10183 5763
rect 1961 5661 1995 5695
rect 2329 5661 2363 5695
rect 3433 5661 3467 5695
rect 3985 5661 4019 5695
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 5825 5661 5859 5695
rect 6285 5661 6319 5695
rect 6929 5661 6963 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 8217 5661 8251 5695
rect 1501 5593 1535 5627
rect 8401 5593 8435 5627
rect 9137 5593 9171 5627
rect 9873 5593 9907 5627
rect 9965 5593 9999 5627
rect 1593 5525 1627 5559
rect 3249 5525 3283 5559
rect 3801 5525 3835 5559
rect 7573 5525 7607 5559
rect 8125 5525 8159 5559
rect 8677 5525 8711 5559
rect 2513 5321 2547 5355
rect 4353 5253 4387 5287
rect 5365 5253 5399 5287
rect 7849 5253 7883 5287
rect 1777 5185 1811 5219
rect 2237 5185 2271 5219
rect 2329 5185 2363 5219
rect 4629 5185 4663 5219
rect 4905 5185 4939 5219
rect 6377 5185 6411 5219
rect 6644 5185 6678 5219
rect 9413 5185 9447 5219
rect 5273 5117 5307 5151
rect 6009 5117 6043 5151
rect 9689 5117 9723 5151
rect 4813 5049 4847 5083
rect 5089 5049 5123 5083
rect 5825 5049 5859 5083
rect 7757 5049 7791 5083
rect 1501 4981 1535 5015
rect 2145 4981 2179 5015
rect 3065 4981 3099 5015
rect 10333 4981 10367 5015
rect 1409 4777 1443 4811
rect 5917 4777 5951 4811
rect 8677 4777 8711 4811
rect 2605 4709 2639 4743
rect 4169 4709 4203 4743
rect 8953 4709 8987 4743
rect 2881 4641 2915 4675
rect 3341 4641 3375 4675
rect 4537 4641 4571 4675
rect 7481 4641 7515 4675
rect 7849 4641 7883 4675
rect 8033 4641 8067 4675
rect 8493 4641 8527 4675
rect 1593 4573 1627 4607
rect 1685 4573 1719 4607
rect 1961 4573 1995 4607
rect 2145 4573 2179 4607
rect 2697 4573 2731 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 6101 4573 6135 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7021 4573 7055 4607
rect 7757 4573 7791 4607
rect 8585 4573 8619 4607
rect 10066 4573 10100 4607
rect 10333 4573 10367 4607
rect 1777 4505 1811 4539
rect 4804 4505 4838 4539
rect 3617 4437 3651 4471
rect 7665 4437 7699 4471
rect 1961 4233 1995 4267
rect 5181 4233 5215 4267
rect 6745 4233 6779 4267
rect 7021 4233 7055 4267
rect 7757 4233 7791 4267
rect 8033 4233 8067 4267
rect 8769 4233 8803 4267
rect 5457 4165 5491 4199
rect 1777 4097 1811 4131
rect 2145 4097 2179 4131
rect 2605 4097 2639 4131
rect 2697 4097 2731 4131
rect 3617 4097 3651 4131
rect 3801 4097 3835 4131
rect 4068 4097 4102 4131
rect 6561 4097 6595 4131
rect 6837 4097 6871 4131
rect 7297 4097 7331 4131
rect 7849 4097 7883 4131
rect 8677 4097 8711 4131
rect 10066 4097 10100 4131
rect 10333 4097 10367 4131
rect 2881 4029 2915 4063
rect 5365 4029 5399 4063
rect 7113 4029 7147 4063
rect 3433 3961 3467 3995
rect 5917 3961 5951 3995
rect 8953 3961 8987 3995
rect 1501 3893 1535 3927
rect 2513 3893 2547 3927
rect 3341 3893 3375 3927
rect 2421 3689 2455 3723
rect 3341 3689 3375 3723
rect 4997 3689 5031 3723
rect 7205 3689 7239 3723
rect 9689 3689 9723 3723
rect 10517 3689 10551 3723
rect 4813 3621 4847 3655
rect 5917 3621 5951 3655
rect 2881 3553 2915 3587
rect 2145 3485 2179 3519
rect 2605 3485 2639 3519
rect 2697 3485 2731 3519
rect 3801 3485 3835 3519
rect 4721 3485 4755 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 7297 3485 7331 3519
rect 9229 3485 9263 3519
rect 9505 3485 9539 3519
rect 9873 3485 9907 3519
rect 1409 3417 1443 3451
rect 1777 3417 1811 3451
rect 2237 3349 2271 3383
rect 3893 3349 3927 3383
rect 9413 3349 9447 3383
rect 1593 3145 1627 3179
rect 2237 3145 2271 3179
rect 3433 3145 3467 3179
rect 3709 3145 3743 3179
rect 3801 3145 3835 3179
rect 8953 3145 8987 3179
rect 9689 3145 9723 3179
rect 9413 3077 9447 3111
rect 1409 3009 1443 3043
rect 1777 3009 1811 3043
rect 2053 3009 2087 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 3525 3009 3559 3043
rect 3985 3009 4019 3043
rect 8769 3009 8803 3043
rect 9045 3009 9079 3043
rect 9965 3009 9999 3043
rect 1869 2805 1903 2839
rect 2697 2805 2731 2839
rect 9229 2805 9263 2839
rect 10241 2805 10275 2839
rect 2697 2601 2731 2635
rect 5641 2601 5675 2635
rect 6837 2601 6871 2635
rect 7849 2601 7883 2635
rect 8769 2601 8803 2635
rect 9505 2601 9539 2635
rect 3249 2533 3283 2567
rect 3985 2533 4019 2567
rect 4445 2533 4479 2567
rect 1777 2397 1811 2431
rect 2237 2397 2271 2431
rect 2513 2397 2547 2431
rect 2973 2397 3007 2431
rect 3065 2397 3099 2431
rect 3341 2397 3375 2431
rect 3801 2397 3835 2431
rect 4261 2397 4295 2431
rect 5457 2397 5491 2431
rect 6653 2397 6687 2431
rect 8033 2397 8067 2431
rect 8585 2397 8619 2431
rect 9045 2397 9079 2431
rect 9321 2397 9355 2431
rect 9689 2397 9723 2431
rect 1409 2329 1443 2363
rect 3433 2329 3467 2363
rect 10149 2329 10183 2363
rect 2145 2261 2179 2295
rect 2789 2261 2823 2295
rect 9229 2261 9263 2295
rect 9873 2261 9907 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 3712 9676 4721 9704
rect 934 9596 940 9648
rect 992 9636 998 9648
rect 1765 9639 1823 9645
rect 1765 9636 1777 9639
rect 992 9608 1777 9636
rect 992 9596 998 9608
rect 1765 9605 1777 9608
rect 1811 9605 1823 9639
rect 1765 9599 1823 9605
rect 2038 9596 2044 9648
rect 2096 9596 2102 9648
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9636 2191 9639
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2179 9608 2973 9636
rect 2179 9605 2191 9608
rect 2133 9599 2191 9605
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 2961 9599 3019 9605
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 2056 9568 2084 9596
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 1535 9540 2084 9568
rect 2608 9540 2697 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 2608 9432 2636 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3252 9568 3280 9596
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3252 9540 3617 9568
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3712 9500 3740 9676
rect 4709 9673 4721 9676
rect 4755 9673 4767 9707
rect 4709 9667 4767 9673
rect 6178 9664 6184 9716
rect 6236 9664 6242 9716
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 8662 9664 8668 9716
rect 8720 9664 8726 9716
rect 9766 9664 9772 9716
rect 9824 9664 9830 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10318 9704 10324 9716
rect 10275 9676 10324 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 3896 9608 4476 9636
rect 3896 9512 3924 9608
rect 4338 9528 4344 9580
rect 4396 9528 4402 9580
rect 4448 9577 4476 9608
rect 4614 9596 4620 9648
rect 4672 9636 4678 9648
rect 4672 9608 4936 9636
rect 4672 9596 4678 9608
rect 4908 9577 4936 9608
rect 6196 9577 6224 9664
rect 7208 9636 7236 9664
rect 6932 9608 7236 9636
rect 6932 9577 6960 9608
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7374 9568 7380 9580
rect 7239 9540 7380 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 7742 9568 7748 9580
rect 7607 9540 7748 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 7834 9528 7840 9580
rect 7892 9528 7898 9580
rect 8680 9568 8708 9664
rect 9784 9577 9812 9664
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8680 9540 8769 9568
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9950 9528 9956 9580
rect 10008 9528 10014 9580
rect 3016 9472 3740 9500
rect 3016 9460 3022 9472
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 4126 9472 4844 9500
rect 4126 9432 4154 9472
rect 2608 9404 4154 9432
rect 4816 9432 4844 9472
rect 5442 9460 5448 9512
rect 5500 9460 5506 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5675 9472 5733 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 5721 9469 5733 9472
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 5960 9472 7880 9500
rect 5960 9460 5966 9472
rect 7101 9435 7159 9441
rect 7101 9432 7113 9435
rect 4816 9404 7113 9432
rect 7101 9401 7113 9404
rect 7147 9401 7159 9435
rect 7852 9432 7880 9472
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 7852 9404 9597 9432
rect 7101 9395 7159 9401
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 1670 9324 1676 9376
rect 1728 9324 1734 9376
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 2774 9364 2780 9376
rect 2639 9336 2780 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3326 9324 3332 9376
rect 3384 9324 3390 9376
rect 3418 9324 3424 9376
rect 3476 9324 3482 9376
rect 4246 9324 4252 9376
rect 4304 9324 4310 9376
rect 4522 9324 4528 9376
rect 4580 9324 4586 9376
rect 4982 9324 4988 9376
rect 5040 9324 5046 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 6178 9364 6184 9376
rect 6043 9336 6184 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6730 9324 6736 9376
rect 6788 9324 6794 9376
rect 7466 9324 7472 9376
rect 7524 9324 7530 9376
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8076 9336 8585 9364
rect 8076 9324 8082 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 1578 9120 1584 9172
rect 1636 9160 1642 9172
rect 1673 9163 1731 9169
rect 1673 9160 1685 9163
rect 1636 9132 1685 9160
rect 1636 9120 1642 9132
rect 1673 9129 1685 9132
rect 1719 9129 1731 9163
rect 1673 9123 1731 9129
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 3418 9160 3424 9172
rect 2556 9132 3424 9160
rect 2556 9120 2562 9132
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4246 9160 4252 9172
rect 3528 9132 4252 9160
rect 3528 9092 3556 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4982 9160 4988 9172
rect 4396 9132 4988 9160
rect 4396 9120 4402 9132
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5132 9132 5825 9160
rect 5132 9120 5138 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 6730 9160 6736 9172
rect 5813 9123 5871 9129
rect 6012 9132 6736 9160
rect 2746 9064 3556 9092
rect 3605 9095 3663 9101
rect 1118 8984 1124 9036
rect 1176 9024 1182 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 1176 8996 2237 9024
rect 1176 8984 1182 8996
rect 2225 8993 2237 8996
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2746 8956 2774 9064
rect 3605 9061 3617 9095
rect 3651 9061 3663 9095
rect 3605 9055 3663 9061
rect 3789 9095 3847 9101
rect 3789 9061 3801 9095
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3620 9024 3648 9055
rect 3108 8996 3188 9024
rect 3108 8984 3114 8996
rect 3160 8965 3188 8996
rect 3344 8996 3648 9024
rect 1995 8928 2774 8956
rect 2869 8959 2927 8965
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 3145 8959 3203 8965
rect 2915 8928 3096 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 2547 8860 3004 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 2682 8780 2688 8832
rect 2740 8780 2746 8832
rect 2976 8829 3004 8860
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8789 3019 8823
rect 3068 8820 3096 8928
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3344 8888 3372 8996
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3804 8956 3832 9055
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 5902 9092 5908 9104
rect 4212 9064 5908 9092
rect 4212 9052 4218 9064
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 4522 8984 4528 9036
rect 4580 8984 4586 9036
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4982 9024 4988 9036
rect 4755 8996 4988 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 3467 8928 3832 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3936 8928 3985 8956
rect 3936 8916 3942 8928
rect 3973 8925 3985 8928
rect 4019 8956 4031 8959
rect 4801 8959 4859 8965
rect 4019 8928 4476 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4448 8888 4476 8928
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4816 8888 4844 8919
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 6012 8965 6040 9132
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7469 9163 7527 9169
rect 7469 9129 7481 9163
rect 7515 9160 7527 9163
rect 7742 9160 7748 9172
rect 7515 9132 7748 9160
rect 7515 9129 7527 9132
rect 7469 9123 7527 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 7892 9132 8309 9160
rect 7892 9120 7898 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 9950 9120 9956 9172
rect 10008 9120 10014 9172
rect 10410 9120 10416 9172
rect 10468 9120 10474 9172
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7432 9064 7941 9092
rect 7432 9052 7438 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 7929 9055 7987 9061
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7524 8996 7757 9024
rect 7524 8984 7530 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 9968 9024 9996 9120
rect 11054 9052 11060 9104
rect 11112 9052 11118 9104
rect 11072 9024 11100 9052
rect 7892 8996 9996 9024
rect 10152 8996 11100 9024
rect 7892 8984 7898 8996
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6135 8928 6914 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 5460 8888 5488 8916
rect 6362 8897 6368 8900
rect 3344 8860 4384 8888
rect 4448 8860 4844 8888
rect 4908 8860 5488 8888
rect 4154 8820 4160 8832
rect 3068 8792 4160 8820
rect 2961 8783 3019 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4356 8820 4384 8860
rect 4908 8820 4936 8860
rect 6356 8851 6368 8897
rect 6362 8848 6368 8851
rect 6420 8848 6426 8900
rect 6886 8888 6914 8928
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 8496 8965 8524 8996
rect 10152 8965 10180 8996
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 9490 8888 9496 8900
rect 6886 8860 9496 8888
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 9876 8888 9904 8919
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 10594 8916 10600 8968
rect 10652 8916 10658 8968
rect 10612 8888 10640 8916
rect 9876 8860 10640 8888
rect 4356 8792 4936 8820
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 9674 8780 9680 8832
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 9824 8792 9965 8820
rect 9824 8780 9830 8792
rect 9953 8789 9965 8792
rect 9999 8789 10011 8823
rect 9953 8783 10011 8789
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 3050 8576 3056 8628
rect 3108 8576 3114 8628
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8616 3295 8619
rect 3878 8616 3884 8628
rect 3283 8588 3884 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4126 8588 6316 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 2700 8548 2728 8576
rect 1811 8520 2728 8548
rect 3068 8548 3096 8576
rect 4126 8548 4154 8588
rect 3068 8520 4154 8548
rect 4976 8551 5034 8557
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 4976 8517 4988 8551
rect 5022 8548 5034 8551
rect 5442 8548 5448 8560
rect 5022 8520 5448 8548
rect 5022 8517 5034 8520
rect 4976 8511 5034 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6288 8548 6316 8588
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7374 8616 7380 8628
rect 7147 8588 7380 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 9248 8551 9306 8557
rect 6288 8520 8892 8548
rect 2682 8480 2688 8492
rect 2148 8452 2688 8480
rect 2148 8421 2176 8452
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 2958 8489 2964 8492
rect 2953 8480 2964 8489
rect 2919 8452 2964 8480
rect 2953 8443 2964 8452
rect 2958 8440 2964 8443
rect 3016 8440 3022 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3970 8480 3976 8492
rect 3099 8452 3976 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4338 8440 4344 8492
rect 4396 8489 4402 8492
rect 4396 8443 4408 8489
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7650 8480 7656 8492
rect 7607 8452 7656 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 4396 8440 4402 8443
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7926 8480 7932 8492
rect 7791 8452 7932 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 8864 8480 8892 8520
rect 9248 8517 9260 8551
rect 9294 8548 9306 8551
rect 9674 8548 9680 8560
rect 9294 8520 9680 8548
rect 9294 8517 9306 8520
rect 9248 8511 9306 8517
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 9766 8480 9772 8492
rect 8864 8452 9772 8480
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 2038 8304 2044 8356
rect 2096 8344 2102 8356
rect 2332 8344 2360 8375
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4672 8384 4721 8412
rect 4672 8372 4678 8384
rect 4709 8381 4721 8384
rect 4755 8381 4767 8415
rect 6362 8412 6368 8424
rect 4709 8375 4767 8381
rect 6104 8384 6368 8412
rect 3142 8344 3148 8356
rect 2096 8316 2360 8344
rect 2608 8316 3148 8344
rect 2096 8304 2102 8316
rect 750 8236 756 8288
rect 808 8276 814 8288
rect 2608 8276 2636 8316
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 6104 8353 6132 8384
rect 6362 8372 6368 8384
rect 6420 8412 6426 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6420 8384 6929 8412
rect 6420 8372 6426 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8313 6147 8347
rect 6089 8307 6147 8313
rect 808 8248 2636 8276
rect 2685 8279 2743 8285
rect 808 8236 814 8248
rect 2685 8245 2697 8279
rect 2731 8276 2743 8279
rect 2866 8276 2872 8288
rect 2731 8248 2872 8276
rect 2731 8245 2743 8248
rect 2685 8239 2743 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8570 8276 8576 8288
rect 8159 8248 8576 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 9677 8279 9735 8285
rect 9677 8245 9689 8279
rect 9723 8276 9735 8279
rect 9858 8276 9864 8288
rect 9723 8248 9864 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 10502 8276 10508 8288
rect 10459 8248 10508 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4396 8044 4445 8072
rect 4396 8032 4402 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 4982 8032 4988 8084
rect 5040 8032 5046 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7558 8072 7564 8084
rect 7331 8044 7564 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7558 8032 7564 8044
rect 7616 8072 7622 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7616 8044 7757 8072
rect 7616 8032 7622 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 9858 8032 9864 8084
rect 9916 8032 9922 8084
rect 3421 8007 3479 8013
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 3467 7976 3832 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 3804 7948 3832 7976
rect 3786 7896 3792 7948
rect 3844 7896 3850 7948
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 6227 7908 7573 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 9876 7936 9904 8032
rect 9815 7908 9904 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2774 7868 2780 7880
rect 2087 7840 2780 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 3292 7840 5181 7868
rect 3292 7828 3298 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6362 7868 6368 7880
rect 6135 7840 6368 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6512 7840 6653 7868
rect 6512 7828 6518 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6788 7840 6837 7868
rect 6788 7828 6794 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 8628 7840 8708 7868
rect 8628 7828 8634 7840
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1397 7803 1455 7809
rect 1397 7800 1409 7803
rect 992 7772 1409 7800
rect 992 7760 998 7772
rect 1397 7769 1409 7772
rect 1443 7769 1455 7803
rect 1397 7763 1455 7769
rect 1765 7803 1823 7809
rect 1765 7769 1777 7803
rect 1811 7769 1823 7803
rect 1765 7763 1823 7769
rect 1780 7732 1808 7763
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2286 7803 2344 7809
rect 2286 7800 2298 7803
rect 2188 7772 2298 7800
rect 2188 7760 2194 7772
rect 2286 7769 2298 7772
rect 2332 7769 2344 7803
rect 2286 7763 2344 7769
rect 8680 7744 8708 7840
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9088 7840 9597 7868
rect 9088 7828 9094 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9907 7840 9996 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 9968 7744 9996 7840
rect 10060 7840 10241 7868
rect 5442 7732 5448 7744
rect 1780 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 8662 7692 8668 7744
rect 8720 7692 8726 7744
rect 8754 7692 8760 7744
rect 8812 7692 8818 7744
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 9950 7692 9956 7744
rect 10008 7692 10014 7744
rect 10060 7741 10088 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2130 7528 2136 7540
rect 2087 7500 2136 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 3292 7500 3525 7528
rect 3292 7488 3298 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 3786 7488 3792 7540
rect 3844 7488 3850 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 4982 7528 4988 7540
rect 4663 7500 4988 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5077 7531 5135 7537
rect 5077 7497 5089 7531
rect 5123 7528 5135 7531
rect 5350 7528 5356 7540
rect 5123 7500 5356 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 9030 7488 9036 7540
rect 9088 7488 9094 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 9180 7500 9229 7528
rect 9180 7488 9186 7500
rect 9217 7497 9229 7500
rect 9263 7497 9275 7531
rect 9217 7491 9275 7497
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 1544 7364 2881 7392
rect 1544 7352 1550 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3804 7392 3832 7488
rect 8018 7460 8024 7472
rect 5920 7432 8024 7460
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3467 7364 3893 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3050 7324 3056 7336
rect 2823 7296 3056 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 2608 7256 2636 7287
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3160 7324 3188 7355
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5920 7401 5948 7432
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 8662 7460 8668 7472
rect 8588 7432 8668 7460
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5675 7364 5917 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6178 7392 6184 7404
rect 6043 7364 6184 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 3160 7296 3740 7324
rect 3712 7265 3740 7296
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4982 7324 4988 7336
rect 4755 7296 4988 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 2961 7259 3019 7265
rect 2961 7256 2973 7259
rect 2608 7228 2973 7256
rect 2961 7225 2973 7228
rect 3007 7225 3019 7259
rect 2961 7219 3019 7225
rect 3329 7259 3387 7265
rect 3329 7225 3341 7259
rect 3375 7256 3387 7259
rect 3697 7259 3755 7265
rect 3375 7228 3648 7256
rect 3375 7225 3387 7228
rect 3329 7219 3387 7225
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2866 7188 2872 7200
rect 2455 7160 2872 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3620 7188 3648 7228
rect 3697 7225 3709 7259
rect 3743 7225 3755 7259
rect 3697 7219 3755 7225
rect 4172 7188 4200 7287
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 6012 7256 6040 7355
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6546 7392 6552 7404
rect 6411 7364 6552 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 8588 7401 8616 7432
rect 8662 7420 8668 7432
rect 8720 7460 8726 7472
rect 8720 7432 10272 7460
rect 8720 7420 8726 7432
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 8573 7395 8631 7401
rect 6687 7364 8432 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7324 6147 7327
rect 6454 7324 6460 7336
rect 6135 7296 6460 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 6454 7284 6460 7296
rect 6512 7324 6518 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6512 7296 6929 7324
rect 6512 7284 6518 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 4356 7228 6040 7256
rect 6549 7259 6607 7265
rect 4356 7200 4384 7228
rect 6549 7225 6561 7259
rect 6595 7256 6607 7259
rect 6730 7256 6736 7268
rect 6595 7228 6736 7256
rect 6595 7225 6607 7228
rect 6549 7219 6607 7225
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 6825 7259 6883 7265
rect 6825 7225 6837 7259
rect 6871 7256 6883 7259
rect 7116 7256 7144 7287
rect 6871 7228 7144 7256
rect 7300 7228 7696 7256
rect 6871 7225 6883 7228
rect 6825 7219 6883 7225
rect 3620 7160 4200 7188
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 5810 7148 5816 7200
rect 5868 7148 5874 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 7300 7188 7328 7228
rect 6696 7160 7328 7188
rect 6696 7148 6702 7160
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 7668 7197 7696 7228
rect 8312 7200 8340 7287
rect 8404 7265 8432 7364
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7225 8447 7259
rect 8389 7219 8447 7225
rect 7653 7191 7711 7197
rect 7653 7157 7665 7191
rect 7699 7157 7711 7191
rect 7653 7151 7711 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8588 7188 8616 7355
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8812 7364 8861 7392
rect 8812 7352 8818 7364
rect 8849 7361 8861 7364
rect 8895 7361 8907 7395
rect 9950 7392 9956 7404
rect 8849 7355 8907 7361
rect 8956 7364 9956 7392
rect 8956 7336 8984 7364
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10244 7401 10272 7432
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9907 7296 10057 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 9692 7256 9720 7287
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 9692 7228 10333 7256
rect 10321 7225 10333 7228
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 8352 7160 8616 7188
rect 8352 7148 8358 7160
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 1486 6984 1492 6996
rect 1443 6956 1492 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 7745 6987 7803 6993
rect 7745 6984 7757 6987
rect 7616 6956 7757 6984
rect 7616 6944 7622 6956
rect 7745 6953 7757 6956
rect 7791 6953 7803 6987
rect 7745 6947 7803 6953
rect 9122 6944 9128 6996
rect 9180 6944 9186 6996
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10134 6984 10140 6996
rect 10091 6956 10140 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 10459 6956 10916 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 4522 6916 4528 6928
rect 4126 6888 4528 6916
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 4126 6848 4154 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6916 5135 6919
rect 5718 6916 5724 6928
rect 5123 6888 5724 6916
rect 5123 6885 5135 6888
rect 5077 6879 5135 6885
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 2832 6820 4154 6848
rect 4709 6851 4767 6857
rect 2832 6808 2838 6820
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 4982 6848 4988 6860
rect 4755 6820 4988 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5810 6848 5816 6860
rect 5491 6820 5816 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 9140 6848 9168 6944
rect 10888 6928 10916 6956
rect 10870 6876 10876 6928
rect 10928 6876 10934 6928
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 9140 6820 9229 6848
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3292 6752 3525 6780
rect 3292 6740 3298 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3988 6752 4537 6780
rect 2532 6715 2590 6721
rect 2532 6681 2544 6715
rect 2578 6712 2590 6715
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2578 6684 2973 6712
rect 2578 6681 2590 6684
rect 2532 6675 2590 6681
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 3988 6653 4016 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5626 6780 5632 6792
rect 5307 6752 5632 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7607 6752 8217 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8619 6752 8984 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4798 6712 4804 6724
rect 4120 6684 4804 6712
rect 4120 6672 4126 6684
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 8312 6712 8340 6740
rect 7944 6684 8340 6712
rect 7944 6656 7972 6684
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6613 4031 6647
rect 3973 6607 4031 6613
rect 6822 6604 6828 6656
rect 6880 6604 6886 6656
rect 7926 6604 7932 6656
rect 7984 6604 7990 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8956 6653 8984 6752
rect 9048 6752 9137 6780
rect 9048 6656 9076 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9364 6752 9413 6780
rect 9364 6740 9370 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 9968 6656 9996 6743
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8720 6616 8769 6644
rect 8720 6604 8726 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9030 6604 9036 6656
rect 9088 6604 9094 6656
rect 9858 6604 9864 6656
rect 9916 6604 9922 6656
rect 9950 6604 9956 6656
rect 10008 6604 10014 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 2096 6412 2145 6440
rect 2096 6400 2102 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 4062 6440 4068 6452
rect 2740 6412 4068 6440
rect 2740 6400 2746 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 4856 6412 5549 6440
rect 4856 6400 4862 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7374 6440 7380 6452
rect 7239 6412 7380 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 9306 6440 9312 6452
rect 8987 6412 9312 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 6365 6375 6423 6381
rect 6365 6372 6377 6375
rect 4580 6344 5028 6372
rect 4580 6332 4586 6344
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 1811 6276 1900 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 1872 6168 1900 6276
rect 1946 6264 1952 6316
rect 2004 6264 2010 6316
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2406 6304 2412 6316
rect 2096 6276 2412 6304
rect 2096 6264 2102 6276
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3160 6276 3433 6304
rect 3160 6248 3188 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4729 6307 4787 6313
rect 4729 6273 4741 6307
rect 4775 6304 4787 6307
rect 4890 6304 4896 6316
rect 4775 6276 4896 6304
rect 4775 6273 4787 6276
rect 4729 6267 4787 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5000 6313 5028 6344
rect 6196 6344 6377 6372
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 3142 6196 3148 6248
rect 3200 6196 3206 6248
rect 3234 6196 3240 6248
rect 3292 6196 3298 6248
rect 5276 6168 5304 6267
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6196 6313 6224 6344
rect 6365 6341 6377 6344
rect 6411 6341 6423 6375
rect 6365 6335 6423 6341
rect 7576 6344 8892 6372
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 5776 6276 6193 6304
rect 5776 6264 5782 6276
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6304 7159 6307
rect 7466 6304 7472 6316
rect 7147 6276 7472 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7576 6313 7604 6344
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 8864 6313 8892 6344
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7708 6276 7849 6304
rect 7708 6264 7714 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 7837 6267 7895 6273
rect 7944 6276 8769 6304
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5408 6208 6009 6236
rect 5408 6196 5414 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6362 6196 6368 6248
rect 6420 6236 6426 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6420 6208 6837 6236
rect 6420 6196 6426 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6972 6208 7021 6236
rect 6972 6196 6978 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7745 6171 7803 6177
rect 1872 6140 4108 6168
rect 5276 6140 5764 6168
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2590 6100 2596 6112
rect 2363 6072 2596 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 2682 6060 2688 6112
rect 2740 6060 2746 6112
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3384 6072 3617 6100
rect 3384 6060 3390 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 4080 6100 4108 6140
rect 5736 6112 5764 6140
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 7944 6168 7972 6276
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 8938 6304 8944 6316
rect 8895 6276 8944 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9263 6276 9965 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10100 6276 10241 6304
rect 10100 6264 10106 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 7791 6140 7972 6168
rect 8036 6168 8064 6199
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 8720 6208 9413 6236
rect 8720 6196 8726 6208
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 8036 6140 8585 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 8573 6131 8631 6137
rect 5074 6100 5080 6112
rect 4080 6072 5080 6100
rect 3605 6063 3663 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5442 6060 5448 6112
rect 5500 6060 5506 6112
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2133 5899 2191 5905
rect 2133 5896 2145 5899
rect 2004 5868 2145 5896
rect 2004 5856 2010 5868
rect 2133 5865 2145 5868
rect 2179 5865 2191 5899
rect 2133 5859 2191 5865
rect 2590 5856 2596 5908
rect 2648 5856 2654 5908
rect 2682 5856 2688 5908
rect 2740 5856 2746 5908
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3786 5896 3792 5908
rect 3651 5868 3792 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4893 5899 4951 5905
rect 4893 5865 4905 5899
rect 4939 5896 4951 5899
rect 4982 5896 4988 5908
rect 4939 5868 4988 5896
rect 4939 5865 4951 5868
rect 4893 5859 4951 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5350 5856 5356 5908
rect 5408 5856 5414 5908
rect 5442 5856 5448 5908
rect 5500 5856 5506 5908
rect 5626 5856 5632 5908
rect 5684 5856 5690 5908
rect 5905 5899 5963 5905
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6362 5896 6368 5908
rect 5951 5868 6368 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 6914 5896 6920 5908
rect 6871 5868 6920 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 10042 5896 10048 5908
rect 7883 5868 10048 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 2501 5831 2559 5837
rect 2501 5797 2513 5831
rect 2547 5797 2559 5831
rect 2501 5791 2559 5797
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1728 5664 1961 5692
rect 1728 5652 1734 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2516 5692 2544 5791
rect 2608 5769 2636 5856
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2700 5760 2728 5856
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2700 5732 2789 5760
rect 2593 5723 2651 5729
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 3252 5692 3280 5856
rect 4709 5831 4767 5837
rect 4709 5797 4721 5831
rect 4755 5828 4767 5831
rect 5368 5828 5396 5856
rect 4755 5800 5396 5828
rect 4755 5797 4767 5800
rect 4709 5791 4767 5797
rect 5460 5760 5488 5856
rect 5644 5828 5672 5856
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 5644 5800 6101 5828
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 8478 5788 8484 5840
rect 8536 5788 8542 5840
rect 8496 5760 8524 5788
rect 8662 5760 8668 5772
rect 5460 5732 6316 5760
rect 8496 5732 8668 5760
rect 2516 5664 3280 5692
rect 2317 5655 2375 5661
rect 1486 5584 1492 5636
rect 1544 5584 1550 5636
rect 2332 5624 2360 5655
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 3384 5664 3433 5692
rect 3384 5652 3390 5664
rect 3421 5661 3433 5664
rect 3467 5692 3479 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3467 5664 3985 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3973 5661 3985 5664
rect 4019 5692 4031 5695
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4019 5664 4629 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5718 5692 5724 5704
rect 5491 5664 5724 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5460 5624 5488 5655
rect 5718 5652 5724 5664
rect 5776 5692 5782 5704
rect 6288 5701 6316 5732
rect 8662 5720 8668 5732
rect 8720 5760 8726 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8720 5732 9045 5760
rect 8720 5720 8726 5732
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9950 5760 9956 5772
rect 9723 5732 9956 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9950 5720 9956 5732
rect 10008 5760 10014 5772
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 10008 5732 10149 5760
rect 10008 5720 10014 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5776 5664 5825 5692
rect 5776 5652 5782 5664
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 2332 5596 3832 5624
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3804 5565 3832 5596
rect 4448 5596 5488 5624
rect 6932 5624 6960 5655
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 8205 5695 8263 5701
rect 7699 5664 7788 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7760 5624 7788 5664
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8251 5664 8524 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 6932 5596 7788 5624
rect 4448 5568 4476 5596
rect 7760 5568 7788 5596
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 8076 5596 8401 5624
rect 8076 5584 8082 5596
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8496 5624 8524 5664
rect 9030 5624 9036 5636
rect 8496 5596 9036 5624
rect 8389 5587 8447 5593
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 9858 5584 9864 5636
rect 9916 5584 9922 5636
rect 9950 5584 9956 5636
rect 10008 5584 10014 5636
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 3200 5528 3249 5556
rect 3200 5516 3206 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 3237 5519 3295 5525
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4430 5516 4436 5568
rect 4488 5516 4494 5568
rect 7558 5516 7564 5568
rect 7616 5516 7622 5568
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 8665 5559 8723 5565
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 10318 5556 10324 5568
rect 8711 5528 10324 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 2498 5312 2504 5364
rect 2556 5312 2562 5364
rect 6822 5352 6828 5364
rect 4356 5324 6828 5352
rect 3234 5284 3240 5296
rect 2240 5256 3240 5284
rect 1762 5176 1768 5228
rect 1820 5176 1826 5228
rect 2240 5225 2268 5256
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 4356 5293 4384 5324
rect 6822 5312 6828 5324
rect 6880 5352 6886 5364
rect 6880 5312 6914 5352
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5253 4399 5287
rect 5353 5287 5411 5293
rect 5353 5284 5365 5287
rect 4341 5247 4399 5253
rect 5092 5256 5365 5284
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4617 5179 4675 5185
rect 4816 5188 4905 5216
rect 2332 5148 2360 5179
rect 4430 5148 4436 5160
rect 1872 5120 4436 5148
rect 1872 5024 1900 5120
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 1854 4972 1860 5024
rect 1912 4972 1918 5024
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2498 5012 2504 5024
rect 2179 4984 2504 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 4522 5012 4528 5024
rect 3099 4984 4528 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 4632 5012 4660 5179
rect 4816 5089 4844 5188
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 5092 5089 5120 5256
rect 5353 5253 5365 5256
rect 5399 5253 5411 5287
rect 6886 5284 6914 5312
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 5353 5247 5411 5253
rect 6380 5256 6776 5284
rect 6886 5256 7849 5284
rect 6380 5225 6408 5256
rect 6638 5225 6644 5228
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6632 5216 6644 5225
rect 6599 5188 6644 5216
rect 6365 5179 6423 5185
rect 6632 5179 6644 5188
rect 6638 5176 6644 5179
rect 6696 5176 6702 5228
rect 6748 5216 6776 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 7837 5247 7895 5253
rect 9398 5216 9404 5228
rect 6748 5188 9404 5216
rect 9398 5176 9404 5188
rect 9456 5216 9462 5228
rect 10226 5216 10232 5228
rect 9456 5188 10232 5216
rect 9456 5176 9462 5188
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5307 5120 6009 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5997 5117 6009 5120
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 9214 5148 9220 5160
rect 7616 5120 9220 5148
rect 7616 5108 7622 5120
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 4801 5083 4859 5089
rect 4801 5049 4813 5083
rect 4847 5049 4859 5083
rect 4801 5043 4859 5049
rect 5077 5083 5135 5089
rect 5077 5049 5089 5083
rect 5123 5049 5135 5083
rect 5077 5043 5135 5049
rect 5813 5083 5871 5089
rect 5813 5049 5825 5083
rect 5859 5080 5871 5083
rect 6178 5080 6184 5092
rect 5859 5052 6184 5080
rect 5859 5049 5871 5052
rect 5813 5043 5871 5049
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 7745 5083 7803 5089
rect 7745 5049 7757 5083
rect 7791 5080 7803 5083
rect 8938 5080 8944 5092
rect 7791 5052 8944 5080
rect 7791 5049 7803 5052
rect 7745 5043 7803 5049
rect 8938 5040 8944 5052
rect 8996 5080 9002 5092
rect 9692 5080 9720 5111
rect 8996 5052 9720 5080
rect 8996 5040 9002 5052
rect 5166 5012 5172 5024
rect 4632 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 10100 4984 10333 5012
rect 10100 4972 10106 4984
rect 10321 4981 10333 4984
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1486 4808 1492 4820
rect 1443 4780 1492 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1486 4768 1492 4780
rect 1544 4768 1550 4820
rect 4338 4808 4344 4820
rect 1596 4780 4344 4808
rect 1596 4613 1624 4780
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5776 4780 5917 4808
rect 5776 4768 5782 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 9122 4808 9128 4820
rect 8711 4780 9128 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 2498 4700 2504 4752
rect 2556 4700 2562 4752
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 4157 4743 4215 4749
rect 4157 4740 4169 4743
rect 2639 4712 4169 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2516 4672 2544 4700
rect 2869 4675 2927 4681
rect 2869 4672 2881 4675
rect 2516 4644 2881 4672
rect 2869 4641 2881 4644
rect 2915 4641 2927 4675
rect 2869 4635 2927 4641
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 1688 4468 1716 4564
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 1964 4536 1992 4567
rect 2038 4564 2044 4616
rect 2096 4604 2102 4616
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 2096 4576 2145 4604
rect 2096 4564 2102 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2976 4604 3004 4712
rect 4157 4709 4169 4712
rect 4203 4709 4215 4743
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 4157 4703 4215 4709
rect 7392 4712 8953 4740
rect 7392 4684 7420 4712
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 3108 4644 3341 4672
rect 3108 4632 3114 4644
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3436 4644 4108 4672
rect 2731 4576 3004 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3436 4613 3464 4644
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3292 4576 3433 4604
rect 3292 4564 3298 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 3878 4604 3884 4616
rect 3835 4576 3884 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 4080 4604 4108 4644
rect 4522 4632 4528 4684
rect 4580 4632 4586 4684
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 7558 4672 7564 4684
rect 7515 4644 7564 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7558 4632 7564 4644
rect 7616 4672 7622 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7616 4644 7849 4672
rect 7616 4632 7622 4644
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 7837 4635 7895 4641
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8110 4672 8116 4684
rect 8067 4644 8116 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 4080 4576 4154 4604
rect 3973 4567 4031 4573
rect 1811 4508 2728 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 2700 4480 2728 4508
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3988 4536 4016 4567
rect 2924 4508 4016 4536
rect 2924 4496 2930 4508
rect 2590 4468 2596 4480
rect 1688 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 2682 4428 2688 4480
rect 2740 4428 2746 4480
rect 3605 4471 3663 4477
rect 3605 4437 3617 4471
rect 3651 4468 3663 4471
rect 3786 4468 3792 4480
rect 3651 4440 3792 4468
rect 3651 4437 3663 4440
rect 3605 4431 3663 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4126 4468 4154 4576
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5132 4576 6101 4604
rect 5132 4564 5138 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6638 4604 6644 4616
rect 6089 4567 6147 4573
rect 6196 4576 6644 4604
rect 4792 4539 4850 4545
rect 4792 4505 4804 4539
rect 4838 4536 4850 4539
rect 4982 4536 4988 4548
rect 4838 4508 4988 4536
rect 4838 4505 4850 4508
rect 4792 4499 4850 4505
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 6196 4468 6224 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 7926 4604 7932 4616
rect 7791 4576 7932 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 7760 4536 7788 4567
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8404 4604 8432 4712
rect 8941 4709 8953 4712
rect 8987 4740 8999 4743
rect 9030 4740 9036 4752
rect 8987 4712 9036 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8662 4672 8668 4684
rect 8527 4644 8668 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8404 4576 8585 4604
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 10042 4564 10048 4616
rect 10100 4613 10106 4616
rect 10100 4604 10112 4613
rect 10100 4576 10145 4604
rect 10100 4567 10112 4576
rect 10100 4564 10106 4567
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10284 4576 10333 4604
rect 10284 4564 10290 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 6886 4508 7788 4536
rect 4126 4440 6224 4468
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6886 4468 6914 4508
rect 6604 4440 6914 4468
rect 6604 4428 6610 4440
rect 7650 4428 7656 4480
rect 7708 4428 7714 4480
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 1949 4267 2007 4273
rect 1949 4264 1961 4267
rect 1820 4236 1961 4264
rect 1820 4224 1826 4236
rect 1949 4233 1961 4236
rect 1995 4233 2007 4267
rect 1949 4227 2007 4233
rect 3234 4224 3240 4276
rect 3292 4224 3298 4276
rect 3786 4264 3792 4276
rect 3620 4236 3792 4264
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2148 3992 2176 4091
rect 2608 4060 2636 4091
rect 2682 4088 2688 4140
rect 2740 4088 2746 4140
rect 3252 4128 3280 4224
rect 3620 4137 3648 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 5074 4224 5080 4276
rect 5132 4224 5138 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 4522 4196 4528 4208
rect 3804 4168 4528 4196
rect 3804 4137 3832 4168
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 2792 4100 3280 4128
rect 3605 4131 3663 4137
rect 2792 4060 2820 4100
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 4056 4131 4114 4137
rect 4056 4097 4068 4131
rect 4102 4128 4114 4131
rect 5092 4128 5120 4224
rect 5442 4156 5448 4208
rect 5500 4156 5506 4208
rect 4102 4100 5120 4128
rect 4102 4097 4114 4100
rect 4056 4091 4114 4097
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6748 4128 6776 4227
rect 7006 4224 7012 4276
rect 7064 4224 7070 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7616 4236 7757 4264
rect 7616 4224 7622 4236
rect 7745 4233 7757 4236
rect 7791 4233 7803 4267
rect 7745 4227 7803 4233
rect 8018 4224 8024 4276
rect 8076 4224 8082 4276
rect 8757 4267 8815 4273
rect 8757 4233 8769 4267
rect 8803 4264 8815 4267
rect 10410 4264 10416 4276
rect 8803 4236 10416 4264
rect 8803 4233 8815 4236
rect 8757 4227 8815 4233
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6748 4100 6837 4128
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7650 4128 7656 4140
rect 7331 4100 7656 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 2608 4032 2820 4060
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 5353 4063 5411 4069
rect 2915 4032 3464 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 2958 3992 2964 4004
rect 2148 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3436 4001 3464 4032
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3961 3479 3995
rect 3421 3955 3479 3961
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 992 3896 1501 3924
rect 992 3884 998 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 2498 3884 2504 3936
rect 2556 3884 2562 3936
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 5368 3924 5396 4023
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7101 4063 7159 4069
rect 7101 4060 7113 4063
rect 6972 4032 7113 4060
rect 6972 4020 6978 4032
rect 7101 4029 7113 4032
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7852 4060 7880 4091
rect 7432 4032 7880 4060
rect 7432 4020 7438 4032
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3961 5963 3995
rect 5905 3955 5963 3961
rect 3384 3896 5396 3924
rect 5920 3924 5948 3955
rect 6178 3924 6184 3936
rect 5920 3896 6184 3924
rect 3384 3884 3390 3896
rect 6178 3884 6184 3896
rect 6236 3924 6242 3936
rect 8680 3924 8708 4091
rect 10042 4088 10048 4140
rect 10100 4137 10106 4140
rect 10100 4091 10112 4137
rect 10100 4088 10106 4091
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10321 4131 10379 4137
rect 10321 4128 10333 4131
rect 10284 4100 10333 4128
rect 10284 4088 10290 4100
rect 10321 4097 10333 4100
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 8938 3952 8944 4004
rect 8996 3952 9002 4004
rect 6236 3896 8708 3924
rect 6236 3884 6242 3896
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 1820 3692 2421 3720
rect 1820 3680 1826 3692
rect 2409 3689 2421 3692
rect 2455 3689 2467 3723
rect 2409 3683 2467 3689
rect 2498 3680 2504 3732
rect 2556 3680 2562 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2866 3720 2872 3732
rect 2648 3692 2872 3720
rect 2648 3680 2654 3692
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3326 3680 3332 3732
rect 3384 3680 3390 3732
rect 4982 3680 4988 3732
rect 5040 3680 5046 3732
rect 5442 3680 5448 3732
rect 5500 3680 5506 3732
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6972 3692 7205 3720
rect 6972 3680 6978 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9677 3723 9735 3729
rect 9088 3692 9628 3720
rect 9088 3680 9094 3692
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 2516 3584 2544 3680
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 4062 3652 4068 3664
rect 3016 3624 4068 3652
rect 3016 3612 3022 3624
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 5460 3652 5488 3680
rect 4847 3624 5488 3652
rect 5905 3655 5963 3661
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 5905 3621 5917 3655
rect 5951 3621 5963 3655
rect 5905 3615 5963 3621
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2004 3556 2268 3584
rect 2516 3556 2881 3584
rect 2004 3544 2010 3556
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 1912 3488 2145 3516
rect 1912 3476 1918 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2240 3516 2268 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 3160 3556 3924 3584
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2240 3488 2605 3516
rect 2133 3479 2191 3485
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 3160 3516 3188 3556
rect 3896 3528 3924 3556
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 5920 3584 5948 3615
rect 4396 3556 5856 3584
rect 5920 3556 9536 3584
rect 4396 3544 4402 3556
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 2731 3488 3188 3516
rect 3252 3488 3801 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 992 3420 1409 3448
rect 992 3408 998 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 1397 3411 1455 3417
rect 1765 3451 1823 3457
rect 1765 3417 1777 3451
rect 1811 3448 1823 3451
rect 2958 3448 2964 3460
rect 1811 3420 2964 3448
rect 1811 3417 1823 3420
rect 1765 3411 1823 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 3252 3392 3280 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3878 3476 3884 3528
rect 3936 3476 3942 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 5166 3516 5172 3528
rect 4755 3488 5172 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 5166 3476 5172 3488
rect 5224 3516 5230 3528
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5224 3488 5549 3516
rect 5224 3476 5230 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5828 3516 5856 3556
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 5828 3488 7297 3516
rect 5721 3479 5779 3485
rect 7285 3485 7297 3488
rect 7331 3516 7343 3519
rect 7331 3488 9076 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 5258 3448 5264 3460
rect 4448 3420 5264 3448
rect 4448 3392 4476 3420
rect 5258 3408 5264 3420
rect 5316 3448 5322 3460
rect 5736 3448 5764 3479
rect 5316 3420 5764 3448
rect 5316 3408 5322 3420
rect 9048 3392 9076 3488
rect 9214 3476 9220 3528
rect 9272 3476 9278 3528
rect 9508 3525 9536 3556
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9600 3516 9628 3692
rect 9677 3689 9689 3723
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 9692 3596 9720 3683
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 10100 3692 10517 3720
rect 10100 3680 10106 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 9674 3544 9680 3596
rect 9732 3544 9738 3596
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9600 3488 9873 3516
rect 9493 3479 9551 3485
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 2314 3380 2320 3392
rect 2271 3352 2320 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 3234 3340 3240 3392
rect 3292 3340 3298 3392
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 9030 3340 9036 3392
rect 9088 3340 9094 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9968 3380 9996 3476
rect 9447 3352 9996 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 1596 3108 1624 3139
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 2096 3148 2237 3176
rect 2096 3136 2102 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 2746 3148 3004 3176
rect 2332 3108 2360 3136
rect 2746 3108 2774 3148
rect 1596 3080 2084 3108
rect 2332 3080 2774 3108
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1443 3012 1777 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1765 3009 1777 3012
rect 1811 3040 1823 3043
rect 1854 3040 1860 3052
rect 1811 3012 1860 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 2056 3049 2084 3080
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 2976 3049 3004 3148
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 3200 3148 3433 3176
rect 3200 3136 3206 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 4062 3176 4068 3188
rect 3835 3148 4068 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 3712 3108 3740 3139
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3145 8999 3179
rect 8941 3139 8999 3145
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 10410 3176 10416 3188
rect 9723 3148 10416 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 8956 3108 8984 3139
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 3160 3080 3648 3108
rect 3712 3080 4154 3108
rect 8956 3080 9413 3108
rect 3160 3052 3188 3080
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 2961 3043 3019 3049
rect 2823 3012 2912 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 2884 2972 2912 3012
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3142 3000 3148 3052
rect 3200 3000 3206 3052
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3292 3012 3525 3040
rect 3292 3000 3298 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3620 3040 3648 3080
rect 3786 3040 3792 3052
rect 3620 3012 3792 3040
rect 3513 3003 3571 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 3970 3000 3976 3052
rect 4028 3000 4034 3052
rect 3896 2972 3924 3000
rect 2884 2944 3924 2972
rect 4126 2972 4154 3080
rect 9401 3077 9413 3080
rect 9447 3077 9459 3111
rect 9401 3071 9459 3077
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 7466 3040 7472 3052
rect 5684 3012 7472 3040
rect 5684 3000 5690 3012
rect 7466 3000 7472 3012
rect 7524 3040 7530 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7524 3012 8769 3040
rect 7524 3000 7530 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 9968 2972 9996 3003
rect 4126 2944 9996 2972
rect 8938 2904 8944 2916
rect 2700 2876 8944 2904
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2836 1915 2839
rect 2590 2836 2596 2848
rect 1903 2808 2596 2836
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 2700 2845 2728 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 9214 2796 9220 2848
rect 9272 2796 9278 2848
rect 10226 2796 10232 2848
rect 10284 2796 10290 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2556 2604 2697 2632
rect 2556 2592 2562 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 2685 2595 2743 2601
rect 2700 2564 2728 2595
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 5534 2632 5540 2644
rect 2832 2604 5540 2632
rect 2832 2592 2838 2604
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7374 2632 7380 2644
rect 6871 2604 7380 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7800 2604 7849 2632
rect 7800 2592 7806 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2632 8815 2635
rect 8846 2632 8852 2644
rect 8803 2604 8852 2632
rect 8803 2601 8815 2604
rect 8757 2595 8815 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9493 2635 9551 2641
rect 9493 2601 9505 2635
rect 9539 2632 9551 2635
rect 10042 2632 10048 2644
rect 9539 2604 10048 2632
rect 9539 2601 9551 2604
rect 9493 2595 9551 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 2700 2536 3188 2564
rect 1780 2468 2636 2496
rect 1780 2437 1808 2468
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 992 2332 1409 2360
rect 992 2320 998 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2130 2252 2136 2304
rect 2188 2252 2194 2304
rect 2240 2292 2268 2391
rect 2498 2388 2504 2440
rect 2556 2388 2562 2440
rect 2608 2428 2636 2468
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 3160 2496 3188 2536
rect 3234 2524 3240 2576
rect 3292 2524 3298 2576
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2564 4031 2567
rect 4338 2564 4344 2576
rect 4019 2536 4344 2564
rect 4019 2533 4031 2536
rect 3973 2527 4031 2533
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 4430 2524 4436 2576
rect 4488 2524 4494 2576
rect 10134 2564 10140 2576
rect 8588 2536 10140 2564
rect 2740 2468 3004 2496
rect 3160 2468 3372 2496
rect 2740 2456 2746 2468
rect 2866 2428 2872 2440
rect 2608 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 2976 2437 3004 2468
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 3142 2388 3148 2440
rect 3200 2388 3206 2440
rect 3344 2437 3372 2468
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 4246 2388 4252 2440
rect 4304 2388 4310 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8588 2437 8616 2536
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 8996 2468 9720 2496
rect 8996 2456 9002 2468
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9692 2437 9720 2468
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9232 2400 9321 2428
rect 3160 2360 3188 2388
rect 3421 2363 3479 2369
rect 3421 2360 3433 2363
rect 2608 2332 3096 2360
rect 3160 2332 3433 2360
rect 2608 2292 2636 2332
rect 2240 2264 2636 2292
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 2958 2292 2964 2304
rect 2823 2264 2964 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 3068 2292 3096 2332
rect 3421 2329 3433 2332
rect 3467 2329 3479 2363
rect 3421 2323 3479 2329
rect 3878 2320 3884 2372
rect 3936 2320 3942 2372
rect 3896 2292 3924 2320
rect 9232 2301 9260 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 9456 2332 10149 2360
rect 9456 2320 9462 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 10137 2323 10195 2329
rect 3068 2264 3924 2292
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9858 2252 9864 2304
rect 9916 2252 9922 2304
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 10502 2292 10508 2304
rect 10459 2264 10508 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 566 2048 572 2100
rect 624 2088 630 2100
rect 3786 2088 3792 2100
rect 624 2060 3792 2088
rect 624 2048 630 2060
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 2130 1980 2136 2032
rect 2188 2020 2194 2032
rect 6822 2020 6828 2032
rect 2188 1992 6828 2020
rect 2188 1980 2194 1992
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 1762 1368 1768 1420
rect 1820 1408 1826 1420
rect 2498 1408 2504 1420
rect 1820 1380 2504 1408
rect 1820 1368 1826 1380
rect 2498 1368 2504 1380
rect 2556 1368 2562 1420
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 940 9596 992 9648
rect 2044 9596 2096 9648
rect 3240 9596 3292 9648
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 2964 9460 3016 9512
rect 6184 9664 6236 9716
rect 7196 9664 7248 9716
rect 8668 9664 8720 9716
rect 9772 9664 9824 9716
rect 10324 9664 10376 9716
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 4620 9596 4672 9648
rect 7380 9528 7432 9580
rect 7748 9528 7800 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 3884 9460 3936 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 5908 9460 5960 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 2780 9324 2832 9376
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 6184 9324 6236 9376
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8024 9324 8076 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 1584 9120 1636 9172
rect 2504 9120 2556 9172
rect 3424 9120 3476 9172
rect 4252 9120 4304 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 4988 9120 5040 9172
rect 5080 9120 5132 9172
rect 1124 8984 1176 9036
rect 3056 8984 3108 9036
rect 2688 8823 2740 8832
rect 2688 8789 2697 8823
rect 2697 8789 2731 8823
rect 2731 8789 2740 8823
rect 2688 8780 2740 8789
rect 4160 9052 4212 9104
rect 5908 9052 5960 9104
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 4988 8984 5040 9036
rect 3884 8916 3936 8968
rect 5448 8916 5500 8968
rect 6736 9120 6788 9172
rect 7748 9120 7800 9172
rect 7840 9120 7892 9172
rect 9956 9120 10008 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 7380 9052 7432 9104
rect 7472 8984 7524 9036
rect 7840 8984 7892 9036
rect 11060 9052 11112 9104
rect 4160 8780 4212 8832
rect 6368 8891 6420 8900
rect 6368 8857 6402 8891
rect 6402 8857 6420 8891
rect 6368 8848 6420 8857
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 9496 8848 9548 8900
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10600 8916 10652 8968
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 9772 8780 9824 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 2688 8576 2740 8628
rect 3056 8576 3108 8628
rect 3884 8576 3936 8628
rect 5448 8508 5500 8560
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 7380 8576 7432 8628
rect 2688 8440 2740 8492
rect 2964 8483 3016 8492
rect 2964 8449 2965 8483
rect 2965 8449 2999 8483
rect 2999 8449 3016 8483
rect 2964 8440 3016 8449
rect 3976 8440 4028 8492
rect 4344 8483 4396 8492
rect 4344 8449 4362 8483
rect 4362 8449 4396 8483
rect 4344 8440 4396 8449
rect 7656 8440 7708 8492
rect 7932 8440 7984 8492
rect 9680 8508 9732 8560
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 2044 8304 2096 8356
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 756 8236 808 8288
rect 3148 8304 3200 8356
rect 6368 8372 6420 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 2872 8236 2924 8288
rect 8576 8236 8628 8288
rect 9864 8236 9916 8288
rect 10508 8236 10560 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 4344 8032 4396 8084
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 7564 8032 7616 8084
rect 9864 8032 9916 8084
rect 3792 7939 3844 7948
rect 3792 7905 3801 7939
rect 3801 7905 3835 7939
rect 3835 7905 3844 7939
rect 3792 7896 3844 7905
rect 2780 7828 2832 7880
rect 3240 7828 3292 7880
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6460 7828 6512 7880
rect 6736 7828 6788 7880
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 940 7760 992 7812
rect 2136 7760 2188 7812
rect 9036 7828 9088 7880
rect 5448 7692 5500 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 8668 7692 8720 7744
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 8760 7692 8812 7701
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9956 7692 10008 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 2136 7488 2188 7540
rect 3240 7488 3292 7540
rect 3792 7488 3844 7540
rect 4988 7488 5040 7540
rect 5356 7488 5408 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 9036 7531 9088 7540
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 9128 7488 9180 7540
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 3056 7284 3108 7336
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 8024 7420 8076 7472
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 2872 7148 2924 7200
rect 4988 7284 5040 7336
rect 6184 7352 6236 7404
rect 6552 7352 6604 7404
rect 8668 7420 8720 7472
rect 6460 7284 6512 7336
rect 6736 7216 6788 7268
rect 4344 7148 4396 7200
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 6644 7148 6696 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 8300 7148 8352 7200
rect 8760 7352 8812 7404
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 8944 7284 8996 7336
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 1492 6944 1544 6996
rect 7564 6944 7616 6996
rect 9128 6944 9180 6996
rect 10140 6944 10192 6996
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 4528 6876 4580 6928
rect 5724 6876 5776 6928
rect 2780 6808 2832 6817
rect 4988 6808 5040 6860
rect 5816 6808 5868 6860
rect 10876 6876 10928 6928
rect 3240 6740 3292 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 5632 6740 5684 6792
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 4068 6715 4120 6724
rect 4068 6681 4077 6715
rect 4077 6681 4111 6715
rect 4111 6681 4120 6715
rect 4068 6672 4120 6681
rect 4804 6672 4856 6724
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7932 6604 7984 6656
rect 8668 6604 8720 6656
rect 9312 6740 9364 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 9036 6604 9088 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 9956 6604 10008 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 2044 6400 2096 6452
rect 2688 6400 2740 6452
rect 4068 6400 4120 6452
rect 4804 6400 4856 6452
rect 7380 6400 7432 6452
rect 9312 6400 9364 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 4528 6332 4580 6384
rect 940 6264 992 6316
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2044 6264 2096 6316
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 4896 6264 4948 6316
rect 3148 6196 3200 6248
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 5724 6264 5776 6316
rect 7472 6264 7524 6316
rect 7656 6264 7708 6316
rect 5356 6196 5408 6248
rect 6368 6196 6420 6248
rect 6920 6196 6972 6248
rect 2596 6060 2648 6112
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3332 6060 3384 6112
rect 8944 6264 8996 6316
rect 10048 6264 10100 6316
rect 8668 6196 8720 6248
rect 5080 6060 5132 6112
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 5724 6060 5776 6112
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1952 5856 2004 5908
rect 2596 5856 2648 5908
rect 2688 5856 2740 5908
rect 3240 5856 3292 5908
rect 3792 5856 3844 5908
rect 4988 5856 5040 5908
rect 5356 5856 5408 5908
rect 5448 5856 5500 5908
rect 5632 5856 5684 5908
rect 6368 5856 6420 5908
rect 6920 5856 6972 5908
rect 10048 5856 10100 5908
rect 1676 5652 1728 5704
rect 8484 5788 8536 5840
rect 1492 5627 1544 5636
rect 1492 5593 1501 5627
rect 1501 5593 1535 5627
rect 1535 5593 1544 5627
rect 1492 5584 1544 5593
rect 3332 5652 3384 5704
rect 5724 5652 5776 5704
rect 8668 5720 8720 5772
rect 9956 5720 10008 5772
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 3148 5516 3200 5568
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 8024 5584 8076 5636
rect 9036 5584 9088 5636
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 9864 5627 9916 5636
rect 9864 5593 9873 5627
rect 9873 5593 9907 5627
rect 9907 5593 9916 5627
rect 9864 5584 9916 5593
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 4436 5516 4488 5568
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 7748 5516 7800 5568
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 10324 5516 10376 5568
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 3240 5244 3292 5296
rect 6828 5312 6880 5364
rect 4436 5108 4488 5160
rect 940 4972 992 5024
rect 1860 4972 1912 5024
rect 2504 4972 2556 5024
rect 4528 4972 4580 5024
rect 6644 5219 6696 5228
rect 6644 5185 6678 5219
rect 6678 5185 6696 5219
rect 6644 5176 6696 5185
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 10232 5176 10284 5228
rect 7564 5108 7616 5160
rect 9220 5108 9272 5160
rect 6184 5040 6236 5092
rect 8944 5040 8996 5092
rect 5172 4972 5224 5024
rect 10048 4972 10100 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 1492 4768 1544 4820
rect 4344 4768 4396 4820
rect 5724 4768 5776 4820
rect 9128 4768 9180 4820
rect 2504 4700 2556 4752
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 2044 4564 2096 4616
rect 3056 4632 3108 4684
rect 3240 4564 3292 4616
rect 3884 4564 3936 4616
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 7380 4632 7432 4684
rect 7564 4632 7616 4684
rect 8116 4632 8168 4684
rect 2872 4496 2924 4548
rect 2596 4428 2648 4480
rect 2688 4428 2740 4480
rect 3792 4428 3844 4480
rect 5080 4564 5132 4616
rect 6644 4607 6696 4616
rect 4988 4496 5040 4548
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7932 4564 7984 4616
rect 9036 4700 9088 4752
rect 8668 4632 8720 4684
rect 10048 4607 10100 4616
rect 10048 4573 10066 4607
rect 10066 4573 10100 4607
rect 10048 4564 10100 4573
rect 10232 4564 10284 4616
rect 6552 4428 6604 4480
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1768 4224 1820 4276
rect 3240 4224 3292 4276
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3792 4224 3844 4276
rect 5080 4224 5132 4276
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 4528 4156 4580 4208
rect 5448 4199 5500 4208
rect 5448 4165 5457 4199
rect 5457 4165 5491 4199
rect 5491 4165 5500 4199
rect 5448 4156 5500 4165
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 7564 4224 7616 4276
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 10416 4224 10468 4276
rect 7656 4088 7708 4140
rect 2964 3952 3016 4004
rect 940 3884 992 3936
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 6920 4020 6972 4072
rect 7380 4020 7432 4072
rect 3332 3884 3384 3893
rect 6184 3884 6236 3936
rect 10048 4131 10100 4140
rect 10048 4097 10066 4131
rect 10066 4097 10100 4131
rect 10048 4088 10100 4097
rect 10232 4088 10284 4140
rect 8944 3995 8996 4004
rect 8944 3961 8953 3995
rect 8953 3961 8987 3995
rect 8987 3961 8996 3995
rect 8944 3952 8996 3961
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 1768 3680 1820 3732
rect 2504 3680 2556 3732
rect 2596 3680 2648 3732
rect 2872 3680 2924 3732
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 5448 3680 5500 3732
rect 6920 3680 6972 3732
rect 9036 3680 9088 3732
rect 1952 3544 2004 3596
rect 2964 3612 3016 3664
rect 4068 3612 4120 3664
rect 1860 3476 1912 3528
rect 4344 3544 4396 3596
rect 940 3408 992 3460
rect 2964 3408 3016 3460
rect 3884 3476 3936 3528
rect 5172 3476 5224 3528
rect 5264 3408 5316 3460
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 10048 3680 10100 3732
rect 9680 3544 9732 3596
rect 9956 3476 10008 3528
rect 2320 3340 2372 3392
rect 3240 3340 3292 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 4436 3340 4488 3392
rect 9036 3340 9088 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 2044 3136 2096 3188
rect 2320 3136 2372 3188
rect 1860 3000 1912 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 3148 3136 3200 3188
rect 4068 3136 4120 3188
rect 10416 3136 10468 3188
rect 3148 3000 3200 3052
rect 3240 3000 3292 3052
rect 3792 3000 3844 3052
rect 3884 3000 3936 3052
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 5632 3000 5684 3052
rect 7472 3000 7524 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 2596 2796 2648 2848
rect 8944 2864 8996 2916
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 2504 2592 2556 2644
rect 2780 2592 2832 2644
rect 5540 2592 5592 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 7380 2592 7432 2644
rect 7748 2592 7800 2644
rect 8852 2592 8904 2644
rect 10048 2592 10100 2644
rect 940 2320 992 2372
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 2688 2456 2740 2508
rect 3240 2567 3292 2576
rect 3240 2533 3249 2567
rect 3249 2533 3283 2567
rect 3283 2533 3292 2567
rect 3240 2524 3292 2533
rect 4344 2524 4396 2576
rect 4436 2567 4488 2576
rect 4436 2533 4445 2567
rect 4445 2533 4479 2567
rect 4479 2533 4488 2567
rect 4436 2524 4488 2533
rect 2872 2388 2924 2440
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3148 2388 3200 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7748 2388 7800 2440
rect 10140 2524 10192 2576
rect 8944 2456 8996 2508
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 2964 2252 3016 2304
rect 3884 2320 3936 2372
rect 9404 2320 9456 2372
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 10508 2252 10560 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 572 2048 624 2100
rect 3792 2048 3844 2100
rect 2136 1980 2188 2032
rect 6828 1980 6880 2032
rect 1768 1368 1820 1420
rect 2504 1368 2556 1420
<< metal2 >>
rect 754 11200 810 12000
rect 2042 11200 2098 12000
rect 2778 11248 2834 11257
rect 768 8294 796 11200
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 940 9648 992 9654
rect 938 9616 940 9625
rect 992 9616 994 9625
rect 938 9551 994 9560
rect 1596 9178 1624 10231
rect 2056 9654 2084 11200
rect 3330 11200 3386 12000
rect 4618 11200 4674 12000
rect 5906 11200 5962 12000
rect 6012 11206 6224 11234
rect 2778 11183 2834 11192
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2792 9382 2820 11183
rect 3344 10010 3372 11200
rect 3252 9982 3372 10010
rect 3252 9654 3280 9982
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 4632 9654 4660 11200
rect 5920 11098 5948 11200
rect 6012 11098 6040 11206
rect 5920 11070 6040 11098
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6196 9722 6224 11206
rect 7194 11200 7250 12000
rect 8482 11200 8538 12000
rect 9770 11200 9826 12000
rect 11058 11200 11114 12000
rect 7208 9722 7236 11200
rect 8496 10282 8524 11200
rect 8496 10254 8708 10282
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8680 9722 8708 10254
rect 9784 9722 9812 11200
rect 10322 10704 10378 10713
rect 10322 10639 10378 10648
rect 10336 9722 10364 10639
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 10598 9616 10654 9625
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 9956 9580 10008 9586
rect 10598 9551 10654 9560
rect 9956 9522 10008 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1124 9036 1176 9042
rect 1124 8978 1176 8984
rect 1136 8809 1164 8978
rect 1122 8800 1178 8809
rect 1122 8735 1178 8744
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 756 8288 808 8294
rect 1504 8265 1532 8298
rect 756 8230 808 8236
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7177 980 7754
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 938 7168 994 7177
rect 938 7103 994 7112
rect 1504 7002 1532 7346
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 938 6352 994 6361
rect 1504 6338 1532 6938
rect 1688 6914 1716 9318
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1688 6886 1808 6914
rect 1504 6310 1716 6338
rect 938 6287 940 6296
rect 992 6287 994 6296
rect 940 6258 992 6264
rect 1688 5710 1716 6310
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1492 5636 1544 5642
rect 1492 5578 1544 5584
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4729 980 4966
rect 1504 4826 1532 5578
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1780 5522 1808 6886
rect 2056 6458 2084 8298
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 7546 2176 7754
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2516 6914 2544 9114
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8634 2728 8774
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2424 6886 2544 6914
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2424 6322 2452 6886
rect 2700 6458 2728 8434
rect 2884 8294 2912 9522
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 8498 3004 9454
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3068 8634 3096 8978
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 6866 2820 7822
rect 2884 7206 2912 8230
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 1964 5914 1992 6258
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5794 2084 6258
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 1582 5471 1638 5480
rect 1688 5494 1808 5522
rect 1964 5766 2084 5794
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1688 4622 1716 5494
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1780 4282 1808 5170
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 940 3936 992 3942
rect 938 3904 940 3913
rect 992 3904 994 3913
rect 938 3839 994 3848
rect 1780 3738 1808 4082
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1872 3534 1900 4966
rect 1964 3602 1992 5766
rect 2516 5370 2544 6258
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2608 5914 2636 6054
rect 2700 5914 2728 6054
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2516 4758 2544 4966
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 938 3088 994 3097
rect 1872 3058 1900 3470
rect 2056 3194 2084 4558
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2504 3936 2556 3942
rect 2608 3924 2636 4422
rect 2700 4146 2728 4422
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2608 3896 2820 3924
rect 2504 3878 2556 3884
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2516 3738 2544 3878
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3194 2360 3334
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 938 3023 994 3032
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2516 2650 2544 2994
rect 2608 2854 2636 3674
rect 2596 2848 2648 2854
rect 2792 2802 2820 3896
rect 2884 3738 2912 4490
rect 2976 4010 3004 8434
rect 3160 8362 3188 9522
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3344 8820 3372 9318
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3896 8974 3924 9454
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4264 9178 4292 9318
rect 4356 9178 4384 9522
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3344 8792 3832 8820
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3804 8106 3832 8792
rect 3896 8634 3924 8910
rect 4172 8838 4200 9046
rect 4540 9042 4568 9318
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 5000 9178 5028 9318
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 3804 8078 3924 8106
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7546 3280 7822
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3804 7546 3832 7890
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6118 3096 7278
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3252 6440 3280 6734
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3252 6412 3372 6440
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 4690 3096 6054
rect 3160 5574 3188 6190
rect 3252 5914 3280 6190
rect 3344 6118 3372 6412
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3344 5710 3372 6054
rect 3804 5914 3832 6734
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3332 5704 3384 5710
rect 3252 5652 3332 5658
rect 3252 5646 3384 5652
rect 3252 5630 3372 5646
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2964 3664 3016 3670
rect 2596 2790 2648 2796
rect 2700 2774 2820 2802
rect 2884 3612 2964 3618
rect 2884 3606 3016 3612
rect 2884 3590 3004 3606
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2700 2514 2728 2774
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2281 980 2314
rect 2136 2304 2188 2310
rect 938 2272 994 2281
rect 2136 2246 2188 2252
rect 938 2207 994 2216
rect 572 2100 624 2106
rect 572 2042 624 2048
rect 584 800 612 2042
rect 2148 2038 2176 2246
rect 2136 2032 2188 2038
rect 2136 1974 2188 1980
rect 2516 1426 2544 2382
rect 2792 1465 2820 2586
rect 2884 2446 2912 3590
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2976 2310 3004 3402
rect 3160 3194 3188 5510
rect 3252 5302 3280 5630
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3896 5012 3924 8078
rect 3988 7342 4016 8434
rect 4356 8090 4384 8434
rect 4620 8424 4672 8430
rect 4540 8372 4620 8378
rect 4540 8366 4672 8372
rect 4540 8350 4660 8366
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4080 6458 4108 6666
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3896 4984 4016 5012
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3252 4282 3280 4558
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3804 4282 3832 4422
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3738 3372 3878
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3896 3534 3924 4558
rect 3884 3528 3936 3534
rect 3804 3476 3884 3482
rect 3804 3470 3936 3476
rect 3804 3454 3924 3470
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3252 3058 3280 3334
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3804 3058 3832 3454
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3988 3058 4016 4984
rect 4356 4826 4384 7142
rect 4540 6934 4568 8350
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 5000 8090 5028 8978
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 7546 5028 8026
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4540 6390 4568 6870
rect 5000 6866 5028 7278
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6458 4844 6666
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5166 4476 5510
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4540 5030 4568 6326
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 6202 4936 6258
rect 4908 6174 5028 6202
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5000 5914 5028 6174
rect 5092 6118 5120 9114
rect 5460 8974 5488 9454
rect 5920 9110 5948 9454
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8566 5488 8774
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 7546 5396 7822
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7546 5488 7686
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 6196 7410 6224 9318
rect 6748 9178 6776 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7392 9110 7420 9522
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6380 8634 6408 8842
rect 7392 8634 7420 9046
rect 7484 9042 7512 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 7886 6408 8366
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7576 8090 7604 8910
rect 7668 8498 7696 9318
rect 7760 9178 7788 9522
rect 7852 9178 7880 9522
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7760 9058 7788 9114
rect 7760 9042 7880 9058
rect 7760 9036 7892 9042
rect 7760 9030 7840 9036
rect 7840 8978 7892 8984
rect 7944 8498 7972 9454
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5184 5794 5212 7346
rect 6472 7342 6500 7822
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7410 6592 7686
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6748 7274 6776 7822
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 5914 5396 6190
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5914 5488 6054
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5184 5766 5304 5794
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4540 4690 4568 4966
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4540 4214 4568 4626
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 5000 3738 5028 4490
rect 5092 4282 5120 4558
rect 5184 4282 5212 4966
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4080 3194 4108 3606
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3160 2446 3188 2994
rect 3252 2582 3280 2994
rect 3988 2774 4016 2994
rect 3896 2746 4016 2774
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2778 1456 2834 1465
rect 1768 1420 1820 1426
rect 1768 1362 1820 1368
rect 2504 1420 2556 1426
rect 2778 1391 2834 1400
rect 2504 1362 2556 1368
rect 1780 800 1808 1362
rect 3068 1306 3096 2382
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3804 2106 3832 2382
rect 3896 2378 3924 2746
rect 4356 2582 4384 3538
rect 5184 3534 5212 4218
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5276 3466 5304 5766
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5460 3738 5488 4150
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 2582 4476 3334
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 5552 2650 5580 6666
rect 5644 5914 5672 6734
rect 5736 6322 5764 6870
rect 5828 6866 5856 7142
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5710 5764 6054
rect 6380 5914 6408 6190
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 4826 5764 5646
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6656 5234 6684 7142
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7392 6798 7420 7822
rect 8036 7478 8064 9318
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 9968 9178 9996 9522
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10428 9081 10456 9114
rect 10414 9072 10470 9081
rect 10414 9007 10470 9016
rect 10612 8974 10640 9551
rect 11072 9110 11100 11200
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 9508 8430 9536 8842
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9692 8566 9720 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9784 8498 9812 8774
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9496 8424 9548 8430
rect 9416 8372 9496 8378
rect 9416 8366 9548 8372
rect 9416 8350 9536 8366
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8588 7886 8616 8230
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8680 7478 8708 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8772 7410 8800 7686
rect 9048 7546 9076 7822
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7546 9168 7686
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7576 7002 7604 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 5370 6868 6598
rect 7392 6458 7420 6734
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 6196 3942 6224 5034
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7392 4690 7420 5646
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 4146 6592 4422
rect 6656 4154 6684 4558
rect 6552 4140 6604 4146
rect 6656 4126 6776 4154
rect 6552 4082 6604 4088
rect 6748 4049 6776 4126
rect 6734 4040 6790 4049
rect 6734 3975 6790 3984
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5644 2650 5672 2994
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4252 2440 4304 2446
rect 4172 2400 4252 2428
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 2976 1278 3096 1306
rect 2976 800 3004 1278
rect 4172 800 4200 2400
rect 5448 2440 5500 2446
rect 4252 2382 4304 2388
rect 5368 2400 5448 2428
rect 5368 800 5396 2400
rect 6644 2440 6696 2446
rect 5448 2382 5500 2388
rect 6564 2400 6644 2428
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6564 800 6592 2400
rect 6644 2382 6696 2388
rect 6840 2038 6868 4558
rect 7024 4282 7052 4558
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 6932 3738 6960 4014
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7392 2650 7420 4014
rect 7484 3058 7512 6258
rect 7576 6202 7604 6938
rect 8312 6798 8340 7142
rect 8956 6914 8984 7278
rect 9140 7002 9168 7482
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8864 6886 8984 6914
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 6202 7696 6258
rect 7576 6174 7696 6202
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7576 5166 7604 5510
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7576 4282 7604 4626
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7668 4146 7696 4422
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7760 2650 7788 5510
rect 7944 4622 7972 6598
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8680 6254 8708 6598
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 5846 8524 6054
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8036 4282 8064 5578
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 4690 8156 5510
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8680 4690 8708 5714
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8864 2650 8892 6886
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9036 6656 9088 6662
rect 8956 6616 9036 6644
rect 8956 6322 8984 6616
rect 9036 6598 9088 6604
rect 9324 6458 9352 6734
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5658 8984 6258
rect 8956 5642 9076 5658
rect 8956 5636 9088 5642
rect 8956 5630 9036 5636
rect 8956 5098 8984 5630
rect 9036 5578 9088 5584
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 9140 4826 9168 5578
rect 9416 5234 9444 8350
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9876 8090 9904 8230
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7410 9996 7686
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 10152 7002 10180 8434
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10244 6914 10272 8910
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10508 8288 10560 8294
rect 10506 8256 10508 8265
rect 10560 8256 10562 8265
rect 10506 8191 10562 8200
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7449 10456 7686
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10414 7440 10470 7449
rect 10414 7375 10470 7384
rect 10876 6928 10928 6934
rect 10244 6886 10364 6914
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9876 6458 9904 6598
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9876 5642 9904 6394
rect 9968 5778 9996 6598
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5914 10088 6258
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8942 4040 8998 4049
rect 8942 3975 8944 3984
rect 8996 3975 8998 3984
rect 8944 3946 8996 3952
rect 9048 3738 9076 4694
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9232 3534 9260 5102
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9678 3632 9734 3641
rect 9678 3567 9680 3576
rect 9732 3567 9734 3576
rect 9680 3538 9732 3544
rect 9968 3534 9996 5578
rect 10244 5352 10272 6734
rect 10336 5658 10364 6886
rect 10876 6870 10928 6876
rect 10888 6769 10916 6870
rect 10874 6760 10930 6769
rect 10874 6695 10930 6704
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5817 10456 6054
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10336 5630 10456 5658
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10152 5324 10272 5352
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4622 10088 4966
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3738 10088 4082
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3058 9076 3334
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8956 2514 8984 2858
rect 9220 2848 9272 2854
rect 9272 2796 9444 2802
rect 9220 2790 9444 2796
rect 9232 2774 9444 2790
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 7760 800 7788 2382
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 9048 1306 9076 2382
rect 9416 2378 9444 2774
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 10152 2666 10180 5324
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 4622 10272 5170
rect 10336 5001 10364 5510
rect 10322 4992 10378 5001
rect 10322 4927 10378 4936
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4146 10272 4558
rect 10428 4282 10456 5630
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10414 4176 10470 4185
rect 10232 4140 10284 4146
rect 10414 4111 10470 4120
rect 10232 4082 10284 4088
rect 10428 3194 10456 4111
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10232 2848 10284 2854
rect 10284 2796 10364 2802
rect 10232 2790 10364 2796
rect 10244 2774 10364 2790
rect 10060 2650 10180 2666
rect 10048 2644 10180 2650
rect 10100 2638 10180 2644
rect 10048 2586 10100 2592
rect 10140 2576 10192 2582
rect 10336 2553 10364 2774
rect 10140 2518 10192 2524
rect 10322 2544 10378 2553
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9876 1737 9904 2246
rect 9862 1728 9918 1737
rect 9862 1663 9918 1672
rect 8956 1278 9076 1306
rect 8956 800 8984 1278
rect 10152 800 10180 2518
rect 10322 2479 10378 2488
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 921 10548 2246
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 10506 912 10562 921
rect 10506 847 10562 856
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
<< via2 >>
rect 1582 10240 1638 10296
rect 938 9596 940 9616
rect 940 9596 992 9616
rect 992 9596 994 9616
rect 938 9560 994 9596
rect 2778 11192 2834 11248
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 10322 10648 10378 10704
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10598 9560 10654 9616
rect 1122 8744 1178 8800
rect 1490 8200 1546 8256
rect 938 7112 994 7168
rect 938 6316 994 6352
rect 938 6296 940 6316
rect 940 6296 992 6316
rect 992 6296 994 6316
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 1582 5480 1638 5516
rect 938 4664 994 4720
rect 938 3884 940 3904
rect 940 3884 992 3904
rect 992 3884 994 3904
rect 938 3848 994 3884
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 938 3032 994 3088
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 938 2216 994 2272
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 2778 1400 2834 1456
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10414 9016 10470 9072
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 6734 3984 6790 4040
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10506 8236 10508 8256
rect 10508 8236 10560 8256
rect 10560 8236 10562 8256
rect 10506 8200 10562 8236
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10414 7384 10470 7440
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 8942 4004 8998 4040
rect 8942 3984 8944 4004
rect 8944 3984 8996 4004
rect 8996 3984 8998 4004
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9678 3596 9734 3632
rect 9678 3576 9680 3596
rect 9680 3576 9732 3596
rect 9732 3576 9734 3596
rect 10874 6704 10930 6760
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10414 5752 10470 5808
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 10322 4936 10378 4992
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10414 4120 10470 4176
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 9862 1672 9918 1728
rect 10322 2488 10378 2544
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 10506 856 10562 912
<< metal3 >>
rect 0 11250 800 11280
rect 2773 11250 2839 11253
rect 0 11248 2839 11250
rect 0 11192 2778 11248
rect 2834 11192 2839 11248
rect 0 11190 2839 11192
rect 0 11160 800 11190
rect 2773 11187 2839 11190
rect 10317 10706 10383 10709
rect 11200 10706 12000 10736
rect 10317 10704 12000 10706
rect 10317 10648 10322 10704
rect 10378 10648 12000 10704
rect 10317 10646 12000 10648
rect 10317 10643 10383 10646
rect 11200 10616 12000 10646
rect 0 10434 800 10464
rect 0 10374 1778 10434
rect 0 10344 800 10374
rect 1577 10298 1643 10301
rect 1718 10298 1778 10374
rect 1577 10296 1778 10298
rect 1577 10240 1582 10296
rect 1638 10240 1778 10296
rect 1577 10238 1778 10240
rect 1577 10235 1643 10238
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 11200 9800 12000 9920
rect 10698 9759 11014 9760
rect 11470 9690 11530 9800
rect 0 9618 800 9648
rect 11102 9630 11530 9690
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 10593 9618 10659 9621
rect 11102 9618 11162 9630
rect 10593 9616 11162 9618
rect 10593 9560 10598 9616
rect 10654 9560 11162 9616
rect 10593 9558 11162 9560
rect 10593 9555 10659 9558
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 10409 9074 10475 9077
rect 11200 9074 12000 9104
rect 10409 9072 12000 9074
rect 10409 9016 10414 9072
rect 10470 9016 12000 9072
rect 10409 9014 12000 9016
rect 10409 9011 10475 9014
rect 11200 8984 12000 9014
rect 0 8802 800 8832
rect 1117 8802 1183 8805
rect 0 8800 1183 8802
rect 0 8744 1122 8800
rect 1178 8744 1183 8800
rect 0 8742 1183 8744
rect 0 8712 800 8742
rect 1117 8739 1183 8742
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 1485 8258 1551 8261
rect 798 8256 1551 8258
rect 798 8200 1490 8256
rect 1546 8200 1551 8256
rect 798 8198 1551 8200
rect 798 8016 858 8198
rect 1485 8195 1551 8198
rect 10501 8258 10567 8261
rect 11200 8258 12000 8288
rect 10501 8256 12000 8258
rect 10501 8200 10506 8256
rect 10562 8200 12000 8256
rect 10501 8198 12000 8200
rect 10501 8195 10567 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 11200 8168 12000 8198
rect 9479 8127 9795 8128
rect 0 7926 858 8016
rect 0 7896 800 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 10409 7442 10475 7445
rect 11200 7442 12000 7472
rect 10409 7440 12000 7442
rect 10409 7384 10414 7440
rect 10470 7384 12000 7440
rect 10409 7382 12000 7384
rect 10409 7379 10475 7382
rect 11200 7352 12000 7382
rect 0 7170 800 7200
rect 933 7170 999 7173
rect 0 7168 999 7170
rect 0 7112 938 7168
rect 994 7112 999 7168
rect 0 7110 999 7112
rect 0 7080 800 7110
rect 933 7107 999 7110
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 10869 6762 10935 6765
rect 10869 6760 11162 6762
rect 10869 6704 10874 6760
rect 10930 6704 11162 6760
rect 10869 6702 11162 6704
rect 10869 6699 10935 6702
rect 11102 6660 11162 6702
rect 11102 6656 11346 6660
rect 11102 6600 12000 6656
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 11200 6536 12000 6600
rect 10698 6495 11014 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 10409 5810 10475 5813
rect 11200 5810 12000 5840
rect 10409 5808 12000 5810
rect 10409 5752 10414 5808
rect 10470 5752 12000 5808
rect 10409 5750 12000 5752
rect 10409 5747 10475 5750
rect 11200 5720 12000 5750
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 10317 4994 10383 4997
rect 11200 4994 12000 5024
rect 10317 4992 12000 4994
rect 10317 4936 10322 4992
rect 10378 4936 12000 4992
rect 10317 4934 12000 4936
rect 10317 4931 10383 4934
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 11200 4904 12000 4934
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 10409 4178 10475 4181
rect 11200 4178 12000 4208
rect 10409 4176 12000 4178
rect 10409 4120 10414 4176
rect 10470 4120 12000 4176
rect 10409 4118 12000 4120
rect 10409 4115 10475 4118
rect 11200 4088 12000 4118
rect 6729 4042 6795 4045
rect 8937 4042 9003 4045
rect 6729 4040 9003 4042
rect 6729 3984 6734 4040
rect 6790 3984 8942 4040
rect 8998 3984 9003 4040
rect 6729 3982 9003 3984
rect 6729 3979 6795 3982
rect 8937 3979 9003 3982
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 9673 3634 9739 3637
rect 9673 3632 11346 3634
rect 9673 3576 9678 3632
rect 9734 3576 11346 3632
rect 9673 3574 11346 3576
rect 9673 3571 9739 3574
rect 11286 3392 11346 3574
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 11200 3272 12000 3392
rect 10698 3231 11014 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 10317 2546 10383 2549
rect 11200 2546 12000 2576
rect 10317 2544 12000 2546
rect 10317 2488 10322 2544
rect 10378 2488 12000 2544
rect 10317 2486 12000 2488
rect 10317 2483 10383 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 933 2274 999 2277
rect 0 2272 999 2274
rect 0 2216 938 2272
rect 994 2216 999 2272
rect 0 2214 999 2216
rect 0 2184 800 2214
rect 933 2211 999 2214
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 9857 1730 9923 1733
rect 11200 1730 12000 1760
rect 9857 1728 12000 1730
rect 9857 1672 9862 1728
rect 9918 1672 12000 1728
rect 9857 1670 12000 1672
rect 9857 1667 9923 1670
rect 11200 1640 12000 1670
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 10501 914 10567 917
rect 11200 914 12000 944
rect 10501 912 12000 914
rect 10501 856 10506 912
rect 10562 856 12000 912
rect 10501 854 12000 856
rect 10501 851 10567 854
rect 11200 824 12000 854
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 7636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1688980957
transform 1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1688980957
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform -1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1688980957
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform -1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform -1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1688980957
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform -1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1688980957
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform -1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1688980957
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1688980957
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1688980957
transform -1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform -1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform -1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform -1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform -1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1688980957
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1688980957
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1688980957
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1688980957
transform -1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1688980957
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1688980957
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1688980957
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1688980957
transform -1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1688980957
transform -1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130_
timestamp 1688980957
transform -1 0 7268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1688980957
transform -1 0 7636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _132_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10396 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _133_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9568 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 1688980957
transform -1 0 2852 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 1688980957
transform -1 0 5060 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _137_
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 1688980957
transform -1 0 10396 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 1688980957
transform -1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp 1688980957
transform 1 0 2024 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _143_
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1688980957
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform -1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform -1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform -1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform -1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform -1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _167__44 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _167_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _168_
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _169_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _170_
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _171_
timestamp 1688980957
transform -1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _172_
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _173_
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _174_
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _175_
timestamp 1688980957
transform -1 0 9936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _176_
timestamp 1688980957
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _177_
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _178_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _179_
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _180__45
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _180_
timestamp 1688980957
transform -1 0 4784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _181_
timestamp 1688980957
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _182_
timestamp 1688980957
transform -1 0 5520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _183_
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _184_
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _185_
timestamp 1688980957
transform -1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _186_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _187_
timestamp 1688980957
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _188_
timestamp 1688980957
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _189_
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _190_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _191__46
timestamp 1688980957
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _191_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _192_
timestamp 1688980957
transform 1 0 2668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _193_
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _194_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _195__47
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _195_
timestamp 1688980957
transform -1 0 5704 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _196_
timestamp 1688980957
transform 1 0 3956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _197_
timestamp 1688980957
transform -1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _198_
timestamp 1688980957
transform -1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _199__48
timestamp 1688980957
transform 1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _199_
timestamp 1688980957
transform -1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _200_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _201_
timestamp 1688980957
transform 1 0 7544 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _202_
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_32
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_80
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_92
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_6
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_13
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_44
timestamp 1688980957
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_32
timestamp 1688980957
transform 1 0 4048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_38
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_68
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_80
timestamp 1688980957
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_12
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_28
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_76
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_36
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_101
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_12
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_24
timestamp 1688980957
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_32
timestamp 1688980957
transform 1 0 4048 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_49
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_57
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_64
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_74
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_26
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_43
timestamp 1688980957
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_87
timestamp 1688980957
transform 1 0 9108 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_79
timestamp 1688980957
transform 1 0 8372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_82
timestamp 1688980957
transform 1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_47
timestamp 1688980957
transform 1 0 5428 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_76
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_80
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_98
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_19
timestamp 1688980957
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_95
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp 1688980957
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_48
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1688980957
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_77
timestamp 1688980957
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_91
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 6716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 10212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 2668 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1688980957
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 2116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 2852 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1688980957
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal3 s 11200 9800 12000 9920 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 11200 10616 12000 10736 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 3 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 4 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 5 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 6 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 7 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 8 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 9 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 10 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 11 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 12 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 13 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 14 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 15 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 16 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 17 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 18 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 19 nsew signal tristate
flabel metal2 s 754 11200 810 12000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 20 nsew signal input
flabel metal2 s 2042 11200 2098 12000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 21 nsew signal input
flabel metal2 s 3330 11200 3386 12000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 22 nsew signal input
flabel metal2 s 4618 11200 4674 12000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 23 nsew signal input
flabel metal2 s 5906 11200 5962 12000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 24 nsew signal input
flabel metal2 s 7194 11200 7250 12000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 25 nsew signal input
flabel metal2 s 8482 11200 8538 12000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 26 nsew signal input
flabel metal2 s 9770 11200 9826 12000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 27 nsew signal input
flabel metal2 s 11058 11200 11114 12000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 28 nsew signal input
flabel metal3 s 11200 824 12000 944 0 FreeSans 480 0 0 0 chany_top_out[0]
port 29 nsew signal tristate
flabel metal3 s 11200 1640 12000 1760 0 FreeSans 480 0 0 0 chany_top_out[1]
port 30 nsew signal tristate
flabel metal3 s 11200 2456 12000 2576 0 FreeSans 480 0 0 0 chany_top_out[2]
port 31 nsew signal tristate
flabel metal3 s 11200 3272 12000 3392 0 FreeSans 480 0 0 0 chany_top_out[3]
port 32 nsew signal tristate
flabel metal3 s 11200 4088 12000 4208 0 FreeSans 480 0 0 0 chany_top_out[4]
port 33 nsew signal tristate
flabel metal3 s 11200 4904 12000 5024 0 FreeSans 480 0 0 0 chany_top_out[5]
port 34 nsew signal tristate
flabel metal3 s 11200 5720 12000 5840 0 FreeSans 480 0 0 0 chany_top_out[6]
port 35 nsew signal tristate
flabel metal3 s 11200 6536 12000 6656 0 FreeSans 480 0 0 0 chany_top_out[7]
port 36 nsew signal tristate
flabel metal3 s 11200 7352 12000 7472 0 FreeSans 480 0 0 0 chany_top_out[8]
port 37 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 38 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 39 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 40 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 41 nsew signal input
flabel metal3 s 11200 8168 12000 8288 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 42 nsew signal tristate
flabel metal3 s 11200 8984 12000 9104 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 43 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 3634 4182 3634 4182 0 _000_
rlabel metal1 4876 5202 4876 5202 0 _001_
rlabel metal1 2070 3060 2070 3060 0 _002_
rlabel metal1 2346 5644 2346 5644 0 _003_
rlabel metal2 2530 5814 2530 5814 0 _004_
rlabel metal1 2070 5882 2070 5882 0 _005_
rlabel metal1 6302 5712 6302 5712 0 _006_
rlabel metal1 3726 5882 3726 5882 0 _007_
rlabel metal1 8372 6290 8372 6290 0 _008_
rlabel metal1 8418 7310 8418 7310 0 _009_
rlabel metal2 9246 4318 9246 4318 0 _010_
rlabel metal1 8832 7378 8832 7378 0 _011_
rlabel metal1 6808 4114 6808 4114 0 _012_
rlabel metal1 8970 6698 8970 6698 0 _013_
rlabel metal1 6486 7378 6486 7378 0 _014_
rlabel metal1 8096 9146 8096 9146 0 _015_
rlabel metal1 3174 7344 3174 7344 0 _016_
rlabel metal1 3634 8942 3634 8942 0 _017_
rlabel metal1 8740 6630 8740 6630 0 _018_
rlabel metal2 7038 4420 7038 4420 0 _019_
rlabel metal1 9706 3366 9706 3366 0 _020_
rlabel metal1 7130 7276 7130 7276 0 _021_
rlabel metal2 9062 7684 9062 7684 0 _022_
rlabel metal1 8050 6188 8050 6188 0 _023_
rlabel metal1 7498 4114 7498 4114 0 _024_
rlabel metal1 7912 6766 7912 6766 0 _025_
rlabel metal1 9706 7276 9706 7276 0 _026_
rlabel metal1 8096 4658 8096 4658 0 _027_
rlabel metal1 9154 6426 9154 6426 0 _028_
rlabel metal1 8924 4794 8924 4794 0 _029_
rlabel metal1 2116 6426 2116 6426 0 _030_
rlabel metal1 4002 6698 4002 6698 0 _031_
rlabel metal1 2530 5746 2530 5746 0 _032_
rlabel metal1 5888 5814 5888 5814 0 _033_
rlabel metal1 2714 5814 2714 5814 0 _034_
rlabel metal1 2162 3162 2162 3162 0 _035_
rlabel metal1 2622 7276 2622 7276 0 _036_
rlabel metal1 5060 5814 5060 5814 0 _037_
rlabel metal1 2530 4692 2530 4692 0 _038_
rlabel metal1 6164 5882 6164 5882 0 _039_
rlabel metal1 2346 3128 2346 3128 0 _040_
rlabel metal1 2254 2822 2254 2822 0 _041_
rlabel metal1 5244 5270 5244 5270 0 _042_
rlabel metal1 3174 4046 3174 4046 0 _043_
rlabel metal1 5152 3638 5152 3638 0 _044_
rlabel metal1 2530 3638 2530 3638 0 _045_
rlabel metal1 3634 9044 3634 9044 0 _046_
rlabel metal1 3634 7208 3634 7208 0 _047_
rlabel metal2 4554 9180 4554 9180 0 _048_
rlabel metal1 3404 7514 3404 7514 0 _049_
rlabel metal1 7636 8466 7636 8466 0 _050_
rlabel metal1 6670 7242 6670 7242 0 _051_
rlabel metal1 7636 9010 7636 9010 0 _052_
rlabel metal1 6900 7922 6900 7922 0 _053_
rlabel metal1 9890 8908 9890 8908 0 ccff_head
rlabel metal1 10304 9690 10304 9690 0 ccff_tail
rlabel metal2 598 1418 598 1418 0 chany_bottom_in[0]
rlabel metal2 1794 1078 1794 1078 0 chany_bottom_in[1]
rlabel metal2 2990 1027 2990 1027 0 chany_bottom_in[2]
rlabel metal2 4186 1588 4186 1588 0 chany_bottom_in[3]
rlabel metal2 5382 1588 5382 1588 0 chany_bottom_in[4]
rlabel metal2 6578 1588 6578 1588 0 chany_bottom_in[5]
rlabel metal2 7774 1588 7774 1588 0 chany_bottom_in[6]
rlabel metal2 8970 1027 8970 1027 0 chany_bottom_in[7]
rlabel metal2 10166 1656 10166 1656 0 chany_bottom_in[8]
rlabel metal3 820 2244 820 2244 0 chany_bottom_out[0]
rlabel metal3 820 3060 820 3060 0 chany_bottom_out[1]
rlabel metal3 820 3876 820 3876 0 chany_bottom_out[2]
rlabel metal3 820 4692 820 4692 0 chany_bottom_out[3]
rlabel metal3 1142 5508 1142 5508 0 chany_bottom_out[4]
rlabel metal3 820 6324 820 6324 0 chany_bottom_out[5]
rlabel metal3 820 7140 820 7140 0 chany_bottom_out[6]
rlabel metal3 751 7956 751 7956 0 chany_bottom_out[7]
rlabel metal3 912 8772 912 8772 0 chany_bottom_out[8]
rlabel metal1 2622 8296 2622 8296 0 chany_top_in[0]
rlabel metal1 1794 9554 1794 9554 0 chany_top_in[1]
rlabel metal1 3450 9554 3450 9554 0 chany_top_in[2]
rlabel metal1 4922 9588 4922 9588 0 chany_top_in[3]
rlabel metal1 6210 9622 6210 9622 0 chany_top_in[4]
rlabel metal1 6946 9588 6946 9588 0 chany_top_in[5]
rlabel metal1 8740 9554 8740 9554 0 chany_top_in[6]
rlabel metal1 9798 9622 9798 9622 0 chany_top_in[7]
rlabel metal1 10166 8976 10166 8976 0 chany_top_in[8]
rlabel metal1 10488 2278 10488 2278 0 chany_top_out[0]
rlabel metal2 9890 1989 9890 1989 0 chany_top_out[1]
rlabel metal3 10818 2516 10818 2516 0 chany_top_out[2]
rlabel metal1 9706 3638 9706 3638 0 chany_top_out[3]
rlabel metal1 10074 3162 10074 3162 0 chany_top_out[4]
rlabel metal1 9522 5542 9522 5542 0 chany_top_out[5]
rlabel metal2 10442 5933 10442 5933 0 chany_top_out[6]
rlabel metal1 10672 6970 10672 6970 0 chany_top_out[7]
rlabel metal2 10442 7565 10442 7565 0 chany_top_out[8]
rlabel metal1 4370 5304 4370 5304 0 clknet_0_prog_clk
rlabel metal1 3818 4148 3818 4148 0 clknet_1_0__leaf_prog_clk
rlabel metal1 6394 5236 6394 5236 0 clknet_1_1__leaf_prog_clk
rlabel metal3 820 9588 820 9588 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal3 1211 10404 1211 10404 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal2 2806 10285 2806 10285 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal2 6578 4284 6578 4284 0 mem_left_ipin_0.DFF_0_.Q
rlabel metal1 8924 6290 8924 6290 0 mem_left_ipin_0.DFF_1_.Q
rlabel metal1 8510 4590 8510 4590 0 mem_left_ipin_0.DFF_2_.Q
rlabel metal1 2622 4080 2622 4080 0 mem_left_ipin_1.DFF_0_.Q
rlabel metal1 5152 3502 5152 3502 0 mem_left_ipin_1.DFF_1_.Q
rlabel metal1 1610 3026 1610 3026 0 mem_right_ipin_0.DFF_0_.Q
rlabel metal1 2254 5236 2254 5236 0 mem_right_ipin_0.DFF_1_.Q
rlabel metal2 1610 6324 1610 6324 0 mem_right_ipin_0.DFF_2_.Q
rlabel metal1 3818 7956 3818 7956 0 mem_right_ipin_1.DFF_0_.Q
rlabel metal1 3956 8942 3956 8942 0 mem_right_ipin_1.DFF_1_.Q
rlabel metal1 6118 8364 6118 8364 0 mem_right_ipin_2.DFF_0_.Q
rlabel metal1 7084 3706 7084 3706 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal2 2162 2142 2162 2142 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 7314 6426 7314 6426 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal1 6578 7854 6578 7854 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 9982 7310 9982 7310 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 9844 7922 9844 7922 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 7682 4658 7682 4658 0 mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7682 6970 7682 6970 0 mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9200 7514 9200 7514 0 mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 8786 5746 8786 5746 0 mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 9890 6528 9890 6528 0 mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 9936 5746 9936 5746 0 mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3312 2346 3312 2346 0 mux_left_ipin_1.INVTX1_0_.out
rlabel metal1 1978 4556 1978 4556 0 mux_left_ipin_1.INVTX1_1_.out
rlabel metal2 3358 3808 3358 3808 0 mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5934 3944 5934 3944 0 mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2852 3026 2852 3026 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal1 2622 5814 2622 5814 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal2 6946 6052 6946 6052 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal1 5658 6834 5658 6834 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 2990 4658 2990 4658 0 mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3220 5542 3220 5542 0 mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 5980 6290 5980 6290 0 mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 3082 5372 3082 5372 0 mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2438 8466 2438 8466 0 mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2898 8908 2898 8908 0 mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 5244 7514 5244 7514 0 mux_right_ipin_1.INVTX1_0_.out
rlabel metal2 4002 7888 4002 7888 0 mux_right_ipin_1.INVTX1_1_.out
rlabel metal2 5014 8534 5014 8534 0 mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4692 9146 4692 9146 0 mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7682 8058 7682 8058 0 mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7268 8602 7268 8602 0 mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9491 8534 9491 8534 0 net1
rlabel metal1 8832 2618 8832 2618 0 net10
rlabel metal1 2254 2346 2254 2346 0 net11
rlabel metal1 1702 4522 1702 4522 0 net12
rlabel metal1 2254 6290 2254 6290 0 net13
rlabel metal1 2162 4046 2162 4046 0 net14
rlabel metal1 1610 4692 1610 4692 0 net15
rlabel metal1 6026 9044 6026 9044 0 net16
rlabel metal1 5934 7412 5934 7412 0 net17
rlabel metal1 2990 8942 2990 8942 0 net18
rlabel metal1 3082 8568 3082 8568 0 net19
rlabel metal1 5842 3536 5842 3536 0 net2
rlabel metal1 8510 8976 8510 8976 0 net20
rlabel metal1 1794 2448 1794 2448 0 net21
rlabel metal1 2898 2278 2898 2278 0 net22
rlabel metal1 2116 3706 2116 3706 0 net23
rlabel metal1 1886 4250 1886 4250 0 net24
rlabel metal1 1472 4794 1472 4794 0 net25
rlabel metal1 1840 6290 1840 6290 0 net26
rlabel metal1 1794 7752 1794 7752 0 net27
rlabel metal1 2254 8534 2254 8534 0 net28
rlabel metal1 2990 8840 2990 8840 0 net29
rlabel metal1 2622 2618 2622 2618 0 net3
rlabel metal1 9798 2346 9798 2346 0 net30
rlabel metal1 2714 2856 2714 2856 0 net31
rlabel metal1 3726 3128 3726 3128 0 net32
rlabel metal1 5934 3604 5934 3604 0 net33
rlabel metal1 9200 3094 9200 3094 0 net34
rlabel metal2 8050 4930 8050 4930 0 net35
rlabel metal1 8970 5882 8970 5882 0 net36
rlabel metal1 9798 2618 9798 2618 0 net37
rlabel metal1 10166 7854 10166 7854 0 net38
rlabel metal1 2576 9622 2576 9622 0 net39
rlabel metal1 3404 3026 3404 3026 0 net4
rlabel metal1 2369 8942 2369 8942 0 net40
rlabel metal1 2622 9486 2622 9486 0 net41
rlabel metal1 10120 6970 10120 6970 0 net42
rlabel metal2 10258 7921 10258 7921 0 net43
rlabel metal1 9614 6290 9614 6290 0 net44
rlabel metal1 4876 6834 4876 6834 0 net45
rlabel metal1 5658 5134 5658 5134 0 net46
rlabel metal1 5704 9486 5704 9486 0 net47
rlabel metal1 7866 8466 7866 8466 0 net48
rlabel metal2 6394 8738 6394 8738 0 net49
rlabel metal1 5750 3468 5750 3468 0 net5
rlabel metal1 5239 8534 5239 8534 0 net50
rlabel metal1 4595 4114 4595 4114 0 net51
rlabel metal1 4416 8058 4416 8058 0 net52
rlabel metal1 4917 4522 4917 4522 0 net53
rlabel metal1 2116 7514 2116 7514 0 net54
rlabel metal1 10304 3706 10304 3706 0 net55
rlabel metal1 4968 5882 4968 5882 0 net56
rlabel via1 6665 5202 6665 5202 0 net57
rlabel metal1 2775 6698 2775 6698 0 net58
rlabel via1 10078 4590 10078 4590 0 net59
rlabel metal2 5658 2822 5658 2822 0 net6
rlabel metal1 7130 2618 7130 2618 0 net7
rlabel metal1 7820 2618 7820 2618 0 net8
rlabel metal1 9292 2414 9292 2414 0 net9
rlabel metal3 1740 1428 1740 1428 0 prog_clk
rlabel metal1 10488 8262 10488 8262 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel metal2 10442 9095 10442 9095 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
