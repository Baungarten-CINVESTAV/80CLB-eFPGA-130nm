* NGSPICE file created from grid_io_top_out.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt grid_io_top_out bottom_width_0_height_0_subtile_0__pin_inpad_0_ bottom_width_0_height_0_subtile_0__pin_outpad_0_
+ ccff_head ccff_tail gfpga_pad_GPIO_PAD prog_clk vdd vss
Xgrid_io_top_out_5 vss vss vdd vdd grid_io_top_out_5/HI bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_27 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_9_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_7_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_4_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput1 bottom_width_0_height_0_subtile_0__pin_outpad_0_ vss vss vdd vdd net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_29 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput2 ccff_head vss vss vdd vdd net2 sky130_fd_sc_hd__clkbuf_1
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_30 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_2_ net1 vss vss vdd vdd net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_0_ prog_clk net2 vss vss vdd vdd net3 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_29 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_8_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_25 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_24 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_26 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XTAP_27 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_28 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_29 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_21 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_23 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput3 net3 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_0_0_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput4 net4 vss vss vdd vdd gfpga_pad_GPIO_PAD sky130_fd_sc_hd__clkbuf_4
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_0_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_6_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
.ends

