magic
tech sky130A
magscale 1 2
timestamp 1712074353
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 750 2128 583450 701808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 754 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583444 703610
rect 754 536 583444 703464
rect 754 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
rect 165022 326 165994 536
rect 166218 326 167098 536
rect 167322 326 168294 536
rect 168518 326 169490 536
rect 169714 326 170686 536
rect 170910 326 171882 536
rect 172106 326 173078 536
rect 173302 326 174182 536
rect 174406 326 175378 536
rect 175602 326 176574 536
rect 176798 326 177770 536
rect 177994 326 178966 536
rect 179190 326 180162 536
rect 180386 326 181358 536
rect 181582 326 182462 536
rect 182686 326 183658 536
rect 183882 326 184854 536
rect 185078 326 186050 536
rect 186274 326 187246 536
rect 187470 326 188442 536
rect 188666 326 189638 536
rect 189862 326 190742 536
rect 190966 326 191938 536
rect 192162 326 193134 536
rect 193358 326 194330 536
rect 194554 326 195526 536
rect 195750 326 196722 536
rect 196946 326 197826 536
rect 198050 326 199022 536
rect 199246 326 200218 536
rect 200442 326 201414 536
rect 201638 326 202610 536
rect 202834 326 203806 536
rect 204030 326 205002 536
rect 205226 326 206106 536
rect 206330 326 207302 536
rect 207526 326 208498 536
rect 208722 326 209694 536
rect 209918 326 210890 536
rect 211114 326 212086 536
rect 212310 326 213282 536
rect 213506 326 214386 536
rect 214610 326 215582 536
rect 215806 326 216778 536
rect 217002 326 217974 536
rect 218198 326 219170 536
rect 219394 326 220366 536
rect 220590 326 221470 536
rect 221694 326 222666 536
rect 222890 326 223862 536
rect 224086 326 225058 536
rect 225282 326 226254 536
rect 226478 326 227450 536
rect 227674 326 228646 536
rect 228870 326 229750 536
rect 229974 326 230946 536
rect 231170 326 232142 536
rect 232366 326 233338 536
rect 233562 326 234534 536
rect 234758 326 235730 536
rect 235954 326 236926 536
rect 237150 326 238030 536
rect 238254 326 239226 536
rect 239450 326 240422 536
rect 240646 326 241618 536
rect 241842 326 242814 536
rect 243038 326 244010 536
rect 244234 326 245114 536
rect 245338 326 246310 536
rect 246534 326 247506 536
rect 247730 326 248702 536
rect 248926 326 249898 536
rect 250122 326 251094 536
rect 251318 326 252290 536
rect 252514 326 253394 536
rect 253618 326 254590 536
rect 254814 326 255786 536
rect 256010 326 256982 536
rect 257206 326 258178 536
rect 258402 326 259374 536
rect 259598 326 260570 536
rect 260794 326 261674 536
rect 261898 326 262870 536
rect 263094 326 264066 536
rect 264290 326 265262 536
rect 265486 326 266458 536
rect 266682 326 267654 536
rect 267878 326 268758 536
rect 268982 326 269954 536
rect 270178 326 271150 536
rect 271374 326 272346 536
rect 272570 326 273542 536
rect 273766 326 274738 536
rect 274962 326 275934 536
rect 276158 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280626 536
rect 280850 326 281822 536
rect 282046 326 283018 536
rect 283242 326 284214 536
rect 284438 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300682 536
rect 300906 326 301878 536
rect 302102 326 303074 536
rect 303298 326 304270 536
rect 304494 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 308962 536
rect 309186 326 310158 536
rect 310382 326 311354 536
rect 311578 326 312550 536
rect 312774 326 313746 536
rect 313970 326 314942 536
rect 315166 326 316138 536
rect 316362 326 317242 536
rect 317466 326 318438 536
rect 318662 326 319634 536
rect 319858 326 320830 536
rect 321054 326 322026 536
rect 322250 326 323222 536
rect 323446 326 324326 536
rect 324550 326 325522 536
rect 325746 326 326718 536
rect 326942 326 327914 536
rect 328138 326 329110 536
rect 329334 326 330306 536
rect 330530 326 331502 536
rect 331726 326 332606 536
rect 332830 326 333802 536
rect 334026 326 334998 536
rect 335222 326 336194 536
rect 336418 326 337390 536
rect 337614 326 338586 536
rect 338810 326 339782 536
rect 340006 326 340886 536
rect 341110 326 342082 536
rect 342306 326 343278 536
rect 343502 326 344474 536
rect 344698 326 345670 536
rect 345894 326 346866 536
rect 347090 326 347970 536
rect 348194 326 349166 536
rect 349390 326 350362 536
rect 350586 326 351558 536
rect 351782 326 352754 536
rect 352978 326 353950 536
rect 354174 326 355146 536
rect 355370 326 356250 536
rect 356474 326 357446 536
rect 357670 326 358642 536
rect 358866 326 359838 536
rect 360062 326 361034 536
rect 361258 326 362230 536
rect 362454 326 363426 536
rect 363650 326 364530 536
rect 364754 326 365726 536
rect 365950 326 366922 536
rect 367146 326 368118 536
rect 368342 326 369314 536
rect 369538 326 370510 536
rect 370734 326 371614 536
rect 371838 326 372810 536
rect 373034 326 374006 536
rect 374230 326 375202 536
rect 375426 326 376398 536
rect 376622 326 377594 536
rect 377818 326 378790 536
rect 379014 326 379894 536
rect 380118 326 381090 536
rect 381314 326 382286 536
rect 382510 326 383482 536
rect 383706 326 384678 536
rect 384902 326 385874 536
rect 386098 326 387070 536
rect 387294 326 388174 536
rect 388398 326 389370 536
rect 389594 326 390566 536
rect 390790 326 391762 536
rect 391986 326 392958 536
rect 393182 326 394154 536
rect 394378 326 395258 536
rect 395482 326 396454 536
rect 396678 326 397650 536
rect 397874 326 398846 536
rect 399070 326 400042 536
rect 400266 326 401238 536
rect 401462 326 402434 536
rect 402658 326 403538 536
rect 403762 326 404734 536
rect 404958 326 405930 536
rect 406154 326 407126 536
rect 407350 326 408322 536
rect 408546 326 409518 536
rect 409742 326 410714 536
rect 410938 326 411818 536
rect 412042 326 413014 536
rect 413238 326 414210 536
rect 414434 326 415406 536
rect 415630 326 416602 536
rect 416826 326 417798 536
rect 418022 326 418902 536
rect 419126 326 420098 536
rect 420322 326 421294 536
rect 421518 326 422490 536
rect 422714 326 423686 536
rect 423910 326 424882 536
rect 425106 326 426078 536
rect 426302 326 427182 536
rect 427406 326 428378 536
rect 428602 326 429574 536
rect 429798 326 430770 536
rect 430994 326 431966 536
rect 432190 326 433162 536
rect 433386 326 434358 536
rect 434582 326 435462 536
rect 435686 326 436658 536
rect 436882 326 437854 536
rect 438078 326 439050 536
rect 439274 326 440246 536
rect 440470 326 441442 536
rect 441666 326 442546 536
rect 442770 326 443742 536
rect 443966 326 444938 536
rect 445162 326 446134 536
rect 446358 326 447330 536
rect 447554 326 448526 536
rect 448750 326 449722 536
rect 449946 326 450826 536
rect 451050 326 452022 536
rect 452246 326 453218 536
rect 453442 326 454414 536
rect 454638 326 455610 536
rect 455834 326 456806 536
rect 457030 326 458002 536
rect 458226 326 459106 536
rect 459330 326 460302 536
rect 460526 326 461498 536
rect 461722 326 462694 536
rect 462918 326 463890 536
rect 464114 326 465086 536
rect 465310 326 466190 536
rect 466414 326 467386 536
rect 467610 326 468582 536
rect 468806 326 469778 536
rect 470002 326 470974 536
rect 471198 326 472170 536
rect 472394 326 473366 536
rect 473590 326 474470 536
rect 474694 326 475666 536
rect 475890 326 476862 536
rect 477086 326 478058 536
rect 478282 326 479254 536
rect 479478 326 480450 536
rect 480674 326 481646 536
rect 481870 326 482750 536
rect 482974 326 483946 536
rect 484170 326 485142 536
rect 485366 326 486338 536
rect 486562 326 487534 536
rect 487758 326 488730 536
rect 488954 326 489834 536
rect 490058 326 491030 536
rect 491254 326 492226 536
rect 492450 326 493422 536
rect 493646 326 494618 536
rect 494842 326 495814 536
rect 496038 326 497010 536
rect 497234 326 498114 536
rect 498338 326 499310 536
rect 499534 326 500506 536
rect 500730 326 501702 536
rect 501926 326 502898 536
rect 503122 326 504094 536
rect 504318 326 505290 536
rect 505514 326 506394 536
rect 506618 326 507590 536
rect 507814 326 508786 536
rect 509010 326 509982 536
rect 510206 326 511178 536
rect 511402 326 512374 536
rect 512598 326 513478 536
rect 513702 326 514674 536
rect 514898 326 515870 536
rect 516094 326 517066 536
rect 517290 326 518262 536
rect 518486 326 519458 536
rect 519682 326 520654 536
rect 520878 326 521758 536
rect 521982 326 522954 536
rect 523178 326 524150 536
rect 524374 326 525346 536
rect 525570 326 526542 536
rect 526766 326 527738 536
rect 527962 326 528934 536
rect 529158 326 530038 536
rect 530262 326 531234 536
rect 531458 326 532430 536
rect 532654 326 533626 536
rect 533850 326 534822 536
rect 535046 326 536018 536
rect 536242 326 537122 536
rect 537346 326 538318 536
rect 538542 326 539514 536
rect 539738 326 540710 536
rect 540934 326 541906 536
rect 542130 326 543102 536
rect 543326 326 544298 536
rect 544522 326 545402 536
rect 545626 326 546598 536
rect 546822 326 547794 536
rect 548018 326 548990 536
rect 549214 326 550186 536
rect 550410 326 551382 536
rect 551606 326 552578 536
rect 552802 326 553682 536
rect 553906 326 554878 536
rect 555102 326 556074 536
rect 556298 326 557270 536
rect 557494 326 558466 536
rect 558690 326 559662 536
rect 559886 326 560766 536
rect 560990 326 561962 536
rect 562186 326 563158 536
rect 563382 326 564354 536
rect 564578 326 565550 536
rect 565774 326 566746 536
rect 566970 326 567942 536
rect 568166 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572634 536
rect 572858 326 573830 536
rect 574054 326 575026 536
rect 575250 326 576222 536
rect 576446 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580914 536
rect 581138 326 582110 536
rect 582334 326 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583520 701793
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 2143 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 994 -7654 1614 711590
rect 4714 -7654 5334 711590
rect 36994 676580 37614 711590
rect 21310 662000 21930 672432
rect 22046 662000 22666 672432
rect 36994 613780 37614 664588
rect 21310 598896 21930 609872
rect 22046 598896 22666 609872
rect 36994 585764 37614 601788
rect 40714 585764 41334 711590
rect 53694 662544 54314 678960
rect 72994 675793 73614 711590
rect 76714 675793 77334 711590
rect 108994 676580 109614 711590
rect 112714 676580 113334 711590
rect 148714 685532 149334 711590
rect 53694 599440 54314 615856
rect 72994 612993 73614 655399
rect 76714 612993 77334 655399
rect 93254 632624 93874 650672
rect 97118 632624 97738 650672
rect 108994 650196 109614 664588
rect 112714 650196 113334 664588
rect 122510 662000 123130 679504
rect 126374 662000 126994 679504
rect 127294 632624 127914 650672
rect 131158 632624 131778 650672
rect 144994 647580 145614 655399
rect 148714 647580 149334 655399
rect 108994 613780 109614 629175
rect 112714 613780 113334 629175
rect 144994 622732 145614 635588
rect 148714 622732 149334 635588
rect 157286 632624 157906 650672
rect 161150 632624 161770 650672
rect 122326 614672 122946 616944
rect 126190 614672 126810 616944
rect 36994 550980 37614 567788
rect 21310 536336 21930 546768
rect 22046 536336 22666 546768
rect 36994 522964 37614 538988
rect 40714 522964 41334 567788
rect 53694 536336 54314 553840
rect 72994 550193 73614 592599
rect 76714 550193 77334 592599
rect 108994 591748 109614 601788
rect 112714 591748 113334 601788
rect 122510 598896 123130 614592
rect 126374 598896 126994 614592
rect 122878 591280 123498 594640
rect 126742 592000 127362 594640
rect 126926 589648 127546 591920
rect 130790 589648 131410 591920
rect 93254 568976 93874 586480
rect 97118 568976 97738 586480
rect 127294 570784 127914 586480
rect 131158 570784 131778 586480
rect 144994 583580 145614 592599
rect 148714 583580 149334 592599
rect 126926 568432 127546 570704
rect 130790 568432 131410 570704
rect 108994 550980 109614 567463
rect 112714 550980 113334 567463
rect 144994 559932 145614 569767
rect 148714 559932 149334 571588
rect 157286 570704 157906 586480
rect 158758 568976 159378 571792
rect 159494 568976 160114 571792
rect 161150 570704 161770 586480
rect 36994 488180 37614 504988
rect 21310 473232 21930 484208
rect 22046 473232 22666 484208
rect 36994 460164 37614 476188
rect 40714 460164 41334 504988
rect 53694 473232 54314 490736
rect 72994 487393 73614 529799
rect 76714 487393 77334 529799
rect 108994 528948 109614 538988
rect 112714 528948 113334 538988
rect 122510 536336 123130 553840
rect 126374 536336 126994 553840
rect 122878 527088 123498 532080
rect 126742 527088 127362 532080
rect 93254 506960 93874 525008
rect 97118 506960 97738 525008
rect 127294 506960 127914 525008
rect 131158 506960 131778 525008
rect 144994 521980 145614 529799
rect 148714 521980 149334 529799
rect 108994 488180 109614 504663
rect 112714 488180 113334 504663
rect 144994 497132 145614 508167
rect 148714 497132 149334 509988
rect 157286 506960 157906 525008
rect 161150 506960 161770 525008
rect 36994 425380 37614 442188
rect 21310 410672 21930 421104
rect 22046 410672 22666 421104
rect 36994 397364 37614 413388
rect 40714 397364 41334 442188
rect 53694 411216 54314 427632
rect 72994 424593 73614 466999
rect 76714 424593 77334 466999
rect 108994 466148 109614 476188
rect 112714 466148 113334 476188
rect 122510 473232 123130 491280
rect 126374 473232 126994 491280
rect 122878 464528 123498 468976
rect 126742 464528 127362 468976
rect 93254 444400 93874 461904
rect 97118 444400 97738 461904
rect 127294 444400 127914 461904
rect 131158 444400 131778 461904
rect 144994 459180 145614 466999
rect 148714 459180 149334 466999
rect 108994 425380 109614 441863
rect 112714 425380 113334 441926
rect 144994 434332 145614 445367
rect 148714 434332 149334 447188
rect 157286 444400 157906 461904
rect 161150 444400 161770 461904
rect 60318 384560 60938 396624
rect 36994 362580 37614 379388
rect 21310 347568 21930 358544
rect 22046 347568 22666 358544
rect 36994 334564 37614 350588
rect 40714 334564 41334 379388
rect 53694 348112 54314 365616
rect 72994 361793 73614 404199
rect 76714 361793 77334 404199
rect 108994 403348 109614 413388
rect 112714 403348 113334 413388
rect 122510 410672 123130 428176
rect 126374 410672 126994 428176
rect 122878 401424 123498 406416
rect 126742 401424 127362 406416
rect 93254 381296 93874 399344
rect 97118 381296 97738 399344
rect 127294 381296 127914 399344
rect 131158 381296 131778 399344
rect 144994 396380 145614 404199
rect 148714 396380 149334 404199
rect 108994 362580 109614 379063
rect 112714 362580 113334 379063
rect 144994 371532 145614 382567
rect 148714 371532 149334 384388
rect 157286 381296 157906 399344
rect 161150 381296 161770 399344
rect 36994 299780 37614 316588
rect 21310 285008 21930 295440
rect 22046 285008 22666 295440
rect 36994 271764 37614 287788
rect 40714 271764 41334 316588
rect 53694 285008 54314 302512
rect 72994 298993 73614 341399
rect 76714 298993 77334 341399
rect 108994 340548 109614 350588
rect 112714 340548 113334 350588
rect 122510 347568 123130 365616
rect 126374 347568 126994 365616
rect 122878 338864 123498 343312
rect 126742 338864 127362 343312
rect 93254 318736 93874 336240
rect 97118 318736 97738 336240
rect 121406 334512 122026 336784
rect 125270 334512 125890 336784
rect 127294 318736 127914 334512
rect 131158 318736 131778 334512
rect 144994 333580 145614 341399
rect 148714 333580 149334 341399
rect 108994 299780 109614 316263
rect 112714 299780 113334 316263
rect 144994 308732 145614 319767
rect 148714 308732 149334 321588
rect 157286 318736 157906 334512
rect 158758 333424 159378 336240
rect 159494 333424 160114 336240
rect 161150 318736 161770 334512
rect 36994 236980 37614 253788
rect 21310 221904 21930 232880
rect 22046 221904 22666 232880
rect 36994 208964 37614 224988
rect 40714 208964 41334 253788
rect 53694 221904 54314 239408
rect 72994 236193 73614 278599
rect 76714 236193 77334 278599
rect 108994 277748 109614 287788
rect 112714 277748 113334 287788
rect 122510 285008 123130 302512
rect 126374 285008 126994 302512
rect 122878 275760 123498 280752
rect 126742 275760 127362 280752
rect 93254 256176 93874 273680
rect 97118 256176 97738 273680
rect 127294 257984 127914 273680
rect 131158 257984 131778 273680
rect 144994 270780 145614 278599
rect 148714 270780 149334 278599
rect 126926 255632 127546 257904
rect 130790 255632 131410 257904
rect 108994 236980 109614 253463
rect 112714 236980 113334 253463
rect 144994 245932 145614 256967
rect 148714 245932 149334 258788
rect 157286 257904 157906 273680
rect 158758 256176 159378 258992
rect 159494 256176 160114 258992
rect 161150 257904 161770 273680
rect 60318 196336 60938 208400
rect 36994 174180 37614 190988
rect 21310 159344 21930 170320
rect 22046 159344 22666 170320
rect 36994 146164 37614 162188
rect 40714 146164 41334 190988
rect 53694 159888 54314 176304
rect 72994 173393 73614 215799
rect 76714 173393 77334 215799
rect 108994 214948 109614 224988
rect 112714 214948 113334 224988
rect 122510 221904 123130 239952
rect 126374 221904 126994 239952
rect 122326 215920 122946 218192
rect 126190 215920 126810 218192
rect 122878 213200 123498 215840
rect 126742 213200 127362 215840
rect 93254 193072 93874 211120
rect 97118 193072 97738 211120
rect 127294 193072 127914 211120
rect 131158 193072 131778 211120
rect 144994 207980 145614 215799
rect 148714 207980 149334 215799
rect 108994 174180 109614 190663
rect 112714 174180 113334 190663
rect 144994 183132 145614 194167
rect 148714 183132 149334 195988
rect 157286 193072 157906 211120
rect 161150 193072 161770 211120
rect 122326 175120 122946 177392
rect 126190 175120 126810 177392
rect 36994 117980 37614 128188
rect 21310 103312 21930 107216
rect 22046 103312 22666 107216
rect 36994 83364 37614 105988
rect 40714 83364 41334 128188
rect 53694 103312 54314 120816
rect 72994 110593 73614 152999
rect 76714 110593 77334 152999
rect 108994 152148 109614 162188
rect 112714 152148 113334 162188
rect 122510 159344 123130 175040
rect 126374 159344 126994 175040
rect 122878 150096 123498 155088
rect 126742 150096 127362 155088
rect 93254 130512 93874 148016
rect 97118 130512 97738 148016
rect 127294 130512 127914 148016
rect 131158 130512 131778 148016
rect 144994 145180 145614 152999
rect 148714 145180 149334 152999
rect 108994 117980 109614 127863
rect 112714 117980 113334 127863
rect 36994 -7654 37614 65388
rect 40714 -7654 41334 65388
rect 66390 36400 67010 48464
rect 72994 -7654 73614 90199
rect 76714 -7654 77334 90199
rect 108994 89348 109614 105988
rect 112714 89348 113334 105988
rect 122510 103312 123130 120816
rect 126374 103312 126994 120816
rect 144994 120332 145614 131367
rect 148714 120332 149334 133188
rect 157286 130512 157906 148016
rect 161150 130512 161770 148016
rect 122878 87536 123498 92528
rect 126742 87536 127362 92528
rect 93254 65232 93874 82736
rect 97118 65232 97738 82736
rect 127294 67408 127914 85456
rect 131158 67408 131778 85456
rect 144994 82380 145614 90199
rect 148714 82380 149334 90199
rect 108994 55596 109614 65063
rect 112714 55596 113334 65063
rect 93254 33136 93874 50640
rect 97118 33136 97738 50640
rect 108994 -7654 109614 35988
rect 112714 -7654 113334 35988
rect 127294 33136 127914 50640
rect 131158 33136 131778 50640
rect 144994 47980 145614 68567
rect 148714 47980 149334 70388
rect 157286 67408 157906 85456
rect 161150 67408 161770 85456
rect 144994 -7654 145614 35988
rect 148714 12780 149334 35988
rect 157286 33136 157906 50640
rect 161150 33136 161770 50640
rect 180994 -7654 181614 711590
rect 184714 -7654 185334 711590
rect 216994 675793 217614 711590
rect 220714 675793 221334 711590
rect 188382 673424 189002 675696
rect 188382 670160 189002 672432
rect 188382 666896 189002 669168
rect 193166 633168 193786 650672
rect 216994 647580 217614 655399
rect 188382 611408 189002 613680
rect 216994 612993 217614 635588
rect 220714 612993 221334 655399
rect 221502 634800 222122 647952
rect 223158 647312 223778 650672
rect 223158 644048 223778 646320
rect 223158 640784 223778 643056
rect 223158 637520 223778 639792
rect 223158 633168 223778 636528
rect 225366 634800 225986 647952
rect 188382 608144 189002 610416
rect 188382 604880 189002 607152
rect 188382 601616 189002 603888
rect 188750 590736 189370 594096
rect 193166 568976 193786 586480
rect 216994 583580 217614 592599
rect 216994 550193 217614 571588
rect 220714 550193 221334 592599
rect 223158 568976 223778 586480
rect 188382 546128 189002 548400
rect 188382 542864 189002 545136
rect 188382 539600 189002 541872
rect 188750 527632 189370 532080
rect 193166 506960 193786 524464
rect 216994 521980 217614 529799
rect 216994 487393 217614 509988
rect 220714 487393 221334 529799
rect 223158 506960 223778 524464
rect 188382 484112 189002 486384
rect 188382 480848 189002 483120
rect 188382 477584 189002 479856
rect 188750 464528 189370 468976
rect 193166 444944 193786 461360
rect 216994 459180 217614 466999
rect 216994 424593 217614 447188
rect 220714 424593 221334 466999
rect 223158 444944 223778 461360
rect 188382 422096 189002 424368
rect 188382 418832 189002 421104
rect 188382 415568 189002 417840
rect 188750 401424 189370 405872
rect 193166 381840 193786 399344
rect 216994 396380 217614 404199
rect 188382 360080 189002 362352
rect 216994 361793 217614 384388
rect 220714 361793 221334 404199
rect 221502 383472 222122 396624
rect 223158 381840 223778 399344
rect 225366 383472 225986 396624
rect 188382 356816 189002 359088
rect 188382 353552 189002 355824
rect 188382 350288 189002 352560
rect 188750 339408 189370 342768
rect 193166 318736 193786 336240
rect 216994 333580 217614 341399
rect 216994 298993 217614 321588
rect 220714 298993 221334 341399
rect 223158 318736 223778 336240
rect 188382 294800 189002 297072
rect 188382 291536 189002 293808
rect 188382 288272 189002 290544
rect 188750 276304 189370 280752
rect 193166 257808 193786 273136
rect 216994 270780 217614 278599
rect 203654 255632 204274 257904
rect 188382 226256 189002 236144
rect 216994 236193 217614 258788
rect 220714 236193 221334 278599
rect 222054 256720 222674 258992
rect 223158 257904 223778 273136
rect 188750 213200 189370 217648
rect 193166 193616 193786 211120
rect 216994 207980 217614 215799
rect 188382 162064 189002 174128
rect 216994 173393 217614 195988
rect 220714 173393 221334 215799
rect 221502 195248 222122 208400
rect 223158 193616 223778 211120
rect 225366 195248 225986 208400
rect 188750 150096 189370 154544
rect 193166 130512 193786 148016
rect 216994 145180 217614 152999
rect 188382 113104 189002 115376
rect 188382 109840 189002 112112
rect 216994 110593 217614 133188
rect 220714 110593 221334 152999
rect 223158 130512 223778 148016
rect 188382 106576 189002 108848
rect 188750 88080 189370 92528
rect 193166 67408 193786 84912
rect 216994 82380 217614 90199
rect 193166 33680 193786 48912
rect 203654 48912 204274 51184
rect 216994 47980 217614 70388
rect 216994 -7654 217614 35988
rect 220714 -7654 221334 90199
rect 223158 67408 223778 84912
rect 221502 35312 222122 48464
rect 223158 47824 223778 50096
rect 223158 43472 223778 46832
rect 223158 38032 223778 41392
rect 223158 33680 223778 35952
rect 225366 35312 225986 48464
rect 252994 -7654 253614 711590
rect 256714 -7654 257334 711590
rect 288994 675793 289614 711590
rect 287190 632624 287810 650128
rect 288994 612993 289614 655399
rect 292714 647257 293334 711590
rect 314238 677776 314858 688208
rect 318102 677776 318722 688208
rect 314606 663808 315226 677696
rect 318470 663808 319090 677696
rect 314238 652752 314858 663728
rect 318102 652752 318722 663728
rect 287190 569520 287810 585936
rect 288994 550193 289614 592599
rect 292714 590713 293334 629175
rect 314238 614672 314858 625648
rect 318102 614672 318722 625648
rect 314606 600704 315226 614592
rect 318470 600704 319090 614592
rect 314238 592912 314858 600624
rect 318102 592912 318722 600624
rect 314790 590192 315410 592832
rect 318654 590192 319274 592832
rect 287190 507504 287810 525008
rect 288994 487393 289614 529799
rect 292714 527913 293334 567463
rect 314238 552112 314858 563088
rect 318102 552112 318722 563088
rect 314606 538144 315226 552032
rect 318470 538144 319090 552032
rect 314238 530352 314858 538064
rect 318102 530352 318722 538064
rect 314790 527088 315410 530272
rect 318654 527088 319274 530272
rect 287190 444400 287810 461904
rect 288994 424593 289614 466999
rect 292714 465113 293334 504663
rect 306878 489552 307498 499984
rect 310742 489552 311362 499984
rect 314606 475040 315226 491280
rect 318470 475040 319090 491280
rect 314238 467248 314858 474960
rect 318102 467248 318722 474960
rect 314790 464528 315410 467168
rect 318654 464528 319274 467168
rect 287190 381296 287810 398800
rect 288994 361793 289614 404199
rect 292714 402313 293334 441926
rect 314238 426448 314858 437424
rect 318102 426448 318722 437424
rect 314606 412480 315226 426368
rect 318470 412480 319090 426368
rect 314238 404688 314858 412400
rect 318102 404688 318722 412400
rect 314790 401424 315410 404608
rect 318654 401424 319274 404608
rect 287190 319280 287810 335696
rect 288994 298993 289614 341399
rect 292714 339513 293334 379063
rect 314238 363888 314858 374320
rect 318102 363888 318722 374320
rect 314606 349376 315226 363808
rect 318470 349376 319090 363808
rect 314238 341584 314858 349296
rect 318102 341584 318722 349296
rect 314790 338864 315410 341504
rect 318654 338864 319274 341504
rect 287190 256176 287810 273680
rect 288994 236193 289614 278599
rect 292714 276713 293334 316263
rect 314238 300784 314858 311760
rect 318102 300784 318722 311760
rect 314606 286816 315226 300704
rect 318470 286816 319090 300704
rect 314238 279024 314858 286736
rect 318102 279024 318722 286736
rect 314790 275760 315410 278944
rect 318654 275760 319274 278944
rect 287190 193072 287810 210576
rect 288994 173393 289614 215799
rect 292714 213913 293334 253463
rect 314238 238224 314858 248656
rect 318102 238224 318722 248656
rect 314606 223712 315226 238144
rect 318470 223712 319090 238144
rect 314238 215920 314858 223632
rect 318102 215920 318722 223632
rect 314790 213200 315410 215840
rect 318654 213200 319274 215840
rect 287190 131056 287810 147472
rect 288994 110593 289614 152999
rect 292714 151113 293334 190663
rect 314238 175120 314858 186096
rect 318102 175120 318722 186096
rect 314606 161152 315226 175040
rect 318470 161152 319090 175040
rect 314238 153360 314858 161072
rect 318102 153360 318722 161072
rect 314790 150096 315410 153280
rect 318654 150096 319274 153280
rect 287190 67952 287810 85456
rect 287190 33136 287810 50640
rect 288994 -7654 289614 90199
rect 292714 88313 293334 127863
rect 314238 119088 314858 122992
rect 318102 119088 318722 122992
rect 314606 105120 315226 119008
rect 318470 105120 319090 119008
rect 314238 90800 314858 105040
rect 318102 90800 318722 105040
rect 314790 87536 315410 90720
rect 318654 87536 319274 90720
rect 292714 -7654 293334 65063
rect 324994 -7654 325614 711590
rect 328714 675793 329334 711590
rect 360994 676580 361614 711590
rect 364714 676580 365334 711590
rect 328714 612993 329334 655399
rect 349382 632624 350002 650672
rect 353246 632624 353866 650672
rect 360994 647257 361614 664588
rect 364714 647257 365334 664588
rect 378454 663808 379074 679504
rect 382318 663808 382938 679504
rect 396994 675793 397614 711590
rect 400714 699892 401334 711590
rect 432994 676580 433614 711590
rect 378270 661456 378890 663728
rect 382134 661456 382754 663728
rect 383422 632624 384042 650672
rect 387286 632624 387906 650672
rect 360994 613780 361614 629175
rect 364714 613780 365334 629175
rect 378270 614672 378890 616944
rect 382134 614672 382754 616944
rect 328714 550193 329334 592599
rect 360994 590713 361614 601788
rect 364714 590713 365334 601788
rect 378454 598896 379074 614592
rect 382318 598896 382938 614592
rect 396994 612993 397614 655399
rect 400714 647580 401334 655399
rect 400714 622732 401334 635588
rect 413414 632624 414034 650672
rect 417278 632624 417898 650672
rect 432994 650196 433614 664588
rect 432994 613780 433614 629175
rect 378822 590192 379442 594640
rect 382686 590192 383306 594640
rect 349382 568976 350002 586480
rect 353246 568976 353866 586480
rect 383422 570784 384042 586480
rect 387286 570784 387906 586480
rect 382870 568432 383490 570704
rect 386734 568432 387354 570704
rect 360994 550980 361614 567463
rect 364714 550980 365334 567463
rect 328714 487393 329334 529799
rect 360994 527913 361614 538988
rect 364714 527913 365334 538988
rect 378454 538144 379074 553840
rect 382318 538144 382938 553840
rect 396994 550193 397614 592599
rect 400714 583580 401334 592599
rect 432994 591748 433614 601788
rect 413414 570704 414034 586480
rect 400714 559932 401334 569767
rect 414886 568976 415506 571792
rect 415622 568976 416242 571792
rect 417278 570704 417898 586480
rect 432994 550980 433614 567463
rect 378270 535792 378890 538064
rect 382134 535792 382754 538064
rect 378822 527088 379442 532080
rect 382686 527088 383306 532080
rect 349382 506960 350002 525008
rect 353246 506960 353866 525008
rect 383422 506960 384042 525008
rect 387286 506960 387906 525008
rect 360994 488180 361614 504663
rect 364714 488180 365334 504663
rect 328714 424593 329334 466999
rect 360994 465113 361614 476188
rect 364714 465113 365334 476188
rect 378454 473232 379074 491280
rect 382318 473232 382938 491280
rect 396994 487393 397614 529799
rect 400714 521980 401334 529799
rect 432994 528948 433614 538988
rect 400714 497132 401334 508167
rect 413414 506960 414034 525008
rect 417278 506960 417898 525008
rect 432994 488180 433614 504663
rect 378822 464528 379442 468976
rect 382686 464528 383306 468976
rect 349382 444400 350002 461904
rect 353246 444400 353866 461904
rect 383422 444400 384042 461904
rect 387286 444400 387906 461904
rect 360994 425380 361614 441863
rect 364714 425380 365334 441926
rect 328714 361793 329334 404199
rect 360994 402313 361614 413388
rect 364714 402313 365334 413388
rect 378454 410672 379074 428176
rect 382318 410672 382938 428176
rect 396994 424593 397614 466999
rect 400714 459180 401334 466999
rect 432994 466148 433614 476188
rect 400714 434332 401334 445367
rect 413414 444400 414034 461904
rect 417278 444400 417898 461904
rect 432994 425380 433614 441863
rect 378822 401424 379442 406416
rect 382686 401424 383306 406416
rect 349382 381296 350002 399344
rect 353246 381296 353866 399344
rect 383422 381296 384042 399344
rect 387286 381296 387906 399344
rect 360994 362580 361614 379063
rect 364714 362580 365334 379063
rect 328714 298993 329334 341399
rect 360994 339513 361614 350588
rect 364714 339513 365334 350588
rect 378454 347568 379074 365616
rect 382318 347568 382938 365616
rect 396994 361793 397614 404199
rect 400714 396380 401334 404199
rect 432994 403348 433614 413388
rect 400714 371532 401334 382567
rect 413414 381296 414034 399344
rect 417278 381296 417898 399344
rect 432994 362580 433614 379063
rect 378822 338864 379442 343312
rect 382686 338864 383306 343312
rect 349382 318736 350002 336240
rect 353246 318736 353866 336240
rect 377350 334512 377970 336784
rect 381214 334512 381834 336784
rect 383422 318736 384042 334512
rect 387286 318736 387906 334512
rect 360994 299780 361614 316263
rect 364714 299780 365334 316263
rect 328714 236193 329334 278599
rect 360994 276713 361614 287788
rect 364714 276713 365334 287788
rect 378454 285008 379074 302512
rect 382318 285008 382938 302512
rect 396994 298993 397614 341399
rect 400714 333580 401334 341399
rect 432994 340548 433614 350588
rect 400714 308732 401334 319767
rect 413414 318736 414034 334512
rect 414886 333424 415506 336240
rect 415622 333424 416242 336240
rect 417278 318736 417898 334512
rect 432994 299780 433614 316263
rect 378822 275760 379442 280752
rect 382686 275760 383306 280752
rect 349382 256176 350002 273680
rect 353246 256176 353866 273680
rect 383422 256176 384042 273680
rect 387286 256176 387906 273680
rect 360994 236980 361614 253463
rect 364714 236980 365334 253463
rect 328714 173393 329334 215799
rect 360994 213913 361614 224988
rect 364714 213913 365334 224988
rect 378454 221904 379074 239952
rect 382318 221904 382938 239952
rect 396994 236193 397614 278599
rect 400714 270780 401334 278599
rect 432994 277748 433614 287788
rect 400714 245932 401334 256967
rect 413414 256176 414034 273680
rect 417278 256176 417898 273680
rect 432994 236980 433614 253463
rect 378270 215920 378890 218192
rect 382134 215920 382754 218192
rect 378822 213200 379442 215840
rect 382686 213200 383306 215840
rect 349382 193072 350002 211120
rect 353246 193072 353866 211120
rect 383422 193072 384042 211120
rect 387286 193072 387906 211120
rect 360994 174180 361614 190663
rect 364714 174180 365334 190663
rect 378270 175120 378890 177392
rect 382134 175120 382754 177392
rect 328714 110593 329334 152999
rect 360994 151113 361614 162188
rect 364714 151113 365334 162188
rect 378454 159344 379074 175040
rect 382318 159344 382938 175040
rect 396994 173393 397614 215799
rect 400714 207980 401334 215799
rect 432994 214948 433614 224988
rect 400714 183132 401334 194167
rect 413414 193072 414034 211120
rect 417278 193072 417898 211120
rect 432994 174180 433614 190663
rect 378822 150096 379442 155088
rect 382686 150096 383306 155088
rect 349382 130512 350002 148016
rect 353246 130512 353866 148016
rect 383422 130512 384042 148016
rect 387286 130512 387906 148016
rect 360994 117980 361614 127863
rect 364714 117980 365334 127863
rect 328714 -7654 329334 90199
rect 360994 88313 361614 105988
rect 364714 88313 365334 105988
rect 378454 103312 379074 120816
rect 382318 103312 382938 120816
rect 396994 110593 397614 152999
rect 400714 145180 401334 152999
rect 432994 152148 433614 162188
rect 400714 120332 401334 131367
rect 413414 130512 414034 148016
rect 417278 130512 417898 148016
rect 432994 117980 433614 127863
rect 378822 87536 379442 92528
rect 382686 87536 383306 92528
rect 349382 67408 350002 85456
rect 353246 67408 353866 85456
rect 383422 67408 384042 85456
rect 387286 67408 387906 85456
rect 349382 33136 350002 50640
rect 353246 33136 353866 50640
rect 360994 -7654 361614 65063
rect 364714 -7654 365334 65063
rect 383422 33136 384042 50640
rect 387286 33136 387906 50640
rect 396994 -7654 397614 90199
rect 400714 82380 401334 90199
rect 432994 89348 433614 105988
rect 400714 47980 401334 68567
rect 413414 67408 414034 85456
rect 417278 67408 417898 85456
rect 432994 55596 433614 65063
rect 400714 -7654 401334 35988
rect 413414 33136 414034 50640
rect 417278 33136 417898 50640
rect 432994 -7654 433614 35988
rect 436714 -7654 437334 711590
rect 468994 685532 469614 711590
rect 472714 685532 473334 711590
rect 442486 663808 443106 679504
rect 446350 663808 446970 679504
rect 442302 661456 442922 663728
rect 446166 661456 446786 663728
rect 447270 632624 447890 650672
rect 451134 632624 451754 650672
rect 468994 647580 469614 655399
rect 472714 647580 473334 655399
rect 468994 622732 469614 635588
rect 472714 622732 473334 635588
rect 477262 632624 477882 650672
rect 481126 632624 481746 650672
rect 442302 614672 442922 616944
rect 446166 614672 446786 616944
rect 442486 598896 443106 614592
rect 446350 598896 446970 614592
rect 442854 590192 443474 594640
rect 446718 590192 447338 594640
rect 447270 568976 447890 586480
rect 451134 568976 451754 586480
rect 468994 583580 469614 592599
rect 472714 583580 473334 592599
rect 468994 559932 469614 571588
rect 472714 559932 473334 571588
rect 477262 568976 477882 586480
rect 481126 568976 481746 586480
rect 442486 536336 443106 553840
rect 446350 536336 446970 553840
rect 442854 527088 443474 532080
rect 446718 527088 447338 532080
rect 447270 506960 447890 525008
rect 451134 506960 451754 525008
rect 468994 521980 469614 529799
rect 472714 521980 473334 529799
rect 468994 497132 469614 509988
rect 472714 497132 473334 509988
rect 477262 506960 477882 525008
rect 481126 506960 481746 525008
rect 442486 473232 443106 491280
rect 446350 473232 446970 491280
rect 442854 464528 443474 468976
rect 446718 464528 447338 468976
rect 447270 444400 447890 461904
rect 451134 444400 451754 461904
rect 468994 459180 469614 466999
rect 472714 459180 473334 466999
rect 468994 434332 469614 447188
rect 472714 434332 473334 447188
rect 477262 444400 477882 461904
rect 481126 444400 481746 461904
rect 442486 410672 443106 428176
rect 446350 410672 446970 428176
rect 442854 401424 443474 406416
rect 446718 401424 447338 406416
rect 447270 381296 447890 399344
rect 451134 381296 451754 399344
rect 468994 396380 469614 404199
rect 472714 396380 473334 404199
rect 468994 371532 469614 384388
rect 472714 371532 473334 384388
rect 477262 381296 477882 399344
rect 481126 381296 481746 399344
rect 442486 347568 443106 365616
rect 446350 347568 446970 365616
rect 442854 338864 443474 343312
rect 446718 338864 447338 343312
rect 441382 334512 442002 336784
rect 445246 334512 445866 336784
rect 447270 318736 447890 334512
rect 451134 318736 451754 334512
rect 468994 333580 469614 341399
rect 472714 333580 473334 341399
rect 468994 308732 469614 321588
rect 472714 308732 473334 321588
rect 477262 318736 477882 334512
rect 478918 333424 479538 336240
rect 479654 333424 480274 336240
rect 481126 318736 481746 334512
rect 442486 285008 443106 302512
rect 446350 285008 446970 302512
rect 442854 275760 443474 280752
rect 446718 275760 447338 280752
rect 447270 256176 447890 273680
rect 451134 256176 451754 273680
rect 468994 270780 469614 278599
rect 472714 270780 473334 278599
rect 468994 245932 469614 258788
rect 472714 245932 473334 258788
rect 477262 256176 477882 273680
rect 481126 256176 481746 273680
rect 442486 221904 443106 239952
rect 446350 221904 446970 239952
rect 442854 213200 443474 217648
rect 446718 213200 447338 217648
rect 447270 193072 447890 211120
rect 451134 193072 451754 211120
rect 468994 207980 469614 215799
rect 472714 207980 473334 215799
rect 468994 183132 469614 195988
rect 472714 183132 473334 195988
rect 477262 193072 477882 211120
rect 481126 193072 481746 211120
rect 437702 175120 438322 177392
rect 441566 175120 442186 177392
rect 442486 159344 443106 175120
rect 446350 159344 446970 175120
rect 442854 150096 443474 155088
rect 446718 150096 447338 155088
rect 447270 130512 447890 148016
rect 451134 130512 451754 148016
rect 468994 145180 469614 152999
rect 472714 145180 473334 152999
rect 442486 103312 443106 120816
rect 446350 103312 446970 120816
rect 468994 120332 469614 133188
rect 472714 120332 473334 133188
rect 477262 130512 477882 148016
rect 481126 130512 481746 148016
rect 442854 87536 443474 92528
rect 446718 87536 447338 92528
rect 447270 67408 447890 85456
rect 451134 67408 451754 85456
rect 468994 82380 469614 90199
rect 472714 82380 473334 90199
rect 447270 33136 447890 50640
rect 451134 33136 451754 50640
rect 468994 47980 469614 70388
rect 472714 47980 473334 70388
rect 477262 67408 477882 85456
rect 481126 67408 481746 85456
rect 468994 12780 469614 35988
rect 472714 -7654 473334 35988
rect 477262 33136 477882 50640
rect 481126 33136 481746 50640
rect 504994 -7654 505614 711590
rect 508714 -7654 509334 711590
rect 540994 675793 541614 711590
rect 544714 675793 545334 711590
rect 566502 663808 567122 674608
rect 567238 663808 567858 674608
rect 540994 612993 541614 655399
rect 544714 612993 545334 655399
rect 565950 652752 566570 663728
rect 566686 652752 567306 663728
rect 566502 600704 567122 611504
rect 567238 600704 567858 611504
rect 540994 550193 541614 592599
rect 544714 550193 545334 592599
rect 565950 590192 566570 600624
rect 566686 590192 567306 600624
rect 566502 538144 567122 548944
rect 567238 538144 567858 548944
rect 540994 487393 541614 529799
rect 543134 509136 543754 522288
rect 544714 487393 545334 529799
rect 565950 527088 566570 538064
rect 566686 527088 567306 538064
rect 540994 424593 541614 466999
rect 544714 424593 545334 466999
rect 562086 464528 562706 474960
rect 565950 464528 566570 474960
rect 567422 473776 568042 485840
rect 568158 473776 568778 485840
rect 566502 412480 567122 423280
rect 567238 412480 567858 423280
rect 540994 361793 541614 404199
rect 544714 361793 545334 404199
rect 565950 401424 566570 412400
rect 566686 401424 567306 412400
rect 540994 298993 541614 341399
rect 543134 320912 543754 334064
rect 544714 298993 545334 341399
rect 562086 338864 562706 349296
rect 565950 338864 566570 349296
rect 567422 347568 568042 360720
rect 568158 347568 568778 360720
rect 566502 286816 567122 297616
rect 567238 286816 567858 297616
rect 540994 236193 541614 278599
rect 544714 236193 545334 278599
rect 565950 275760 566570 286736
rect 566686 275760 567306 286736
rect 540994 173393 541614 215799
rect 544714 173393 545334 215799
rect 562086 213200 562706 223632
rect 565950 213200 566570 223632
rect 567422 222448 568042 235056
rect 568158 222448 568778 235056
rect 566502 161152 567122 171952
rect 567238 161152 567858 171952
rect 540994 110593 541614 152999
rect 544714 110593 545334 152999
rect 565950 150096 566570 161072
rect 566686 150096 567306 161072
rect 566502 105120 567122 109392
rect 567238 105120 567858 109392
rect 540994 -7654 541614 90199
rect 543134 69584 543754 82736
rect 544714 -7654 545334 90199
rect 565950 87536 566570 105040
rect 566686 87536 567306 105040
rect 576994 -7654 577614 711590
rect 579750 652752 580370 674608
rect 579750 590736 580370 611504
rect 579750 527632 580370 548400
rect 579750 464528 580370 485296
rect 579750 401424 580370 423280
rect 579750 339408 580370 360176
rect 579750 276304 580370 297072
rect 579750 213200 580370 235056
rect 579750 150096 580370 171952
rect 579750 88080 580370 108848
rect 580714 -7654 581334 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 13415 676500 36914 697752
rect 37694 676500 40634 697752
rect 13415 672512 40634 676500
rect 13415 661920 21230 672512
rect 22746 664668 40634 672512
rect 22746 661920 36914 664668
rect 13415 613700 36914 661920
rect 37694 613700 40634 664668
rect 13415 609952 40634 613700
rect 13415 598816 21230 609952
rect 22746 601868 40634 609952
rect 22746 598816 36914 601868
rect 13415 585684 36914 598816
rect 37694 585684 40634 601868
rect 41414 679040 72914 697752
rect 41414 662464 53614 679040
rect 54394 675713 72914 679040
rect 73694 675713 76634 697752
rect 77414 676500 108914 697752
rect 109694 676500 112634 697752
rect 113414 685452 148634 697752
rect 149414 685452 180914 697752
rect 113414 679584 180914 685452
rect 113414 676500 122430 679584
rect 77414 675713 122430 676500
rect 54394 664668 122430 675713
rect 54394 662464 108914 664668
rect 41414 655479 108914 662464
rect 41414 615936 72914 655479
rect 41414 599360 53614 615936
rect 54394 612913 72914 615936
rect 73694 612913 76634 655479
rect 77414 650752 108914 655479
rect 77414 632544 93174 650752
rect 93954 632544 97038 650752
rect 97818 650116 108914 650752
rect 109694 650116 112634 664668
rect 113414 661920 122430 664668
rect 123210 661920 126294 679584
rect 127074 661920 180914 679584
rect 113414 655479 180914 661920
rect 113414 650752 144914 655479
rect 113414 650116 127214 650752
rect 97818 632544 127214 650116
rect 127994 632544 131078 650752
rect 131858 647500 144914 650752
rect 145694 647500 148634 655479
rect 149414 650752 180914 655479
rect 149414 647500 157206 650752
rect 131858 635668 157206 647500
rect 131858 632544 144914 635668
rect 77414 629255 144914 632544
rect 77414 613700 108914 629255
rect 109694 613700 112634 629255
rect 113414 622652 144914 629255
rect 145694 622652 148634 635668
rect 149414 632544 157206 635668
rect 157986 632544 161070 650752
rect 161850 632544 180914 650752
rect 149414 622652 180914 632544
rect 113414 617024 180914 622652
rect 113414 614592 122246 617024
rect 123026 614672 126110 617024
rect 126890 614672 180914 617024
rect 123210 614592 126110 614672
rect 113414 613700 122430 614592
rect 77414 612913 122430 613700
rect 54394 601868 122430 612913
rect 54394 599360 108914 601868
rect 41414 592679 108914 599360
rect 41414 585684 72914 592679
rect 13415 567868 72914 585684
rect 13415 550900 36914 567868
rect 37694 550900 40634 567868
rect 13415 546848 40634 550900
rect 13415 536256 21230 546848
rect 22746 539068 40634 546848
rect 22746 536256 36914 539068
rect 13415 522884 36914 536256
rect 37694 522884 40634 539068
rect 41414 553920 72914 567868
rect 41414 536256 53614 553920
rect 54394 550113 72914 553920
rect 73694 550113 76634 592679
rect 77414 591668 108914 592679
rect 109694 591668 112634 601868
rect 113414 598816 122430 601868
rect 123210 598816 126294 614592
rect 127074 598816 180914 614672
rect 113414 594720 180914 598816
rect 113414 591668 122798 594720
rect 77414 591200 122798 591668
rect 123578 591920 126662 594720
rect 127442 592679 180914 594720
rect 127442 592000 144914 592679
rect 123578 591200 126846 591920
rect 77414 589568 126846 591200
rect 127626 589568 130710 592000
rect 131490 589568 144914 592000
rect 77414 586560 144914 589568
rect 77414 568896 93174 586560
rect 93954 568896 97038 586560
rect 97818 570784 127214 586560
rect 127994 570784 131078 586560
rect 131858 583500 144914 586560
rect 145694 583500 148634 592679
rect 149414 586560 180914 592679
rect 149414 583500 157206 586560
rect 131858 571668 157206 583500
rect 97818 568896 126846 570784
rect 127994 570704 130710 570784
rect 131858 570704 148634 571668
rect 77414 568352 126846 568896
rect 127626 568352 130710 570704
rect 131490 569847 148634 570704
rect 131490 568352 144914 569847
rect 77414 567543 144914 568352
rect 77414 550900 108914 567543
rect 109694 550900 112634 567543
rect 113414 559852 144914 567543
rect 145694 559852 148634 569847
rect 149414 570624 157206 571668
rect 157986 571872 161070 586560
rect 157986 570624 158678 571872
rect 149414 568896 158678 570624
rect 160194 570624 161070 571872
rect 161850 570624 180914 586560
rect 160194 568896 180914 570624
rect 149414 559852 180914 568896
rect 113414 553920 180914 559852
rect 113414 550900 122430 553920
rect 77414 550113 122430 550900
rect 54394 539068 122430 550113
rect 54394 536256 108914 539068
rect 41414 529879 108914 536256
rect 41414 522884 72914 529879
rect 13415 505068 72914 522884
rect 13415 488100 36914 505068
rect 37694 488100 40634 505068
rect 13415 484288 40634 488100
rect 13415 473152 21230 484288
rect 22746 476268 40634 484288
rect 22746 473152 36914 476268
rect 13415 460084 36914 473152
rect 37694 460084 40634 476268
rect 41414 490816 72914 505068
rect 41414 473152 53614 490816
rect 54394 487313 72914 490816
rect 73694 487313 76634 529879
rect 77414 528868 108914 529879
rect 109694 528868 112634 539068
rect 113414 536256 122430 539068
rect 123210 536256 126294 553920
rect 127074 536256 180914 553920
rect 113414 532160 180914 536256
rect 113414 528868 122798 532160
rect 77414 527008 122798 528868
rect 123578 527008 126662 532160
rect 127442 529879 180914 532160
rect 127442 527008 144914 529879
rect 77414 525088 144914 527008
rect 77414 506880 93174 525088
rect 93954 506880 97038 525088
rect 97818 506880 127214 525088
rect 127994 506880 131078 525088
rect 131858 521900 144914 525088
rect 145694 521900 148634 529879
rect 149414 525088 180914 529879
rect 149414 521900 157206 525088
rect 131858 510068 157206 521900
rect 131858 508247 148634 510068
rect 131858 506880 144914 508247
rect 77414 504743 144914 506880
rect 77414 488100 108914 504743
rect 109694 488100 112634 504743
rect 113414 497052 144914 504743
rect 145694 497052 148634 508247
rect 149414 506880 157206 510068
rect 157986 506880 161070 525088
rect 161850 506880 180914 525088
rect 149414 497052 180914 506880
rect 113414 491360 180914 497052
rect 113414 488100 122430 491360
rect 77414 487313 122430 488100
rect 54394 476268 122430 487313
rect 54394 473152 108914 476268
rect 41414 467079 108914 473152
rect 41414 460084 72914 467079
rect 13415 442268 72914 460084
rect 13415 425300 36914 442268
rect 37694 425300 40634 442268
rect 13415 421184 40634 425300
rect 13415 410592 21230 421184
rect 22746 413468 40634 421184
rect 22746 410592 36914 413468
rect 13415 397284 36914 410592
rect 37694 397284 40634 413468
rect 41414 427712 72914 442268
rect 41414 411136 53614 427712
rect 54394 424513 72914 427712
rect 73694 424513 76634 467079
rect 77414 466068 108914 467079
rect 109694 466068 112634 476268
rect 113414 473152 122430 476268
rect 123210 473152 126294 491360
rect 127074 473152 180914 491360
rect 113414 469056 180914 473152
rect 113414 466068 122798 469056
rect 77414 464448 122798 466068
rect 123578 464448 126662 469056
rect 127442 467079 180914 469056
rect 127442 464448 144914 467079
rect 77414 461984 144914 464448
rect 77414 444320 93174 461984
rect 93954 444320 97038 461984
rect 97818 444320 127214 461984
rect 127994 444320 131078 461984
rect 131858 459100 144914 461984
rect 145694 459100 148634 467079
rect 149414 461984 180914 467079
rect 149414 459100 157206 461984
rect 131858 447268 157206 459100
rect 131858 445447 148634 447268
rect 131858 444320 144914 445447
rect 77414 442006 144914 444320
rect 77414 441943 112634 442006
rect 77414 425300 108914 441943
rect 109694 425300 112634 441943
rect 113414 434252 144914 442006
rect 145694 434252 148634 445447
rect 149414 444320 157206 447268
rect 157986 444320 161070 461984
rect 161850 444320 180914 461984
rect 149414 434252 180914 444320
rect 113414 428256 180914 434252
rect 113414 425300 122430 428256
rect 77414 424513 122430 425300
rect 54394 413468 122430 424513
rect 54394 411136 108914 413468
rect 41414 404279 108914 411136
rect 41414 397284 72914 404279
rect 13415 396704 72914 397284
rect 13415 384480 60238 396704
rect 61018 384480 72914 396704
rect 13415 379468 72914 384480
rect 13415 362500 36914 379468
rect 37694 362500 40634 379468
rect 13415 358624 40634 362500
rect 13415 347488 21230 358624
rect 22746 350668 40634 358624
rect 22746 347488 36914 350668
rect 13415 334484 36914 347488
rect 37694 334484 40634 350668
rect 41414 365696 72914 379468
rect 41414 348032 53614 365696
rect 54394 361713 72914 365696
rect 73694 361713 76634 404279
rect 77414 403268 108914 404279
rect 109694 403268 112634 413468
rect 113414 410592 122430 413468
rect 123210 410592 126294 428256
rect 127074 410592 180914 428256
rect 113414 406496 180914 410592
rect 113414 403268 122798 406496
rect 77414 401344 122798 403268
rect 123578 401344 126662 406496
rect 127442 404279 180914 406496
rect 127442 401344 144914 404279
rect 77414 399424 144914 401344
rect 77414 381216 93174 399424
rect 93954 381216 97038 399424
rect 97818 381216 127214 399424
rect 127994 381216 131078 399424
rect 131858 396300 144914 399424
rect 145694 396300 148634 404279
rect 149414 399424 180914 404279
rect 149414 396300 157206 399424
rect 131858 384468 157206 396300
rect 131858 382647 148634 384468
rect 131858 381216 144914 382647
rect 77414 379143 144914 381216
rect 77414 362500 108914 379143
rect 109694 362500 112634 379143
rect 113414 371452 144914 379143
rect 145694 371452 148634 382647
rect 149414 381216 157206 384468
rect 157986 381216 161070 399424
rect 161850 381216 180914 399424
rect 149414 371452 180914 381216
rect 113414 365696 180914 371452
rect 113414 362500 122430 365696
rect 77414 361713 122430 362500
rect 54394 350668 122430 361713
rect 54394 348032 108914 350668
rect 41414 341479 108914 348032
rect 41414 334484 72914 341479
rect 13415 316668 72914 334484
rect 13415 299700 36914 316668
rect 37694 299700 40634 316668
rect 13415 295520 40634 299700
rect 13415 284928 21230 295520
rect 22746 287868 40634 295520
rect 22746 284928 36914 287868
rect 13415 271684 36914 284928
rect 37694 271684 40634 287868
rect 41414 302592 72914 316668
rect 41414 284928 53614 302592
rect 54394 298913 72914 302592
rect 73694 298913 76634 341479
rect 77414 340468 108914 341479
rect 109694 340468 112634 350668
rect 113414 347488 122430 350668
rect 123210 347488 126294 365696
rect 127074 347488 180914 365696
rect 113414 343392 180914 347488
rect 113414 340468 122798 343392
rect 77414 338784 122798 340468
rect 123578 338784 126662 343392
rect 127442 341479 180914 343392
rect 127442 338784 144914 341479
rect 77414 336864 144914 338784
rect 77414 336320 121326 336864
rect 77414 318656 93174 336320
rect 93954 318656 97038 336320
rect 97818 334432 121326 336320
rect 122106 334432 125190 336864
rect 125970 334592 144914 336864
rect 125970 334432 127214 334592
rect 97818 318656 127214 334432
rect 127994 318656 131078 334592
rect 131858 333500 144914 334592
rect 145694 333500 148634 341479
rect 149414 336320 180914 341479
rect 149414 334592 158678 336320
rect 149414 333500 157206 334592
rect 131858 321668 157206 333500
rect 131858 319847 148634 321668
rect 131858 318656 144914 319847
rect 77414 316343 144914 318656
rect 77414 299700 108914 316343
rect 109694 299700 112634 316343
rect 113414 308652 144914 316343
rect 145694 308652 148634 319847
rect 149414 318656 157206 321668
rect 157986 333344 158678 334592
rect 160194 334592 180914 336320
rect 160194 333344 161070 334592
rect 157986 318656 161070 333344
rect 161850 318656 180914 334592
rect 149414 308652 180914 318656
rect 113414 302592 180914 308652
rect 113414 299700 122430 302592
rect 77414 298913 122430 299700
rect 54394 287868 122430 298913
rect 54394 284928 108914 287868
rect 41414 278679 108914 284928
rect 41414 271684 72914 278679
rect 13415 253868 72914 271684
rect 13415 236900 36914 253868
rect 37694 236900 40634 253868
rect 13415 232960 40634 236900
rect 13415 221824 21230 232960
rect 22746 225068 40634 232960
rect 22746 221824 36914 225068
rect 13415 208884 36914 221824
rect 37694 208884 40634 225068
rect 41414 239488 72914 253868
rect 41414 221824 53614 239488
rect 54394 236113 72914 239488
rect 73694 236113 76634 278679
rect 77414 277668 108914 278679
rect 109694 277668 112634 287868
rect 113414 284928 122430 287868
rect 123210 284928 126294 302592
rect 127074 284928 180914 302592
rect 113414 280832 180914 284928
rect 113414 277668 122798 280832
rect 77414 275680 122798 277668
rect 123578 275680 126662 280832
rect 127442 278679 180914 280832
rect 127442 275680 144914 278679
rect 77414 273760 144914 275680
rect 77414 256096 93174 273760
rect 93954 256096 97038 273760
rect 97818 257984 127214 273760
rect 127994 257984 131078 273760
rect 131858 270700 144914 273760
rect 145694 270700 148634 278679
rect 149414 273760 180914 278679
rect 149414 270700 157206 273760
rect 131858 258868 157206 270700
rect 97818 256096 126846 257984
rect 127994 257904 130710 257984
rect 131858 257904 148634 258868
rect 77414 255552 126846 256096
rect 127626 255552 130710 257904
rect 131490 257047 148634 257904
rect 131490 255552 144914 257047
rect 77414 253543 144914 255552
rect 77414 236900 108914 253543
rect 109694 236900 112634 253543
rect 113414 245852 144914 253543
rect 145694 245852 148634 257047
rect 149414 257824 157206 258868
rect 157986 259072 161070 273760
rect 157986 257824 158678 259072
rect 149414 256096 158678 257824
rect 160194 257824 161070 259072
rect 161850 257824 180914 273760
rect 160194 256096 180914 257824
rect 149414 245852 180914 256096
rect 113414 240032 180914 245852
rect 113414 236900 122430 240032
rect 77414 236113 122430 236900
rect 54394 225068 122430 236113
rect 54394 221824 108914 225068
rect 41414 215879 108914 221824
rect 41414 208884 72914 215879
rect 13415 208480 72914 208884
rect 13415 196256 60238 208480
rect 61018 196256 72914 208480
rect 13415 191068 72914 196256
rect 13415 174100 36914 191068
rect 37694 174100 40634 191068
rect 13415 170400 40634 174100
rect 13415 159264 21230 170400
rect 22746 162268 40634 170400
rect 22746 159264 36914 162268
rect 13415 146084 36914 159264
rect 37694 146084 40634 162268
rect 41414 176384 72914 191068
rect 41414 159808 53614 176384
rect 54394 173313 72914 176384
rect 73694 173313 76634 215879
rect 77414 214868 108914 215879
rect 109694 214868 112634 225068
rect 113414 221824 122430 225068
rect 123210 221824 126294 240032
rect 127074 221824 180914 240032
rect 113414 218272 180914 221824
rect 113414 215840 122246 218272
rect 123026 215920 126110 218272
rect 126890 215920 180914 218272
rect 123578 215840 126110 215920
rect 127442 215879 180914 215920
rect 113414 214868 122798 215840
rect 77414 213120 122798 214868
rect 123578 213120 126662 215840
rect 127442 213120 144914 215879
rect 77414 211200 144914 213120
rect 77414 192992 93174 211200
rect 93954 192992 97038 211200
rect 97818 192992 127214 211200
rect 127994 192992 131078 211200
rect 131858 207900 144914 211200
rect 145694 207900 148634 215879
rect 149414 211200 180914 215879
rect 149414 207900 157206 211200
rect 131858 196068 157206 207900
rect 131858 194247 148634 196068
rect 131858 192992 144914 194247
rect 77414 190743 144914 192992
rect 77414 174100 108914 190743
rect 109694 174100 112634 190743
rect 113414 183052 144914 190743
rect 145694 183052 148634 194247
rect 149414 192992 157206 196068
rect 157986 192992 161070 211200
rect 161850 192992 180914 211200
rect 149414 183052 180914 192992
rect 113414 177472 180914 183052
rect 113414 175040 122246 177472
rect 123026 175120 126110 177472
rect 126890 175120 180914 177472
rect 123210 175040 126110 175120
rect 113414 174100 122430 175040
rect 77414 173313 122430 174100
rect 54394 162268 122430 173313
rect 54394 159808 108914 162268
rect 41414 153079 108914 159808
rect 41414 146084 72914 153079
rect 13415 128268 72914 146084
rect 13415 117900 36914 128268
rect 37694 117900 40634 128268
rect 13415 107296 40634 117900
rect 13415 103232 21230 107296
rect 22746 106068 40634 107296
rect 22746 103232 36914 106068
rect 13415 83284 36914 103232
rect 37694 83284 40634 106068
rect 41414 120896 72914 128268
rect 41414 103232 53614 120896
rect 54394 110513 72914 120896
rect 73694 110513 76634 153079
rect 77414 152068 108914 153079
rect 109694 152068 112634 162268
rect 113414 159264 122430 162268
rect 123210 159264 126294 175040
rect 127074 159264 180914 175120
rect 113414 155168 180914 159264
rect 113414 152068 122798 155168
rect 77414 150016 122798 152068
rect 123578 150016 126662 155168
rect 127442 153079 180914 155168
rect 127442 150016 144914 153079
rect 77414 148096 144914 150016
rect 77414 130432 93174 148096
rect 93954 130432 97038 148096
rect 97818 130432 127214 148096
rect 127994 130432 131078 148096
rect 131858 145100 144914 148096
rect 145694 145100 148634 153079
rect 149414 148096 180914 153079
rect 149414 145100 157206 148096
rect 131858 133268 157206 145100
rect 131858 131447 148634 133268
rect 131858 130432 144914 131447
rect 77414 127943 144914 130432
rect 77414 117900 108914 127943
rect 109694 117900 112634 127943
rect 113414 120896 144914 127943
rect 113414 117900 122430 120896
rect 77414 110513 122430 117900
rect 54394 106068 122430 110513
rect 54394 103232 108914 106068
rect 41414 90279 108914 103232
rect 41414 83284 72914 90279
rect 13415 65468 72914 83284
rect 13415 2928 36914 65468
rect 37694 2928 40634 65468
rect 41414 48544 72914 65468
rect 41414 36320 66310 48544
rect 67090 36320 72914 48544
rect 41414 2928 72914 36320
rect 73694 2928 76634 90279
rect 77414 89268 108914 90279
rect 109694 89268 112634 106068
rect 113414 103232 122430 106068
rect 123210 103232 126294 120896
rect 127074 120252 144914 120896
rect 145694 120252 148634 131447
rect 149414 130432 157206 133268
rect 157986 130432 161070 148096
rect 161850 130432 180914 148096
rect 149414 120252 180914 130432
rect 127074 103232 180914 120252
rect 113414 92608 180914 103232
rect 113414 89268 122798 92608
rect 77414 87456 122798 89268
rect 123578 87456 126662 92608
rect 127442 90279 180914 92608
rect 127442 87456 144914 90279
rect 77414 85536 144914 87456
rect 77414 82816 127214 85536
rect 77414 65152 93174 82816
rect 93954 65152 97038 82816
rect 97818 67328 127214 82816
rect 127994 67328 131078 85536
rect 131858 82300 144914 85536
rect 145694 82300 148634 90279
rect 149414 85536 180914 90279
rect 149414 82300 157206 85536
rect 131858 70468 157206 82300
rect 131858 68647 148634 70468
rect 131858 67328 144914 68647
rect 97818 65152 144914 67328
rect 77414 65143 144914 65152
rect 77414 55516 108914 65143
rect 109694 55516 112634 65143
rect 113414 55516 144914 65143
rect 77414 50720 144914 55516
rect 77414 33056 93174 50720
rect 93954 33056 97038 50720
rect 97818 36068 127214 50720
rect 97818 33056 108914 36068
rect 77414 2928 108914 33056
rect 109694 2928 112634 36068
rect 113414 33056 127214 36068
rect 127994 33056 131078 50720
rect 131858 47900 144914 50720
rect 145694 47900 148634 68647
rect 149414 67328 157206 70468
rect 157986 67328 161070 85536
rect 161850 67328 180914 85536
rect 149414 50720 180914 67328
rect 149414 47900 157206 50720
rect 131858 36068 157206 47900
rect 131858 33056 144914 36068
rect 113414 2928 144914 33056
rect 145694 12700 148634 36068
rect 149414 33056 157206 36068
rect 157986 33056 161070 50720
rect 161850 33056 180914 50720
rect 149414 12700 180914 33056
rect 145694 2928 180914 12700
rect 181694 2928 184634 697752
rect 185414 675776 216914 697752
rect 185414 673344 188302 675776
rect 189082 675713 216914 675776
rect 217694 675713 220634 697752
rect 221414 675713 252914 697752
rect 189082 673344 252914 675713
rect 185414 672512 252914 673344
rect 185414 670080 188302 672512
rect 189082 670080 252914 672512
rect 185414 669248 252914 670080
rect 185414 666816 188302 669248
rect 189082 666816 252914 669248
rect 185414 655479 252914 666816
rect 185414 650752 216914 655479
rect 185414 633088 193086 650752
rect 193866 647500 216914 650752
rect 217694 647500 220634 655479
rect 193866 635668 220634 647500
rect 193866 633088 216914 635668
rect 185414 613760 216914 633088
rect 185414 611328 188302 613760
rect 189082 612913 216914 613760
rect 217694 612913 220634 635668
rect 221414 650752 252914 655479
rect 221414 648032 223078 650752
rect 221414 634720 221422 648032
rect 222202 647232 223078 648032
rect 223858 648032 252914 650752
rect 223858 647232 225286 648032
rect 222202 646400 225286 647232
rect 222202 643968 223078 646400
rect 223858 643968 225286 646400
rect 222202 643136 225286 643968
rect 222202 640704 223078 643136
rect 223858 640704 225286 643136
rect 222202 639872 225286 640704
rect 222202 637440 223078 639872
rect 223858 637440 225286 639872
rect 222202 636608 225286 637440
rect 222202 634720 223078 636608
rect 221414 633088 223078 634720
rect 223858 634720 225286 636608
rect 226066 634720 252914 648032
rect 223858 633088 252914 634720
rect 221414 612913 252914 633088
rect 189082 611328 252914 612913
rect 185414 610496 252914 611328
rect 185414 608064 188302 610496
rect 189082 608064 252914 610496
rect 185414 607232 252914 608064
rect 185414 604800 188302 607232
rect 189082 604800 252914 607232
rect 185414 603968 252914 604800
rect 185414 601536 188302 603968
rect 189082 601536 252914 603968
rect 185414 594176 252914 601536
rect 185414 590656 188670 594176
rect 189450 592679 252914 594176
rect 189450 590656 216914 592679
rect 185414 586560 216914 590656
rect 185414 568896 193086 586560
rect 193866 583500 216914 586560
rect 217694 583500 220634 592679
rect 193866 571668 220634 583500
rect 193866 568896 216914 571668
rect 185414 550113 216914 568896
rect 217694 550113 220634 571668
rect 221414 586560 252914 592679
rect 221414 568896 223078 586560
rect 223858 568896 252914 586560
rect 221414 550113 252914 568896
rect 185414 548480 252914 550113
rect 185414 546048 188302 548480
rect 189082 546048 252914 548480
rect 185414 545216 252914 546048
rect 185414 542784 188302 545216
rect 189082 542784 252914 545216
rect 185414 541952 252914 542784
rect 185414 539520 188302 541952
rect 189082 539520 252914 541952
rect 185414 532160 252914 539520
rect 185414 527552 188670 532160
rect 189450 529879 252914 532160
rect 189450 527552 216914 529879
rect 185414 524544 216914 527552
rect 185414 506880 193086 524544
rect 193866 521900 216914 524544
rect 217694 521900 220634 529879
rect 193866 510068 220634 521900
rect 193866 506880 216914 510068
rect 185414 487313 216914 506880
rect 217694 487313 220634 510068
rect 221414 524544 252914 529879
rect 221414 506880 223078 524544
rect 223858 506880 252914 524544
rect 221414 487313 252914 506880
rect 185414 486464 252914 487313
rect 185414 484032 188302 486464
rect 189082 484032 252914 486464
rect 185414 483200 252914 484032
rect 185414 480768 188302 483200
rect 189082 480768 252914 483200
rect 185414 479936 252914 480768
rect 185414 477504 188302 479936
rect 189082 477504 252914 479936
rect 185414 469056 252914 477504
rect 185414 464448 188670 469056
rect 189450 467079 252914 469056
rect 189450 464448 216914 467079
rect 185414 461440 216914 464448
rect 185414 444864 193086 461440
rect 193866 459100 216914 461440
rect 217694 459100 220634 467079
rect 193866 447268 220634 459100
rect 193866 444864 216914 447268
rect 185414 424513 216914 444864
rect 217694 424513 220634 447268
rect 221414 461440 252914 467079
rect 221414 444864 223078 461440
rect 223858 444864 252914 461440
rect 221414 424513 252914 444864
rect 185414 424448 252914 424513
rect 185414 422016 188302 424448
rect 189082 422016 252914 424448
rect 185414 421184 252914 422016
rect 185414 418752 188302 421184
rect 189082 418752 252914 421184
rect 185414 417920 252914 418752
rect 185414 415488 188302 417920
rect 189082 415488 252914 417920
rect 185414 405952 252914 415488
rect 185414 401344 188670 405952
rect 189450 404279 252914 405952
rect 189450 401344 216914 404279
rect 185414 399424 216914 401344
rect 185414 381760 193086 399424
rect 193866 396300 216914 399424
rect 217694 396300 220634 404279
rect 193866 384468 220634 396300
rect 193866 381760 216914 384468
rect 185414 362432 216914 381760
rect 185414 360000 188302 362432
rect 189082 361713 216914 362432
rect 217694 361713 220634 384468
rect 221414 399424 252914 404279
rect 221414 396704 223078 399424
rect 221414 383392 221422 396704
rect 222202 383392 223078 396704
rect 221414 381760 223078 383392
rect 223858 396704 252914 399424
rect 223858 383392 225286 396704
rect 226066 383392 252914 396704
rect 223858 381760 252914 383392
rect 221414 361713 252914 381760
rect 189082 360000 252914 361713
rect 185414 359168 252914 360000
rect 185414 356736 188302 359168
rect 189082 356736 252914 359168
rect 185414 355904 252914 356736
rect 185414 353472 188302 355904
rect 189082 353472 252914 355904
rect 185414 352640 252914 353472
rect 185414 350208 188302 352640
rect 189082 350208 252914 352640
rect 185414 342848 252914 350208
rect 185414 339328 188670 342848
rect 189450 341479 252914 342848
rect 189450 339328 216914 341479
rect 185414 336320 216914 339328
rect 185414 318656 193086 336320
rect 193866 333500 216914 336320
rect 217694 333500 220634 341479
rect 193866 321668 220634 333500
rect 193866 318656 216914 321668
rect 185414 298913 216914 318656
rect 217694 298913 220634 321668
rect 221414 336320 252914 341479
rect 221414 318656 223078 336320
rect 223858 318656 252914 336320
rect 221414 298913 252914 318656
rect 185414 297152 252914 298913
rect 185414 294720 188302 297152
rect 189082 294720 252914 297152
rect 185414 293888 252914 294720
rect 185414 291456 188302 293888
rect 189082 291456 252914 293888
rect 185414 290624 252914 291456
rect 185414 288192 188302 290624
rect 189082 288192 252914 290624
rect 185414 280832 252914 288192
rect 185414 276224 188670 280832
rect 189450 278679 252914 280832
rect 189450 276224 216914 278679
rect 185414 273216 216914 276224
rect 185414 257728 193086 273216
rect 193866 270700 216914 273216
rect 217694 270700 220634 278679
rect 193866 258868 220634 270700
rect 193866 257984 216914 258868
rect 193866 257728 203574 257984
rect 185414 255552 203574 257728
rect 204354 255552 216914 257984
rect 185414 236224 216914 255552
rect 185414 226176 188302 236224
rect 189082 236113 216914 236224
rect 217694 236113 220634 258868
rect 221414 273216 252914 278679
rect 221414 259072 223078 273216
rect 221414 256640 221974 259072
rect 222754 257824 223078 259072
rect 223858 257824 252914 273216
rect 222754 256640 252914 257824
rect 221414 236113 252914 256640
rect 189082 226176 252914 236113
rect 185414 217728 252914 226176
rect 185414 213120 188670 217728
rect 189450 215879 252914 217728
rect 189450 213120 216914 215879
rect 185414 211200 216914 213120
rect 185414 193536 193086 211200
rect 193866 207900 216914 211200
rect 217694 207900 220634 215879
rect 193866 196068 220634 207900
rect 193866 193536 216914 196068
rect 185414 174208 216914 193536
rect 185414 161984 188302 174208
rect 189082 173313 216914 174208
rect 217694 173313 220634 196068
rect 221414 211200 252914 215879
rect 221414 208480 223078 211200
rect 221414 195168 221422 208480
rect 222202 195168 223078 208480
rect 221414 193536 223078 195168
rect 223858 208480 252914 211200
rect 223858 195168 225286 208480
rect 226066 195168 252914 208480
rect 223858 193536 252914 195168
rect 221414 173313 252914 193536
rect 189082 161984 252914 173313
rect 185414 154624 252914 161984
rect 185414 150016 188670 154624
rect 189450 153079 252914 154624
rect 189450 150016 216914 153079
rect 185414 148096 216914 150016
rect 185414 130432 193086 148096
rect 193866 145100 216914 148096
rect 217694 145100 220634 153079
rect 193866 133268 220634 145100
rect 193866 130432 216914 133268
rect 185414 115456 216914 130432
rect 185414 113024 188302 115456
rect 189082 113024 216914 115456
rect 185414 112192 216914 113024
rect 185414 109760 188302 112192
rect 189082 110513 216914 112192
rect 217694 110513 220634 133268
rect 221414 148096 252914 153079
rect 221414 130432 223078 148096
rect 223858 130432 252914 148096
rect 221414 110513 252914 130432
rect 189082 109760 252914 110513
rect 185414 108928 252914 109760
rect 185414 106496 188302 108928
rect 189082 106496 252914 108928
rect 185414 92608 252914 106496
rect 185414 88000 188670 92608
rect 189450 90279 252914 92608
rect 189450 88000 216914 90279
rect 185414 84992 216914 88000
rect 185414 67328 193086 84992
rect 193866 82300 216914 84992
rect 217694 82300 220634 90279
rect 193866 70468 220634 82300
rect 193866 67328 216914 70468
rect 185414 51264 216914 67328
rect 185414 48992 203574 51264
rect 185414 33600 193086 48992
rect 193866 48832 203574 48992
rect 204354 48832 216914 51264
rect 193866 47900 216914 48832
rect 217694 47900 220634 70468
rect 193866 36068 220634 47900
rect 193866 33600 216914 36068
rect 185414 2928 216914 33600
rect 217694 2928 220634 36068
rect 221414 84992 252914 90279
rect 221414 67328 223078 84992
rect 223858 67328 252914 84992
rect 221414 50176 252914 67328
rect 221414 48544 223078 50176
rect 221414 35232 221422 48544
rect 222202 47744 223078 48544
rect 223858 48544 252914 50176
rect 223858 47744 225286 48544
rect 222202 46912 225286 47744
rect 222202 43392 223078 46912
rect 223858 43392 225286 46912
rect 222202 41472 225286 43392
rect 222202 37952 223078 41472
rect 223858 37952 225286 41472
rect 222202 36032 225286 37952
rect 222202 35232 223078 36032
rect 221414 33600 223078 35232
rect 223858 35232 225286 36032
rect 226066 35232 252914 48544
rect 223858 33600 252914 35232
rect 221414 2928 252914 33600
rect 253694 2928 256634 697752
rect 257414 675713 288914 697752
rect 289694 675713 292634 697752
rect 257414 655479 292634 675713
rect 257414 650208 288914 655479
rect 257414 632544 287110 650208
rect 287890 632544 288914 650208
rect 257414 612913 288914 632544
rect 289694 647177 292634 655479
rect 293414 688288 324914 697752
rect 293414 677696 314158 688288
rect 314938 677776 318022 688288
rect 318802 677776 324914 688288
rect 315306 677696 318022 677776
rect 293414 663808 314526 677696
rect 315306 663808 318390 677696
rect 293414 652672 314158 663808
rect 315306 663728 318022 663808
rect 319170 663728 324914 677776
rect 314938 652672 318022 663728
rect 318802 652672 324914 663728
rect 293414 647177 324914 652672
rect 289694 629255 324914 647177
rect 289694 612913 292634 629255
rect 257414 592679 292634 612913
rect 257414 586016 288914 592679
rect 257414 569440 287110 586016
rect 287890 569440 288914 586016
rect 257414 550113 288914 569440
rect 289694 590633 292634 592679
rect 293414 625728 324914 629255
rect 293414 614592 314158 625728
rect 314938 614672 318022 625728
rect 318802 614672 324914 625728
rect 315306 614592 318022 614672
rect 293414 600704 314526 614592
rect 315306 600704 318390 614592
rect 293414 592832 314158 600704
rect 315306 600624 318022 600704
rect 319170 600624 324914 614672
rect 314938 592912 318022 600624
rect 318802 592912 324914 600624
rect 315490 592832 318022 592912
rect 293414 590633 314710 592832
rect 289694 590112 314710 590633
rect 315490 590112 318574 592832
rect 319354 590112 324914 592912
rect 289694 567543 324914 590112
rect 289694 550113 292634 567543
rect 257414 529879 292634 550113
rect 257414 525088 288914 529879
rect 257414 507424 287110 525088
rect 287890 507424 288914 525088
rect 257414 487313 288914 507424
rect 289694 527833 292634 529879
rect 293414 563168 324914 567543
rect 293414 552032 314158 563168
rect 314938 552112 318022 563168
rect 318802 552112 324914 563168
rect 315306 552032 318022 552112
rect 293414 538144 314526 552032
rect 315306 538144 318390 552032
rect 293414 530272 314158 538144
rect 315306 538064 318022 538144
rect 319170 538064 324914 552112
rect 314938 530352 318022 538064
rect 318802 530352 324914 538064
rect 315490 530272 318022 530352
rect 293414 527833 314710 530272
rect 289694 527008 314710 527833
rect 315490 527008 318574 530272
rect 319354 527008 324914 530352
rect 289694 504743 324914 527008
rect 289694 487313 292634 504743
rect 257414 467079 292634 487313
rect 257414 461984 288914 467079
rect 257414 444320 287110 461984
rect 287890 444320 288914 461984
rect 257414 424513 288914 444320
rect 289694 465033 292634 467079
rect 293414 500064 324914 504743
rect 293414 489472 306798 500064
rect 307578 489472 310662 500064
rect 311442 491360 324914 500064
rect 311442 489472 314526 491360
rect 293414 475040 314526 489472
rect 315306 475040 318390 491360
rect 293414 467168 314158 475040
rect 315306 474960 318022 475040
rect 319170 474960 324914 491360
rect 314938 467248 318022 474960
rect 318802 467248 324914 474960
rect 315490 467168 318022 467248
rect 293414 465033 314710 467168
rect 289694 464448 314710 465033
rect 315490 464448 318574 467168
rect 319354 464448 324914 467248
rect 289694 442006 324914 464448
rect 289694 424513 292634 442006
rect 257414 404279 292634 424513
rect 257414 398880 288914 404279
rect 257414 381216 287110 398880
rect 287890 381216 288914 398880
rect 257414 361713 288914 381216
rect 289694 402233 292634 404279
rect 293414 437504 324914 442006
rect 293414 426368 314158 437504
rect 314938 426448 318022 437504
rect 318802 426448 324914 437504
rect 315306 426368 318022 426448
rect 293414 412480 314526 426368
rect 315306 412480 318390 426368
rect 293414 404608 314158 412480
rect 315306 412400 318022 412480
rect 319170 412400 324914 426448
rect 314938 404688 318022 412400
rect 318802 404688 324914 412400
rect 315490 404608 318022 404688
rect 293414 402233 314710 404608
rect 289694 401344 314710 402233
rect 315490 401344 318574 404608
rect 319354 401344 324914 404688
rect 289694 379143 324914 401344
rect 289694 361713 292634 379143
rect 257414 341479 292634 361713
rect 257414 335776 288914 341479
rect 257414 319200 287110 335776
rect 287890 319200 288914 335776
rect 257414 298913 288914 319200
rect 289694 339433 292634 341479
rect 293414 374400 324914 379143
rect 293414 363808 314158 374400
rect 314938 363888 318022 374400
rect 318802 363888 324914 374400
rect 315306 363808 318022 363888
rect 293414 349376 314526 363808
rect 315306 349376 318390 363808
rect 293414 341504 314158 349376
rect 315306 349296 318022 349376
rect 319170 349296 324914 363888
rect 314938 341584 318022 349296
rect 318802 341584 324914 349296
rect 315490 341504 318022 341584
rect 293414 339433 314710 341504
rect 289694 338784 314710 339433
rect 315490 338784 318574 341504
rect 319354 338784 324914 341584
rect 289694 316343 324914 338784
rect 289694 298913 292634 316343
rect 257414 278679 292634 298913
rect 257414 273760 288914 278679
rect 257414 256096 287110 273760
rect 287890 256096 288914 273760
rect 257414 236113 288914 256096
rect 289694 276633 292634 278679
rect 293414 311840 324914 316343
rect 293414 300704 314158 311840
rect 314938 300784 318022 311840
rect 318802 300784 324914 311840
rect 315306 300704 318022 300784
rect 293414 286816 314526 300704
rect 315306 286816 318390 300704
rect 293414 278944 314158 286816
rect 315306 286736 318022 286816
rect 319170 286736 324914 300784
rect 314938 279024 318022 286736
rect 318802 279024 324914 286736
rect 315490 278944 318022 279024
rect 293414 276633 314710 278944
rect 289694 275680 314710 276633
rect 315490 275680 318574 278944
rect 319354 275680 324914 279024
rect 289694 253543 324914 275680
rect 289694 236113 292634 253543
rect 257414 215879 292634 236113
rect 257414 210656 288914 215879
rect 257414 192992 287110 210656
rect 287890 192992 288914 210656
rect 257414 173313 288914 192992
rect 289694 213833 292634 215879
rect 293414 248736 324914 253543
rect 293414 238144 314158 248736
rect 314938 238224 318022 248736
rect 318802 238224 324914 248736
rect 315306 238144 318022 238224
rect 293414 223712 314526 238144
rect 315306 223712 318390 238144
rect 293414 215840 314158 223712
rect 315306 223632 318022 223712
rect 319170 223632 324914 238224
rect 314938 215920 318022 223632
rect 318802 215920 324914 223632
rect 315490 215840 318022 215920
rect 293414 213833 314710 215840
rect 289694 213120 314710 213833
rect 315490 213120 318574 215840
rect 319354 213120 324914 215920
rect 289694 190743 324914 213120
rect 289694 173313 292634 190743
rect 257414 153079 292634 173313
rect 257414 147552 288914 153079
rect 257414 130976 287110 147552
rect 287890 130976 288914 147552
rect 257414 110513 288914 130976
rect 289694 151033 292634 153079
rect 293414 186176 324914 190743
rect 293414 175040 314158 186176
rect 314938 175120 318022 186176
rect 318802 175120 324914 186176
rect 315306 175040 318022 175120
rect 293414 161152 314526 175040
rect 315306 161152 318390 175040
rect 293414 153280 314158 161152
rect 315306 161072 318022 161152
rect 319170 161072 324914 175120
rect 314938 153360 318022 161072
rect 318802 153360 324914 161072
rect 315490 153280 318022 153360
rect 293414 151033 314710 153280
rect 289694 150016 314710 151033
rect 315490 150016 318574 153280
rect 319354 150016 324914 153360
rect 289694 127943 324914 150016
rect 289694 110513 292634 127943
rect 257414 90279 292634 110513
rect 257414 85536 288914 90279
rect 257414 67872 287110 85536
rect 287890 67872 288914 85536
rect 257414 50720 288914 67872
rect 257414 33056 287110 50720
rect 287890 33056 288914 50720
rect 257414 2928 288914 33056
rect 289694 88233 292634 90279
rect 293414 123072 324914 127943
rect 293414 119008 314158 123072
rect 314938 119088 318022 123072
rect 318802 119088 324914 123072
rect 315306 119008 318022 119088
rect 293414 105120 314526 119008
rect 315306 105120 318390 119008
rect 293414 90720 314158 105120
rect 315306 105040 318022 105120
rect 319170 105040 324914 119088
rect 314938 90800 318022 105040
rect 318802 90800 324914 105040
rect 315490 90720 318022 90800
rect 293414 88233 314710 90720
rect 289694 87456 314710 88233
rect 315490 87456 318574 90720
rect 319354 87456 324914 90800
rect 289694 65143 324914 87456
rect 289694 2928 292634 65143
rect 293414 2928 324914 65143
rect 325694 675713 328634 697752
rect 329414 676500 360914 697752
rect 361694 676500 364634 697752
rect 365414 679584 396914 697752
rect 365414 676500 378374 679584
rect 329414 675713 378374 676500
rect 325694 664668 378374 675713
rect 325694 655479 360914 664668
rect 325694 612913 328634 655479
rect 329414 650752 360914 655479
rect 329414 632544 349302 650752
rect 350082 632544 353166 650752
rect 353946 647177 360914 650752
rect 361694 647177 364634 664668
rect 365414 663808 378374 664668
rect 379154 663808 382238 679584
rect 383018 675713 396914 679584
rect 397694 676500 432914 697752
rect 433694 676500 436634 697752
rect 397694 675713 436634 676500
rect 383018 664668 436634 675713
rect 365414 661376 378190 663808
rect 379154 663728 382054 663808
rect 383018 663728 432914 664668
rect 378970 661376 382054 663728
rect 382834 661376 432914 663728
rect 365414 655479 432914 661376
rect 365414 650752 396914 655479
rect 365414 647177 383342 650752
rect 353946 632544 383342 647177
rect 384122 632544 387206 650752
rect 387986 632544 396914 650752
rect 329414 629255 396914 632544
rect 329414 613700 360914 629255
rect 361694 613700 364634 629255
rect 365414 617024 396914 629255
rect 365414 614592 378190 617024
rect 378970 614672 382054 617024
rect 382834 614672 396914 617024
rect 379154 614592 382054 614672
rect 365414 613700 378374 614592
rect 329414 612913 378374 613700
rect 325694 601868 378374 612913
rect 325694 592679 360914 601868
rect 325694 550113 328634 592679
rect 329414 590633 360914 592679
rect 361694 590633 364634 601868
rect 365414 598816 378374 601868
rect 379154 598816 382238 614592
rect 383018 612913 396914 614672
rect 397694 647500 400634 655479
rect 401414 650752 432914 655479
rect 401414 647500 413334 650752
rect 397694 635668 413334 647500
rect 397694 622652 400634 635668
rect 401414 632544 413334 635668
rect 414114 632544 417198 650752
rect 417978 650116 432914 650752
rect 433694 650116 436634 664668
rect 417978 632544 436634 650116
rect 401414 629255 436634 632544
rect 401414 622652 432914 629255
rect 397694 613700 432914 622652
rect 433694 613700 436634 629255
rect 397694 612913 436634 613700
rect 383018 601868 436634 612913
rect 383018 598816 432914 601868
rect 365414 594720 432914 598816
rect 365414 590633 378742 594720
rect 329414 590112 378742 590633
rect 379522 590112 382606 594720
rect 383386 592679 432914 594720
rect 383386 590112 396914 592679
rect 329414 586560 396914 590112
rect 329414 568896 349302 586560
rect 350082 568896 353166 586560
rect 353946 570784 383342 586560
rect 384122 570784 387206 586560
rect 353946 568896 382790 570784
rect 384122 570704 386654 570784
rect 387986 570704 396914 586560
rect 329414 568352 382790 568896
rect 383570 568352 386654 570704
rect 387434 568352 396914 570704
rect 329414 567543 396914 568352
rect 329414 550900 360914 567543
rect 361694 550900 364634 567543
rect 365414 553920 396914 567543
rect 365414 550900 378374 553920
rect 329414 550113 378374 550900
rect 325694 539068 378374 550113
rect 325694 529879 360914 539068
rect 325694 487313 328634 529879
rect 329414 527833 360914 529879
rect 361694 527833 364634 539068
rect 365414 538144 378374 539068
rect 379154 538144 382238 553920
rect 383018 550113 396914 553920
rect 397694 583500 400634 592679
rect 401414 591668 432914 592679
rect 433694 591668 436634 601868
rect 401414 586560 436634 591668
rect 401414 583500 413334 586560
rect 397694 570624 413334 583500
rect 414114 571872 417198 586560
rect 414114 570624 414806 571872
rect 397694 569847 414806 570624
rect 397694 559852 400634 569847
rect 401414 568896 414806 569847
rect 416322 570624 417198 571872
rect 417978 570624 436634 586560
rect 416322 568896 436634 570624
rect 401414 567543 436634 568896
rect 401414 559852 432914 567543
rect 397694 550900 432914 559852
rect 433694 550900 436634 567543
rect 397694 550113 436634 550900
rect 383018 539068 436634 550113
rect 365414 535712 378190 538144
rect 379154 538064 382054 538144
rect 383018 538064 432914 539068
rect 378970 535712 382054 538064
rect 382834 535712 432914 538064
rect 365414 532160 432914 535712
rect 365414 527833 378742 532160
rect 329414 527008 378742 527833
rect 379522 527008 382606 532160
rect 383386 529879 432914 532160
rect 383386 527008 396914 529879
rect 329414 525088 396914 527008
rect 329414 506880 349302 525088
rect 350082 506880 353166 525088
rect 353946 506880 383342 525088
rect 384122 506880 387206 525088
rect 387986 506880 396914 525088
rect 329414 504743 396914 506880
rect 329414 488100 360914 504743
rect 361694 488100 364634 504743
rect 365414 491360 396914 504743
rect 365414 488100 378374 491360
rect 329414 487313 378374 488100
rect 325694 476268 378374 487313
rect 325694 467079 360914 476268
rect 325694 424513 328634 467079
rect 329414 465033 360914 467079
rect 361694 465033 364634 476268
rect 365414 473152 378374 476268
rect 379154 473152 382238 491360
rect 383018 487313 396914 491360
rect 397694 521900 400634 529879
rect 401414 528868 432914 529879
rect 433694 528868 436634 539068
rect 401414 525088 436634 528868
rect 401414 521900 413334 525088
rect 397694 508247 413334 521900
rect 397694 497052 400634 508247
rect 401414 506880 413334 508247
rect 414114 506880 417198 525088
rect 417978 506880 436634 525088
rect 401414 504743 436634 506880
rect 401414 497052 432914 504743
rect 397694 488100 432914 497052
rect 433694 488100 436634 504743
rect 397694 487313 436634 488100
rect 383018 476268 436634 487313
rect 383018 473152 432914 476268
rect 365414 469056 432914 473152
rect 365414 465033 378742 469056
rect 329414 464448 378742 465033
rect 379522 464448 382606 469056
rect 383386 467079 432914 469056
rect 383386 464448 396914 467079
rect 329414 461984 396914 464448
rect 329414 444320 349302 461984
rect 350082 444320 353166 461984
rect 353946 444320 383342 461984
rect 384122 444320 387206 461984
rect 387986 444320 396914 461984
rect 329414 442006 396914 444320
rect 329414 441943 364634 442006
rect 329414 425300 360914 441943
rect 361694 425300 364634 441943
rect 365414 428256 396914 442006
rect 365414 425300 378374 428256
rect 329414 424513 378374 425300
rect 325694 413468 378374 424513
rect 325694 404279 360914 413468
rect 325694 361713 328634 404279
rect 329414 402233 360914 404279
rect 361694 402233 364634 413468
rect 365414 410592 378374 413468
rect 379154 410592 382238 428256
rect 383018 424513 396914 428256
rect 397694 459100 400634 467079
rect 401414 466068 432914 467079
rect 433694 466068 436634 476268
rect 401414 461984 436634 466068
rect 401414 459100 413334 461984
rect 397694 445447 413334 459100
rect 397694 434252 400634 445447
rect 401414 444320 413334 445447
rect 414114 444320 417198 461984
rect 417978 444320 436634 461984
rect 401414 441943 436634 444320
rect 401414 434252 432914 441943
rect 397694 425300 432914 434252
rect 433694 425300 436634 441943
rect 397694 424513 436634 425300
rect 383018 413468 436634 424513
rect 383018 410592 432914 413468
rect 365414 406496 432914 410592
rect 365414 402233 378742 406496
rect 329414 401344 378742 402233
rect 379522 401344 382606 406496
rect 383386 404279 432914 406496
rect 383386 401344 396914 404279
rect 329414 399424 396914 401344
rect 329414 381216 349302 399424
rect 350082 381216 353166 399424
rect 353946 381216 383342 399424
rect 384122 381216 387206 399424
rect 387986 381216 396914 399424
rect 329414 379143 396914 381216
rect 329414 362500 360914 379143
rect 361694 362500 364634 379143
rect 365414 365696 396914 379143
rect 365414 362500 378374 365696
rect 329414 361713 378374 362500
rect 325694 350668 378374 361713
rect 325694 341479 360914 350668
rect 325694 298913 328634 341479
rect 329414 339433 360914 341479
rect 361694 339433 364634 350668
rect 365414 347488 378374 350668
rect 379154 347488 382238 365696
rect 383018 361713 396914 365696
rect 397694 396300 400634 404279
rect 401414 403268 432914 404279
rect 433694 403268 436634 413468
rect 401414 399424 436634 403268
rect 401414 396300 413334 399424
rect 397694 382647 413334 396300
rect 397694 371452 400634 382647
rect 401414 381216 413334 382647
rect 414114 381216 417198 399424
rect 417978 381216 436634 399424
rect 401414 379143 436634 381216
rect 401414 371452 432914 379143
rect 397694 362500 432914 371452
rect 433694 362500 436634 379143
rect 397694 361713 436634 362500
rect 383018 350668 436634 361713
rect 383018 347488 432914 350668
rect 365414 343392 432914 347488
rect 365414 339433 378742 343392
rect 329414 338784 378742 339433
rect 379522 338784 382606 343392
rect 383386 341479 432914 343392
rect 383386 338784 396914 341479
rect 329414 336864 396914 338784
rect 329414 336320 377270 336864
rect 329414 318656 349302 336320
rect 350082 318656 353166 336320
rect 353946 334432 377270 336320
rect 378050 334432 381134 336864
rect 381914 334592 396914 336864
rect 381914 334432 383342 334592
rect 353946 318656 383342 334432
rect 384122 318656 387206 334592
rect 387986 318656 396914 334592
rect 329414 316343 396914 318656
rect 329414 299700 360914 316343
rect 361694 299700 364634 316343
rect 365414 302592 396914 316343
rect 365414 299700 378374 302592
rect 329414 298913 378374 299700
rect 325694 287868 378374 298913
rect 325694 278679 360914 287868
rect 325694 236113 328634 278679
rect 329414 276633 360914 278679
rect 361694 276633 364634 287868
rect 365414 284928 378374 287868
rect 379154 284928 382238 302592
rect 383018 298913 396914 302592
rect 397694 333500 400634 341479
rect 401414 340468 432914 341479
rect 433694 340468 436634 350668
rect 401414 336320 436634 340468
rect 401414 334592 414806 336320
rect 401414 333500 413334 334592
rect 397694 319847 413334 333500
rect 397694 308652 400634 319847
rect 401414 318656 413334 319847
rect 414114 333344 414806 334592
rect 416322 334592 436634 336320
rect 416322 333344 417198 334592
rect 414114 318656 417198 333344
rect 417978 318656 436634 334592
rect 401414 316343 436634 318656
rect 401414 308652 432914 316343
rect 397694 299700 432914 308652
rect 433694 299700 436634 316343
rect 397694 298913 436634 299700
rect 383018 287868 436634 298913
rect 383018 284928 432914 287868
rect 365414 280832 432914 284928
rect 365414 276633 378742 280832
rect 329414 275680 378742 276633
rect 379522 275680 382606 280832
rect 383386 278679 432914 280832
rect 383386 275680 396914 278679
rect 329414 273760 396914 275680
rect 329414 256096 349302 273760
rect 350082 256096 353166 273760
rect 353946 256096 383342 273760
rect 384122 256096 387206 273760
rect 387986 256096 396914 273760
rect 329414 253543 396914 256096
rect 329414 236900 360914 253543
rect 361694 236900 364634 253543
rect 365414 240032 396914 253543
rect 365414 236900 378374 240032
rect 329414 236113 378374 236900
rect 325694 225068 378374 236113
rect 325694 215879 360914 225068
rect 325694 173313 328634 215879
rect 329414 213833 360914 215879
rect 361694 213833 364634 225068
rect 365414 221824 378374 225068
rect 379154 221824 382238 240032
rect 383018 236113 396914 240032
rect 397694 270700 400634 278679
rect 401414 277668 432914 278679
rect 433694 277668 436634 287868
rect 401414 273760 436634 277668
rect 401414 270700 413334 273760
rect 397694 257047 413334 270700
rect 397694 245852 400634 257047
rect 401414 256096 413334 257047
rect 414114 256096 417198 273760
rect 417978 256096 436634 273760
rect 401414 253543 436634 256096
rect 401414 245852 432914 253543
rect 397694 236900 432914 245852
rect 433694 236900 436634 253543
rect 397694 236113 436634 236900
rect 383018 225068 436634 236113
rect 383018 221824 432914 225068
rect 365414 218272 432914 221824
rect 365414 215840 378190 218272
rect 378970 215920 382054 218272
rect 382834 215920 432914 218272
rect 379522 215840 382054 215920
rect 383386 215879 432914 215920
rect 365414 213833 378742 215840
rect 329414 213120 378742 213833
rect 379522 213120 382606 215840
rect 383386 213120 396914 215879
rect 329414 211200 396914 213120
rect 329414 192992 349302 211200
rect 350082 192992 353166 211200
rect 353946 192992 383342 211200
rect 384122 192992 387206 211200
rect 387986 192992 396914 211200
rect 329414 190743 396914 192992
rect 329414 174100 360914 190743
rect 361694 174100 364634 190743
rect 365414 177472 396914 190743
rect 365414 175040 378190 177472
rect 378970 175120 382054 177472
rect 382834 175120 396914 177472
rect 379154 175040 382054 175120
rect 365414 174100 378374 175040
rect 329414 173313 378374 174100
rect 325694 162268 378374 173313
rect 325694 153079 360914 162268
rect 325694 110513 328634 153079
rect 329414 151033 360914 153079
rect 361694 151033 364634 162268
rect 365414 159264 378374 162268
rect 379154 159264 382238 175040
rect 383018 173313 396914 175120
rect 397694 207900 400634 215879
rect 401414 214868 432914 215879
rect 433694 214868 436634 225068
rect 401414 211200 436634 214868
rect 401414 207900 413334 211200
rect 397694 194247 413334 207900
rect 397694 183052 400634 194247
rect 401414 192992 413334 194247
rect 414114 192992 417198 211200
rect 417978 192992 436634 211200
rect 401414 190743 436634 192992
rect 401414 183052 432914 190743
rect 397694 174100 432914 183052
rect 433694 174100 436634 190743
rect 397694 173313 436634 174100
rect 383018 162268 436634 173313
rect 383018 159264 432914 162268
rect 365414 155168 432914 159264
rect 365414 151033 378742 155168
rect 329414 150016 378742 151033
rect 379522 150016 382606 155168
rect 383386 153079 432914 155168
rect 383386 150016 396914 153079
rect 329414 148096 396914 150016
rect 329414 130432 349302 148096
rect 350082 130432 353166 148096
rect 353946 130432 383342 148096
rect 384122 130432 387206 148096
rect 387986 130432 396914 148096
rect 329414 127943 396914 130432
rect 329414 117900 360914 127943
rect 361694 117900 364634 127943
rect 365414 120896 396914 127943
rect 365414 117900 378374 120896
rect 329414 110513 378374 117900
rect 325694 106068 378374 110513
rect 325694 90279 360914 106068
rect 325694 2928 328634 90279
rect 329414 88233 360914 90279
rect 361694 88233 364634 106068
rect 365414 103232 378374 106068
rect 379154 103232 382238 120896
rect 383018 110513 396914 120896
rect 397694 145100 400634 153079
rect 401414 152068 432914 153079
rect 433694 152068 436634 162268
rect 401414 148096 436634 152068
rect 401414 145100 413334 148096
rect 397694 131447 413334 145100
rect 397694 120252 400634 131447
rect 401414 130432 413334 131447
rect 414114 130432 417198 148096
rect 417978 130432 436634 148096
rect 401414 127943 436634 130432
rect 401414 120252 432914 127943
rect 397694 117900 432914 120252
rect 433694 117900 436634 127943
rect 397694 110513 436634 117900
rect 383018 106068 436634 110513
rect 383018 103232 432914 106068
rect 365414 92608 432914 103232
rect 365414 88233 378742 92608
rect 329414 87456 378742 88233
rect 379522 87456 382606 92608
rect 383386 90279 432914 92608
rect 383386 87456 396914 90279
rect 329414 85536 396914 87456
rect 329414 67328 349302 85536
rect 350082 67328 353166 85536
rect 353946 67328 383342 85536
rect 384122 67328 387206 85536
rect 387986 67328 396914 85536
rect 329414 65143 396914 67328
rect 329414 50720 360914 65143
rect 329414 33056 349302 50720
rect 350082 33056 353166 50720
rect 353946 33056 360914 50720
rect 329414 2928 360914 33056
rect 361694 2928 364634 65143
rect 365414 50720 396914 65143
rect 365414 33056 383342 50720
rect 384122 33056 387206 50720
rect 387986 33056 396914 50720
rect 365414 2928 396914 33056
rect 397694 82300 400634 90279
rect 401414 89268 432914 90279
rect 433694 89268 436634 106068
rect 401414 85536 436634 89268
rect 401414 82300 413334 85536
rect 397694 68647 413334 82300
rect 397694 47900 400634 68647
rect 401414 67328 413334 68647
rect 414114 67328 417198 85536
rect 417978 67328 436634 85536
rect 401414 65143 436634 67328
rect 401414 55516 432914 65143
rect 433694 55516 436634 65143
rect 401414 50720 436634 55516
rect 401414 47900 413334 50720
rect 397694 36068 413334 47900
rect 397694 2928 400634 36068
rect 401414 33056 413334 36068
rect 414114 33056 417198 50720
rect 417978 36068 436634 50720
rect 417978 33056 432914 36068
rect 401414 2928 432914 33056
rect 433694 2928 436634 36068
rect 437414 685452 468914 697752
rect 469694 685452 472634 697752
rect 473414 685452 504914 697752
rect 437414 679584 504914 685452
rect 437414 663808 442406 679584
rect 443186 663808 446270 679584
rect 437414 661376 442222 663808
rect 443186 663728 446086 663808
rect 447050 663728 504914 679584
rect 443002 661376 446086 663728
rect 446866 661376 504914 663728
rect 437414 655479 504914 661376
rect 437414 650752 468914 655479
rect 437414 632544 447190 650752
rect 447970 632544 451054 650752
rect 451834 647500 468914 650752
rect 469694 647500 472634 655479
rect 473414 650752 504914 655479
rect 473414 647500 477182 650752
rect 451834 635668 477182 647500
rect 451834 632544 468914 635668
rect 437414 622652 468914 632544
rect 469694 622652 472634 635668
rect 473414 632544 477182 635668
rect 477962 632544 481046 650752
rect 481826 632544 504914 650752
rect 473414 622652 504914 632544
rect 437414 617024 504914 622652
rect 437414 614592 442222 617024
rect 443002 614672 446086 617024
rect 446866 614672 504914 617024
rect 443186 614592 446086 614672
rect 437414 598816 442406 614592
rect 443186 598816 446270 614592
rect 447050 598816 504914 614672
rect 437414 594720 504914 598816
rect 437414 590112 442774 594720
rect 443554 590112 446638 594720
rect 447418 592679 504914 594720
rect 447418 590112 468914 592679
rect 437414 586560 468914 590112
rect 437414 568896 447190 586560
rect 447970 568896 451054 586560
rect 451834 583500 468914 586560
rect 469694 583500 472634 592679
rect 473414 586560 504914 592679
rect 473414 583500 477182 586560
rect 451834 571668 477182 583500
rect 451834 568896 468914 571668
rect 437414 559852 468914 568896
rect 469694 559852 472634 571668
rect 473414 568896 477182 571668
rect 477962 568896 481046 586560
rect 481826 568896 504914 586560
rect 473414 559852 504914 568896
rect 437414 553920 504914 559852
rect 437414 536256 442406 553920
rect 443186 536256 446270 553920
rect 447050 536256 504914 553920
rect 437414 532160 504914 536256
rect 437414 527008 442774 532160
rect 443554 527008 446638 532160
rect 447418 529879 504914 532160
rect 447418 527008 468914 529879
rect 437414 525088 468914 527008
rect 437414 506880 447190 525088
rect 447970 506880 451054 525088
rect 451834 521900 468914 525088
rect 469694 521900 472634 529879
rect 473414 525088 504914 529879
rect 473414 521900 477182 525088
rect 451834 510068 477182 521900
rect 451834 506880 468914 510068
rect 437414 497052 468914 506880
rect 469694 497052 472634 510068
rect 473414 506880 477182 510068
rect 477962 506880 481046 525088
rect 481826 506880 504914 525088
rect 473414 497052 504914 506880
rect 437414 491360 504914 497052
rect 437414 473152 442406 491360
rect 443186 473152 446270 491360
rect 447050 473152 504914 491360
rect 437414 469056 504914 473152
rect 437414 464448 442774 469056
rect 443554 464448 446638 469056
rect 447418 467079 504914 469056
rect 447418 464448 468914 467079
rect 437414 461984 468914 464448
rect 437414 444320 447190 461984
rect 447970 444320 451054 461984
rect 451834 459100 468914 461984
rect 469694 459100 472634 467079
rect 473414 461984 504914 467079
rect 473414 459100 477182 461984
rect 451834 447268 477182 459100
rect 451834 444320 468914 447268
rect 437414 434252 468914 444320
rect 469694 434252 472634 447268
rect 473414 444320 477182 447268
rect 477962 444320 481046 461984
rect 481826 444320 504914 461984
rect 473414 434252 504914 444320
rect 437414 428256 504914 434252
rect 437414 410592 442406 428256
rect 443186 410592 446270 428256
rect 447050 410592 504914 428256
rect 437414 406496 504914 410592
rect 437414 401344 442774 406496
rect 443554 401344 446638 406496
rect 447418 404279 504914 406496
rect 447418 401344 468914 404279
rect 437414 399424 468914 401344
rect 437414 381216 447190 399424
rect 447970 381216 451054 399424
rect 451834 396300 468914 399424
rect 469694 396300 472634 404279
rect 473414 399424 504914 404279
rect 473414 396300 477182 399424
rect 451834 384468 477182 396300
rect 451834 381216 468914 384468
rect 437414 371452 468914 381216
rect 469694 371452 472634 384468
rect 473414 381216 477182 384468
rect 477962 381216 481046 399424
rect 481826 381216 504914 399424
rect 473414 371452 504914 381216
rect 437414 365696 504914 371452
rect 437414 347488 442406 365696
rect 443186 347488 446270 365696
rect 447050 347488 504914 365696
rect 437414 343392 504914 347488
rect 437414 338784 442774 343392
rect 443554 338784 446638 343392
rect 447418 341479 504914 343392
rect 447418 338784 468914 341479
rect 437414 336864 468914 338784
rect 437414 334432 441302 336864
rect 442082 334432 445166 336864
rect 445946 334592 468914 336864
rect 445946 334432 447190 334592
rect 437414 318656 447190 334432
rect 447970 318656 451054 334592
rect 451834 333500 468914 334592
rect 469694 333500 472634 341479
rect 473414 336320 504914 341479
rect 473414 334592 478838 336320
rect 473414 333500 477182 334592
rect 451834 321668 477182 333500
rect 451834 318656 468914 321668
rect 437414 308652 468914 318656
rect 469694 308652 472634 321668
rect 473414 318656 477182 321668
rect 477962 333344 478838 334592
rect 480354 334592 504914 336320
rect 480354 333344 481046 334592
rect 477962 318656 481046 333344
rect 481826 318656 504914 334592
rect 473414 308652 504914 318656
rect 437414 302592 504914 308652
rect 437414 284928 442406 302592
rect 443186 284928 446270 302592
rect 447050 284928 504914 302592
rect 437414 280832 504914 284928
rect 437414 275680 442774 280832
rect 443554 275680 446638 280832
rect 447418 278679 504914 280832
rect 447418 275680 468914 278679
rect 437414 273760 468914 275680
rect 437414 256096 447190 273760
rect 447970 256096 451054 273760
rect 451834 270700 468914 273760
rect 469694 270700 472634 278679
rect 473414 273760 504914 278679
rect 473414 270700 477182 273760
rect 451834 258868 477182 270700
rect 451834 256096 468914 258868
rect 437414 245852 468914 256096
rect 469694 245852 472634 258868
rect 473414 256096 477182 258868
rect 477962 256096 481046 273760
rect 481826 256096 504914 273760
rect 473414 245852 504914 256096
rect 437414 240032 504914 245852
rect 437414 221824 442406 240032
rect 443186 221824 446270 240032
rect 447050 221824 504914 240032
rect 437414 217728 504914 221824
rect 437414 213120 442774 217728
rect 443554 213120 446638 217728
rect 447418 215879 504914 217728
rect 447418 213120 468914 215879
rect 437414 211200 468914 213120
rect 437414 192992 447190 211200
rect 447970 192992 451054 211200
rect 451834 207900 468914 211200
rect 469694 207900 472634 215879
rect 473414 211200 504914 215879
rect 473414 207900 477182 211200
rect 451834 196068 477182 207900
rect 451834 192992 468914 196068
rect 437414 183052 468914 192992
rect 469694 183052 472634 196068
rect 473414 192992 477182 196068
rect 477962 192992 481046 211200
rect 481826 192992 504914 211200
rect 473414 183052 504914 192992
rect 437414 177472 504914 183052
rect 437414 175040 437622 177472
rect 438402 175040 441486 177472
rect 442266 175200 504914 177472
rect 442266 175040 442406 175200
rect 437414 159264 442406 175040
rect 443186 159264 446270 175200
rect 447050 159264 504914 175200
rect 437414 155168 504914 159264
rect 437414 150016 442774 155168
rect 443554 150016 446638 155168
rect 447418 153079 504914 155168
rect 447418 150016 468914 153079
rect 437414 148096 468914 150016
rect 437414 130432 447190 148096
rect 447970 130432 451054 148096
rect 451834 145100 468914 148096
rect 469694 145100 472634 153079
rect 473414 148096 504914 153079
rect 473414 145100 477182 148096
rect 451834 133268 477182 145100
rect 451834 130432 468914 133268
rect 437414 120896 468914 130432
rect 437414 103232 442406 120896
rect 443186 103232 446270 120896
rect 447050 120252 468914 120896
rect 469694 120252 472634 133268
rect 473414 130432 477182 133268
rect 477962 130432 481046 148096
rect 481826 130432 504914 148096
rect 473414 120252 504914 130432
rect 447050 103232 504914 120252
rect 437414 92608 504914 103232
rect 437414 87456 442774 92608
rect 443554 87456 446638 92608
rect 447418 90279 504914 92608
rect 447418 87456 468914 90279
rect 437414 85536 468914 87456
rect 437414 67328 447190 85536
rect 447970 67328 451054 85536
rect 451834 82300 468914 85536
rect 469694 82300 472634 90279
rect 473414 85536 504914 90279
rect 473414 82300 477182 85536
rect 451834 70468 477182 82300
rect 451834 67328 468914 70468
rect 437414 50720 468914 67328
rect 437414 33056 447190 50720
rect 447970 33056 451054 50720
rect 451834 47900 468914 50720
rect 469694 47900 472634 70468
rect 473414 67328 477182 70468
rect 477962 67328 481046 85536
rect 481826 67328 504914 85536
rect 473414 50720 504914 67328
rect 473414 47900 477182 50720
rect 451834 36068 477182 47900
rect 451834 33056 468914 36068
rect 437414 12700 468914 33056
rect 469694 12700 472634 36068
rect 437414 2928 472634 12700
rect 473414 33056 477182 36068
rect 477962 33056 481046 50720
rect 481826 33056 504914 50720
rect 473414 2928 504914 33056
rect 505694 2928 508634 697752
rect 509414 675713 540914 697752
rect 541694 675713 544634 697752
rect 545414 675713 576035 697752
rect 509414 674688 576035 675713
rect 509414 663808 566422 674688
rect 509414 655479 565870 663808
rect 567938 663728 576035 674688
rect 509414 612913 540914 655479
rect 541694 612913 544634 655479
rect 545414 652672 565870 655479
rect 567386 652672 576035 663728
rect 545414 612913 576035 652672
rect 509414 611584 576035 612913
rect 509414 600704 566422 611584
rect 509414 592679 565870 600704
rect 567938 600624 576035 611584
rect 509414 550113 540914 592679
rect 541694 550113 544634 592679
rect 545414 590112 565870 592679
rect 567386 590112 576035 600624
rect 545414 550113 576035 590112
rect 509414 549024 576035 550113
rect 509414 538144 566422 549024
rect 509414 529879 565870 538144
rect 567938 538064 576035 549024
rect 509414 487313 540914 529879
rect 541694 522368 544634 529879
rect 541694 509056 543054 522368
rect 543834 509056 544634 522368
rect 541694 487313 544634 509056
rect 545414 527008 565870 529879
rect 567386 527008 576035 538064
rect 545414 487313 576035 527008
rect 509414 485920 576035 487313
rect 509414 475040 567342 485920
rect 509414 467079 562006 475040
rect 509414 424513 540914 467079
rect 541694 424513 544634 467079
rect 545414 464448 562006 467079
rect 562786 464448 565870 475040
rect 566650 473696 567342 475040
rect 568858 473696 576035 485920
rect 566650 464448 576035 473696
rect 545414 424513 576035 464448
rect 509414 423360 576035 424513
rect 509414 412480 566422 423360
rect 509414 404279 565870 412480
rect 567938 412400 576035 423360
rect 509414 361713 540914 404279
rect 541694 361713 544634 404279
rect 545414 401344 565870 404279
rect 567386 401344 576035 412400
rect 545414 361713 576035 401344
rect 509414 360800 576035 361713
rect 509414 349376 567342 360800
rect 509414 341479 562006 349376
rect 509414 298913 540914 341479
rect 541694 334144 544634 341479
rect 541694 320832 543054 334144
rect 543834 320832 544634 334144
rect 541694 298913 544634 320832
rect 545414 338784 562006 341479
rect 562786 338784 565870 349376
rect 566650 347488 567342 349376
rect 568858 347488 576035 360800
rect 566650 338784 576035 347488
rect 545414 298913 576035 338784
rect 509414 297696 576035 298913
rect 509414 286816 566422 297696
rect 509414 278679 565870 286816
rect 567938 286736 576035 297696
rect 509414 236113 540914 278679
rect 541694 236113 544634 278679
rect 545414 275680 565870 278679
rect 567386 275680 576035 286736
rect 545414 236113 576035 275680
rect 509414 235136 576035 236113
rect 509414 223712 567342 235136
rect 509414 215879 562006 223712
rect 509414 173313 540914 215879
rect 541694 173313 544634 215879
rect 545414 213120 562006 215879
rect 562786 213120 565870 223712
rect 566650 222368 567342 223712
rect 568858 222368 576035 235136
rect 566650 213120 576035 222368
rect 545414 173313 576035 213120
rect 509414 172032 576035 173313
rect 509414 161152 566422 172032
rect 509414 153079 565870 161152
rect 567938 161072 576035 172032
rect 509414 110513 540914 153079
rect 541694 110513 544634 153079
rect 545414 150016 565870 153079
rect 567386 150016 576035 161072
rect 545414 110513 576035 150016
rect 509414 109472 576035 110513
rect 509414 105120 566422 109472
rect 509414 90279 565870 105120
rect 567938 105040 576035 109472
rect 509414 2928 540914 90279
rect 541694 82816 544634 90279
rect 541694 69504 543054 82816
rect 543834 69504 544634 82816
rect 541694 2928 544634 69504
rect 545414 87456 565870 90279
rect 567386 87456 576035 105040
rect 545414 2928 576035 87456
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 699306 592650 699926
rect -8726 698066 592650 698686
rect -8726 693306 592650 693926
rect -8726 692066 592650 692686
rect -8726 687306 592650 687926
rect -8726 686066 592650 686686
rect -8726 681306 592650 681926
rect -8726 680066 592650 680686
rect -8726 675306 592650 675926
rect -8726 674066 592650 674686
rect -8726 669306 592650 669926
rect -8726 668066 592650 668686
rect -8726 663306 592650 663926
rect -8726 662066 592650 662686
rect -8726 657306 592650 657926
rect -8726 656066 592650 656686
rect -8726 651306 592650 651926
rect -8726 650066 592650 650686
rect -8726 645306 592650 645926
rect -8726 644066 592650 644686
rect -8726 639306 592650 639926
rect -8726 638066 592650 638686
rect -8726 633306 592650 633926
rect -8726 632066 592650 632686
rect -8726 627306 592650 627926
rect -8726 626066 592650 626686
rect -8726 621306 592650 621926
rect -8726 620066 592650 620686
rect -8726 615306 592650 615926
rect -8726 614066 592650 614686
rect -8726 609306 592650 609926
rect -8726 608066 592650 608686
rect -8726 603306 592650 603926
rect -8726 602066 592650 602686
rect -8726 597306 592650 597926
rect -8726 596066 592650 596686
rect -8726 591306 592650 591926
rect -8726 590066 592650 590686
rect -8726 585306 592650 585926
rect -8726 584066 592650 584686
rect -8726 579306 592650 579926
rect -8726 578066 592650 578686
rect -8726 573306 592650 573926
rect -8726 572066 592650 572686
rect -8726 567306 592650 567926
rect -8726 566066 592650 566686
rect -8726 561306 592650 561926
rect -8726 560066 592650 560686
rect -8726 555306 592650 555926
rect -8726 554066 592650 554686
rect -8726 549306 592650 549926
rect -8726 548066 592650 548686
rect -8726 543306 592650 543926
rect -8726 542066 592650 542686
rect -8726 537306 592650 537926
rect -8726 536066 592650 536686
rect -8726 531306 592650 531926
rect -8726 530066 592650 530686
rect -8726 525306 592650 525926
rect -8726 524066 592650 524686
rect -8726 519306 592650 519926
rect -8726 518066 592650 518686
rect -8726 513306 592650 513926
rect -8726 512066 592650 512686
rect -8726 507306 592650 507926
rect -8726 506066 592650 506686
rect -8726 501306 592650 501926
rect -8726 500066 592650 500686
rect -8726 495306 592650 495926
rect -8726 494066 592650 494686
rect -8726 489306 592650 489926
rect -8726 488066 592650 488686
rect -8726 483306 592650 483926
rect -8726 482066 592650 482686
rect -8726 477306 592650 477926
rect -8726 476066 592650 476686
rect -8726 471306 592650 471926
rect -8726 470066 592650 470686
rect -8726 465306 592650 465926
rect -8726 464066 592650 464686
rect -8726 459306 592650 459926
rect -8726 458066 592650 458686
rect -8726 453306 592650 453926
rect -8726 452066 592650 452686
rect -8726 447306 592650 447926
rect -8726 446066 592650 446686
rect -8726 441306 592650 441926
rect -8726 440066 592650 440686
rect -8726 435306 592650 435926
rect -8726 434066 592650 434686
rect -8726 429306 592650 429926
rect -8726 428066 592650 428686
rect -8726 423306 592650 423926
rect -8726 422066 592650 422686
rect -8726 417306 592650 417926
rect -8726 416066 592650 416686
rect -8726 411306 592650 411926
rect -8726 410066 592650 410686
rect -8726 405306 592650 405926
rect -8726 404066 592650 404686
rect -8726 399306 592650 399926
rect -8726 398066 592650 398686
rect -8726 393306 592650 393926
rect -8726 392066 592650 392686
rect -8726 387306 592650 387926
rect -8726 386066 592650 386686
rect -8726 381306 592650 381926
rect -8726 380066 592650 380686
rect -8726 375306 592650 375926
rect -8726 374066 592650 374686
rect -8726 369306 592650 369926
rect -8726 368066 592650 368686
rect -8726 363306 592650 363926
rect -8726 362066 592650 362686
rect -8726 357306 592650 357926
rect -8726 356066 592650 356686
rect -8726 351306 592650 351926
rect -8726 350066 592650 350686
rect -8726 345306 592650 345926
rect -8726 344066 592650 344686
rect -8726 339306 592650 339926
rect -8726 338066 592650 338686
rect -8726 333306 592650 333926
rect -8726 332066 592650 332686
rect -8726 327306 592650 327926
rect -8726 326066 592650 326686
rect -8726 321306 592650 321926
rect -8726 320066 592650 320686
rect -8726 315306 592650 315926
rect -8726 314066 592650 314686
rect -8726 309306 592650 309926
rect -8726 308066 592650 308686
rect -8726 303306 592650 303926
rect -8726 302066 592650 302686
rect -8726 297306 592650 297926
rect -8726 296066 592650 296686
rect -8726 291306 592650 291926
rect -8726 290066 592650 290686
rect -8726 285306 592650 285926
rect -8726 284066 592650 284686
rect -8726 279306 592650 279926
rect -8726 278066 592650 278686
rect -8726 273306 592650 273926
rect -8726 272066 592650 272686
rect -8726 267306 592650 267926
rect -8726 266066 592650 266686
rect -8726 261306 592650 261926
rect -8726 260066 592650 260686
rect -8726 255306 592650 255926
rect -8726 254066 592650 254686
rect -8726 249306 592650 249926
rect -8726 248066 592650 248686
rect -8726 243306 592650 243926
rect -8726 242066 592650 242686
rect -8726 237306 592650 237926
rect -8726 236066 592650 236686
rect -8726 231306 592650 231926
rect -8726 230066 592650 230686
rect -8726 225306 592650 225926
rect -8726 224066 592650 224686
rect -8726 219306 592650 219926
rect -8726 218066 592650 218686
rect -8726 213306 592650 213926
rect -8726 212066 592650 212686
rect -8726 207306 592650 207926
rect -8726 206066 592650 206686
rect -8726 201306 592650 201926
rect -8726 200066 592650 200686
rect -8726 195306 592650 195926
rect -8726 194066 592650 194686
rect -8726 189306 592650 189926
rect -8726 188066 592650 188686
rect -8726 183306 592650 183926
rect -8726 182066 592650 182686
rect -8726 177306 592650 177926
rect -8726 176066 592650 176686
rect -8726 171306 592650 171926
rect -8726 170066 592650 170686
rect -8726 165306 592650 165926
rect -8726 164066 592650 164686
rect -8726 159306 592650 159926
rect -8726 158066 592650 158686
rect -8726 153306 592650 153926
rect -8726 152066 592650 152686
rect -8726 147306 592650 147926
rect -8726 146066 592650 146686
rect -8726 141306 592650 141926
rect -8726 140066 592650 140686
rect -8726 135306 592650 135926
rect -8726 134066 592650 134686
rect -8726 129306 592650 129926
rect -8726 128066 592650 128686
rect -8726 123306 592650 123926
rect -8726 122066 592650 122686
rect -8726 117306 592650 117926
rect -8726 116066 592650 116686
rect -8726 111306 592650 111926
rect -8726 110066 592650 110686
rect -8726 105306 592650 105926
rect -8726 104066 592650 104686
rect -8726 99306 592650 99926
rect -8726 98066 592650 98686
rect -8726 93306 592650 93926
rect -8726 92066 592650 92686
rect -8726 87306 592650 87926
rect -8726 86066 592650 86686
rect -8726 81306 592650 81926
rect -8726 80066 592650 80686
rect -8726 75306 592650 75926
rect -8726 74066 592650 74686
rect -8726 69306 592650 69926
rect -8726 68066 592650 68686
rect -8726 63306 592650 63926
rect -8726 62066 592650 62686
rect -8726 57306 592650 57926
rect -8726 56066 592650 56686
rect -8726 51306 592650 51926
rect -8726 50066 592650 50686
rect -8726 45306 592650 45926
rect -8726 44066 592650 44686
rect -8726 39306 592650 39926
rect -8726 38066 592650 38686
rect -8726 33306 592650 33926
rect -8726 32066 592650 32686
rect -8726 27306 592650 27926
rect -8726 26066 592650 26686
rect -8726 21306 592650 21926
rect -8726 20066 592650 20686
rect -8726 15306 592650 15926
rect -8726 14066 592650 14686
rect -8726 9306 592650 9926
rect -8726 8066 592650 8686
rect -8726 3306 592650 3926
rect -8726 2066 592650 2686
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 4714 -7654 5334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 -7654 41334 65388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 83364 41334 128188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 146164 41334 190988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 208964 41334 253788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 271764 41334 316588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 334564 41334 379388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 397364 41334 442188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 460164 41334 504988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 522964 41334 567788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 40714 585764 41334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 -7654 77334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 110593 77334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 173393 77334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 236193 77334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 298993 77334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 361793 77334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 424593 77334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 487393 77334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 550193 77334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 612993 77334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 76714 675793 77334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 -7654 113334 35988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 55596 113334 65063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 89348 113334 105988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 117980 113334 127863 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 152148 113334 162188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 174180 113334 190663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 214948 113334 224988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 236980 113334 253463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 277748 113334 287788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 299780 113334 316263 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 340548 113334 350588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 362580 113334 379063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 403348 113334 413388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 425380 113334 441926 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 466148 113334 476188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 488180 113334 504663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 528948 113334 538988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 550980 113334 567463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 591748 113334 601788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 613780 113334 629175 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 650196 113334 664588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 112714 676580 113334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 12780 149334 35988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 47980 149334 70388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 82380 149334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 120332 149334 133188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 145180 149334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 183132 149334 195988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 207980 149334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 245932 149334 258788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 270780 149334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 308732 149334 321588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 333580 149334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 371532 149334 384388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 396380 149334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 434332 149334 447188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 459180 149334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 497132 149334 509988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 521980 149334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 559932 149334 571588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 583580 149334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 622732 149334 635588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 647580 149334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 148714 685532 149334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 184714 -7654 185334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 -7654 221334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 110593 221334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 173393 221334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 236193 221334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 298993 221334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 361793 221334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 424593 221334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 487393 221334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 550193 221334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 612993 221334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 220714 675793 221334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 256714 -7654 257334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 -7654 293334 65063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 88313 293334 127863 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 151113 293334 190663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 213913 293334 253463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 276713 293334 316263 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 339513 293334 379063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 402313 293334 441926 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 465113 293334 504663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 527913 293334 567463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 590713 293334 629175 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 292714 647257 293334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 -7654 329334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 110593 329334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 173393 329334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 236193 329334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 298993 329334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 361793 329334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 424593 329334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 487393 329334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 550193 329334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 612993 329334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 328714 675793 329334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 -7654 365334 65063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 88313 365334 105988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 117980 365334 127863 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 151113 365334 162188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 174180 365334 190663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 213913 365334 224988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 236980 365334 253463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 276713 365334 287788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 299780 365334 316263 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 339513 365334 350588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 362580 365334 379063 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 402313 365334 413388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 425380 365334 441926 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 465113 365334 476188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 488180 365334 504663 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 527913 365334 538988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 550980 365334 567463 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 590713 365334 601788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 613780 365334 629175 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 647257 365334 664588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 364714 676580 365334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 -7654 401334 35988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 47980 401334 68567 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 82380 401334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 120332 401334 131367 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 145180 401334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 183132 401334 194167 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 207980 401334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 245932 401334 256967 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 270780 401334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 308732 401334 319767 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 333580 401334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 371532 401334 382567 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 396380 401334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 434332 401334 445367 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 459180 401334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 497132 401334 508167 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 521980 401334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 559932 401334 569767 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 583580 401334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 622732 401334 635588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 647580 401334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 400714 699892 401334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 436714 -7654 437334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 -7654 473334 35988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 47980 473334 70388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 82380 473334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 120332 473334 133188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 145180 473334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 183132 473334 195988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 207980 473334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 245932 473334 258788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 270780 473334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 308732 473334 321588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 333580 473334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 371532 473334 384388 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 396380 473334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 434332 473334 447188 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 459180 473334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 497132 473334 509988 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 521980 473334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 559932 473334 571588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 583580 473334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 622732 473334 635588 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 647580 473334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 472714 685532 473334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 508714 -7654 509334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 -7654 545334 90199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 110593 545334 152999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 173393 545334 215799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 236193 545334 278599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 298993 545334 341399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 361793 545334 404199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 424593 545334 466999 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 487393 545334 529799 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 550193 545334 592599 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 612993 545334 655399 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 544714 675793 545334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 580714 -7654 581334 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 3306 592650 3926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 9306 592650 9926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 15306 592650 15926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 21306 592650 21926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 27306 592650 27926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 33306 592650 33926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 39306 592650 39926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 45306 592650 45926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 51306 592650 51926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 57306 592650 57926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 63306 592650 63926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 69306 592650 69926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 75306 592650 75926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 81306 592650 81926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 87306 592650 87926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 93306 592650 93926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 99306 592650 99926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 105306 592650 105926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 111306 592650 111926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 117306 592650 117926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 123306 592650 123926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 129306 592650 129926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 135306 592650 135926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 141306 592650 141926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 147306 592650 147926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 153306 592650 153926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 159306 592650 159926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 165306 592650 165926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 171306 592650 171926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 177306 592650 177926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 183306 592650 183926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 189306 592650 189926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 195306 592650 195926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 201306 592650 201926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 207306 592650 207926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 213306 592650 213926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 219306 592650 219926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 225306 592650 225926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 231306 592650 231926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 237306 592650 237926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 243306 592650 243926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 249306 592650 249926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 255306 592650 255926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 261306 592650 261926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 267306 592650 267926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 273306 592650 273926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 279306 592650 279926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 285306 592650 285926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 291306 592650 291926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 297306 592650 297926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 303306 592650 303926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 309306 592650 309926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 315306 592650 315926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 321306 592650 321926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 327306 592650 327926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 333306 592650 333926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 339306 592650 339926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 345306 592650 345926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 351306 592650 351926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 357306 592650 357926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 363306 592650 363926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 369306 592650 369926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 375306 592650 375926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 381306 592650 381926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 387306 592650 387926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 393306 592650 393926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 399306 592650 399926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 405306 592650 405926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 411306 592650 411926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 417306 592650 417926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 423306 592650 423926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 429306 592650 429926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 435306 592650 435926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 441306 592650 441926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 447306 592650 447926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 453306 592650 453926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 459306 592650 459926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 465306 592650 465926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 471306 592650 471926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 477306 592650 477926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 483306 592650 483926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 489306 592650 489926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 495306 592650 495926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 501306 592650 501926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 507306 592650 507926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 513306 592650 513926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 519306 592650 519926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 525306 592650 525926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 531306 592650 531926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 537306 592650 537926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 543306 592650 543926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 549306 592650 549926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 555306 592650 555926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 561306 592650 561926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 567306 592650 567926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 573306 592650 573926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 579306 592650 579926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 585306 592650 585926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 591306 592650 591926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 597306 592650 597926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 603306 592650 603926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 609306 592650 609926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 615306 592650 615926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 621306 592650 621926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 627306 592650 627926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 633306 592650 633926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 639306 592650 639926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 645306 592650 645926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 651306 592650 651926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 657306 592650 657926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 663306 592650 663926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 669306 592650 669926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 675306 592650 675926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 681306 592650 681926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 687306 592650 687926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 693306 592650 693926 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 699306 592650 699926 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 103312 21930 107216 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 33136 93874 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122326 215920 122946 218192 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 67408 157906 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 221502 195248 222122 208400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 131056 287810 147472 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 119088 314858 122992 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 256176 350002 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378270 535792 378890 538064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 318736 414034 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442302 614672 442922 616944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 381296 477882 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 275760 566570 286736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 159344 21930 170320 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 65232 93874 82736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122326 175120 122946 177392 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 33136 157906 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 221502 383472 222122 396624 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 193072 287810 210576 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 215920 314858 223632 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 130512 350002 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378270 614672 378890 616944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 256176 414034 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442302 661456 442922 663728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 318736 477882 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 562086 338864 562706 349296 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 221904 21930 232880 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 130512 93874 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122326 614672 122946 616944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 193072 157906 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 221502 35312 222122 48464 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 67952 287810 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 90800 314858 105040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 318736 350002 336240 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378270 175120 378890 177392 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 381296 414034 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 159344 443106 175120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 256176 477882 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 401424 566570 412400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 285008 21930 295440 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 193072 93874 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 103312 123130 120816 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 130512 157906 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 221502 634800 222122 647952 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 33136 287810 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 153360 314858 161072 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 67408 350002 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378270 215920 378890 218192 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 444400 414034 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437702 175120 438322 177392 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 506960 477882 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 562086 464528 562706 474960 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 347568 21930 358544 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 256176 93874 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 159344 123130 175040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 318736 157906 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 381296 287810 398800 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 238224 314858 248656 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 193072 350002 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378270 661456 378890 663728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 67408 414034 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 285008 443106 302512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 130512 477882 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 87536 566570 105040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 410672 21930 421104 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 318736 93874 336240 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 221904 123130 239952 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 257904 157906 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 444400 287810 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 175120 314858 186096 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 381296 350002 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 103312 379074 120816 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 130512 414034 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 473232 443106 491280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 67408 477882 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 150096 566570 161072 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 473232 21930 484208 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 381296 93874 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 285008 123130 302512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 444400 157906 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 256176 287810 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 341584 314858 349296 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 506960 350002 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 159344 379074 175040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 193072 414034 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 103312 443106 120816 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 568976 477882 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 562086 213200 562706 223632 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 536336 21930 546768 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 444400 93874 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 347568 123130 365616 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 381296 157906 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 319280 287810 335696 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 279024 314858 286736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 33136 350002 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 221904 379074 239952 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 506960 414034 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 410672 443106 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 193072 477882 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 590192 566570 600624 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 598896 21930 609872 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 506960 93874 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 410672 123130 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 570704 157906 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 632624 287810 650128 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 300784 314858 311760 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 444400 350002 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 347568 379074 365616 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 33136 414034 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 221904 443106 239952 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 527088 566570 538064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 21310 662000 21930 672432 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 568976 93874 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 473232 123130 491280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 506960 157906 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 363888 314858 374320 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 632624 350002 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 285008 379074 302512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 536336 443106 553840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 33136 477882 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 105120 567122 109392 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 60318 196336 60938 208400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 93254 632624 93874 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 536336 123130 553840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 507504 287810 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 404688 314858 412400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 349382 568976 350002 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 473232 379074 491280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 598896 443106 614592 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 444400 477882 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 565950 652752 566570 663728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 60318 384560 60938 396624 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 598896 123130 614592 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157286 632624 157906 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 287190 569520 287810 585936 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 426448 314858 437424 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 538144 379074 553840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 663808 443106 679504 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 161152 567122 171952 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 66390 36400 67010 48464 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122510 662000 123130 679504 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 467248 314858 474960 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 598896 379074 614592 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 570704 414034 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442486 347568 443106 365616 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477262 632624 477882 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 567422 222448 568042 235056 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 33136 127914 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 306878 489552 307498 499984 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 663808 379074 679504 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 413414 632624 414034 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 67408 447890 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 286816 567122 297616 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 67408 127914 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 530352 314858 538064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 33136 384042 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 87536 443474 92528 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 567422 347568 568042 360720 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 87536 123498 92528 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 552112 314858 563088 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378454 410672 379074 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 33136 447890 50640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 538144 567122 548944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 130512 127914 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 592912 314858 600624 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 67408 384042 85456 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 150096 443474 155088 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 412480 567122 423280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 150096 123498 155088 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 614672 314858 625648 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 87536 379442 92528 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 130512 447890 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 600704 567122 611504 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 193072 127914 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 652752 314858 663728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 130512 384042 148016 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 213200 443474 217648 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 567422 473776 568042 485840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 213200 123498 215840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314238 677776 314858 688208 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 150096 379442 155088 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 193072 447890 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 566502 663808 567122 674608 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 126926 255632 127546 257904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 105120 315226 119008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 193072 384042 211120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 275760 443474 280752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 257984 127914 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 161152 315226 175040 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 213200 379442 215840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 318736 447890 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 275760 123498 280752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 158758 256176 159378 258992 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 223712 315226 238144 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 318736 384042 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 441382 334512 442002 336784 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 318736 127914 334512 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 286816 315226 300704 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 256176 384042 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 338864 443474 343312 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121406 334512 122026 336784 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 349376 315226 363808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 275760 379442 280752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 256176 447890 273680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 338864 123498 343312 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 158758 333424 159378 336240 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 412480 315226 426368 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 381296 384042 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 401424 443474 406416 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 381296 127914 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 475040 315226 491280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 377350 334512 377970 336784 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 444400 447890 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 401424 123498 406416 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 538144 315226 552032 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 338864 379442 343312 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 414886 333424 415506 336240 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 381296 447890 399344 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 444400 127914 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 600704 315226 614592 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 401424 379442 406416 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 464528 443474 468976 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 478918 333424 479538 336240 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 464528 123498 468976 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314606 663808 315226 677696 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 444400 384042 461904 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 506960 447890 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 506960 127914 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 87536 315410 90720 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 464528 379442 468976 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 527088 443474 532080 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 527088 123498 532080 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 150096 315410 153280 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 506960 384042 525008 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 568976 447890 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 126926 568432 127546 570704 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 213200 315410 215840 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 527088 379442 532080 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 442854 590192 443474 594640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 570784 127914 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 275760 315410 278944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 378822 590192 379442 594640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 447270 632624 447890 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 126926 589648 127546 591920 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 338864 315410 341504 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 382870 568432 383490 570704 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 122878 591280 123498 594640 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 158758 568976 159378 571792 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 401424 315410 404608 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 632624 384042 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127294 632624 127914 650672 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 464528 315410 467168 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 383422 570784 384042 586480 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 527088 315410 530272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 414886 568976 415506 571792 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 314790 590192 315410 592832 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 994 -7654 1614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 -7654 37614 65388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 83364 37614 105988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 117980 37614 128188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 146164 37614 162188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 174180 37614 190988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 208964 37614 224988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 236980 37614 253788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 271764 37614 287788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 299780 37614 316588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 334564 37614 350588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 362580 37614 379388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 397364 37614 413388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 425380 37614 442188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 460164 37614 476188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 488180 37614 504988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 522964 37614 538988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 550980 37614 567788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 585764 37614 601788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 613780 37614 664588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 36994 676580 37614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 -7654 73614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 110593 73614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 173393 73614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 236193 73614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 298993 73614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 361793 73614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 424593 73614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 487393 73614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 550193 73614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 612993 73614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72994 675793 73614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 -7654 109614 35988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 55596 109614 65063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 89348 109614 105988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 117980 109614 127863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 152148 109614 162188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 174180 109614 190663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 214948 109614 224988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 236980 109614 253463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 277748 109614 287788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 299780 109614 316263 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 340548 109614 350588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 362580 109614 379063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 403348 109614 413388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 425380 109614 441863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 466148 109614 476188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 488180 109614 504663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 528948 109614 538988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 550980 109614 567463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 591748 109614 601788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 613780 109614 629175 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 650196 109614 664588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 108994 676580 109614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 -7654 145614 35988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 47980 145614 68567 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 82380 145614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 120332 145614 131367 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 145180 145614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 183132 145614 194167 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 207980 145614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 245932 145614 256967 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 270780 145614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 308732 145614 319767 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 333580 145614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 371532 145614 382567 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 396380 145614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 434332 145614 445367 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 459180 145614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 497132 145614 508167 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 521980 145614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 559932 145614 569767 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 583580 145614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 622732 145614 635588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 144994 647580 145614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 180994 -7654 181614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 -7654 217614 35988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 47980 217614 70388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 82380 217614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 110593 217614 133188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 145180 217614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 173393 217614 195988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 207980 217614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 236193 217614 258788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 270780 217614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 298993 217614 321588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 333580 217614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 361793 217614 384388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 396380 217614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 424593 217614 447188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 459180 217614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 487393 217614 509988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 521980 217614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 550193 217614 571588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 583580 217614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 612993 217614 635588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 647580 217614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 216994 675793 217614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 252994 -7654 253614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 -7654 289614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 110593 289614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 173393 289614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 236193 289614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 298993 289614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 361793 289614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 424593 289614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 487393 289614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 550193 289614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 612993 289614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 288994 675793 289614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 324994 -7654 325614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 -7654 361614 65063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 88313 361614 105988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 117980 361614 127863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 151113 361614 162188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 174180 361614 190663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 213913 361614 224988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 236980 361614 253463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 276713 361614 287788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 299780 361614 316263 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 339513 361614 350588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 362580 361614 379063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 402313 361614 413388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 425380 361614 441863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 465113 361614 476188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 488180 361614 504663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 527913 361614 538988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 550980 361614 567463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 590713 361614 601788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 613780 361614 629175 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 647257 361614 664588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 360994 676580 361614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 -7654 397614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 110593 397614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 173393 397614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 236193 397614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 298993 397614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 361793 397614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 424593 397614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 487393 397614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 550193 397614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 612993 397614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 396994 675793 397614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 -7654 433614 35988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 55596 433614 65063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 89348 433614 105988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 117980 433614 127863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 152148 433614 162188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 174180 433614 190663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 214948 433614 224988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 236980 433614 253463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 277748 433614 287788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 299780 433614 316263 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 340548 433614 350588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 362580 433614 379063 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 403348 433614 413388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 425380 433614 441863 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 466148 433614 476188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 488180 433614 504663 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 528948 433614 538988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 550980 433614 567463 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 591748 433614 601788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 613780 433614 629175 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 650196 433614 664588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 432994 676580 433614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 12780 469614 35988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 47980 469614 70388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 82380 469614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 120332 469614 133188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 145180 469614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 183132 469614 195988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 207980 469614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 245932 469614 258788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 270780 469614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 308732 469614 321588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 333580 469614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 371532 469614 384388 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 396380 469614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 434332 469614 447188 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 459180 469614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 497132 469614 509988 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 521980 469614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 559932 469614 571588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 583580 469614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 622732 469614 635588 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 647580 469614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 468994 685532 469614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 504994 -7654 505614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 -7654 541614 90199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 110593 541614 152999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 173393 541614 215799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 236193 541614 278599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 298993 541614 341399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 361793 541614 404199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 424593 541614 466999 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 487393 541614 529799 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 550193 541614 592599 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 612993 541614 655399 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 540994 675793 541614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 576994 -7654 577614 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 2066 592650 2686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 8066 592650 8686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 14066 592650 14686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 20066 592650 20686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 26066 592650 26686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 32066 592650 32686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 38066 592650 38686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 44066 592650 44686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 50066 592650 50686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 56066 592650 56686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 62066 592650 62686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 68066 592650 68686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 74066 592650 74686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 80066 592650 80686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 86066 592650 86686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 92066 592650 92686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 98066 592650 98686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 104066 592650 104686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 110066 592650 110686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 116066 592650 116686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 122066 592650 122686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 128066 592650 128686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 134066 592650 134686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 140066 592650 140686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 146066 592650 146686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 152066 592650 152686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 158066 592650 158686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 164066 592650 164686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 170066 592650 170686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 176066 592650 176686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 182066 592650 182686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 188066 592650 188686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 194066 592650 194686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 200066 592650 200686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 206066 592650 206686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 212066 592650 212686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 218066 592650 218686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 224066 592650 224686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 230066 592650 230686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 236066 592650 236686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 242066 592650 242686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 248066 592650 248686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 254066 592650 254686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 260066 592650 260686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 266066 592650 266686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 272066 592650 272686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 278066 592650 278686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 284066 592650 284686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 290066 592650 290686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 296066 592650 296686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 302066 592650 302686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 308066 592650 308686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 314066 592650 314686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 320066 592650 320686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 326066 592650 326686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 332066 592650 332686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 338066 592650 338686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 344066 592650 344686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 350066 592650 350686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 356066 592650 356686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 362066 592650 362686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 368066 592650 368686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 374066 592650 374686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 380066 592650 380686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 386066 592650 386686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 392066 592650 392686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 398066 592650 398686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 404066 592650 404686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 410066 592650 410686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 416066 592650 416686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 422066 592650 422686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 428066 592650 428686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 434066 592650 434686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 440066 592650 440686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 446066 592650 446686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 452066 592650 452686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 458066 592650 458686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 464066 592650 464686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 470066 592650 470686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 476066 592650 476686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 482066 592650 482686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 488066 592650 488686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 494066 592650 494686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 500066 592650 500686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 506066 592650 506686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 512066 592650 512686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 518066 592650 518686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 524066 592650 524686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 530066 592650 530686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 536066 592650 536686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 542066 592650 542686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 548066 592650 548686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 554066 592650 554686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 560066 592650 560686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 566066 592650 566686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 572066 592650 572686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 578066 592650 578686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 584066 592650 584686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 590066 592650 590686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 596066 592650 596686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 602066 592650 602686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 608066 592650 608686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 614066 592650 614686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 620066 592650 620686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 626066 592650 626686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 632066 592650 632686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 638066 592650 638686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 644066 592650 644686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 650066 592650 650686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 656066 592650 656686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 662066 592650 662686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 668066 592650 668686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 674066 592650 674686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 680066 592650 680686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 686066 592650 686686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 692066 592650 692686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 698066 592650 698686 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 103312 22666 107216 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 159888 54314 176304 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 33136 97738 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126190 215920 126810 218192 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 67408 161770 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 109840 189002 112112 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 225366 195248 225986 208400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 119088 318722 122992 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 256176 353866 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382134 535792 382754 538064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 318736 417898 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446166 614672 446786 616944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 381296 481746 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 543134 509136 543754 522288 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 275760 567306 286736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 339408 580370 360176 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 159344 22666 170320 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 103312 54314 120816 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 65232 97738 82736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126190 175120 126810 177392 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 33136 161770 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 226256 189002 236144 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 225366 383472 225986 396624 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 215920 318722 223632 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 130512 353866 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382134 614672 382754 616944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 256176 417898 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446166 661456 446786 663728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 318736 481746 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 565950 338864 566570 349296 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 276304 580370 297072 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 221904 22666 232880 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 285008 54314 302512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 130512 97738 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126190 614672 126810 616944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 193072 161770 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 106576 189002 108848 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 225366 35312 225986 48464 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 90800 318722 105040 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 318736 353866 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382134 175120 382754 177392 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 381296 417898 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 159344 446970 175120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 256176 481746 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 401424 567306 412400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 464528 580370 485296 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 285008 22666 295440 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 221904 54314 239408 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 193072 97738 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 103312 126994 120816 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 130512 161770 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 162064 189002 174128 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 225366 634800 225986 647952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 153360 318722 161072 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 67408 353866 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382134 215920 382754 218192 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 444400 417898 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 441566 175120 442186 177392 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 506960 481746 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 543134 320912 543754 334064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 565950 464528 566570 474960 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 401424 580370 423280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 347568 22666 358544 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 411216 54314 427632 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 256176 97738 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 159344 126994 175040 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 318736 161770 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 113104 189002 115376 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 33680 223778 35952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 238224 318722 248656 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 193072 353866 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382134 661456 382754 663728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 67408 417898 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 285008 446970 302512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 130512 481746 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 87536 567306 105040 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 213200 580370 235056 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 410672 22666 421104 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 348112 54314 365616 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 318736 97738 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 221904 126994 239952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 257904 161770 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 288272 189002 290544 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 38032 223778 41392 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 175120 318722 186096 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 381296 353866 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 103312 382938 120816 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 130512 417898 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 473232 446970 491280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 67408 481746 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 150096 567306 161072 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 527632 580370 548400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 473232 22666 484208 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 536336 54314 553840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 381296 97738 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 285008 126994 302512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 444400 161770 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 350288 189002 352560 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 43472 223778 46832 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 341584 318722 349296 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 506960 353866 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 159344 382938 175040 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 193072 417898 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 103312 446970 120816 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 568976 481746 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 543134 69584 543754 82736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 565950 213200 566570 223632 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 590736 580370 611504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 536336 22666 546768 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 473232 54314 490736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 444400 97738 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 347568 126994 365616 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 381296 161770 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 291536 189002 293808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 67408 223778 84912 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 279024 318722 286736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 33136 353866 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 221904 382938 239952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 506960 417898 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 410672 446970 428176 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 193072 481746 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 590192 567306 600624 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 88080 580370 108848 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 598896 22666 609872 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 662544 54314 678960 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 506960 97738 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 410672 126994 428176 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 570704 161770 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 294800 189002 297072 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 130512 223778 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 300784 318722 311760 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 444400 353866 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 347568 382938 365616 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 33136 417898 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 221904 446970 239952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 527088 567306 538064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 150096 580370 171952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22046 662000 22666 672432 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 53694 599440 54314 615856 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 568976 97738 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 473232 126994 491280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 506960 161770 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 353552 189002 355824 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 193616 223778 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 363888 318722 374320 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 632624 353866 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 285008 382938 302512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 536336 446970 553840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 33136 481746 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 105120 567858 109392 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 97118 632624 97738 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 536336 126994 553840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 356816 189002 359088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 257904 223778 273136 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 404688 318722 412400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 353246 568976 353866 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 473232 382938 491280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 598896 446970 614592 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 444400 481746 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 566686 652752 567306 663728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 598896 126994 614592 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 161150 632624 161770 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 360080 189002 362352 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 318736 223778 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 426448 318722 437424 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 538144 382938 553840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 663808 446970 679504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 161152 567858 171952 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126374 662000 126994 679504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 415568 189002 417840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 381840 223778 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 467248 318722 474960 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 598896 382938 614592 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 570704 417898 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446350 347568 446970 365616 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 481126 632624 481746 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 568158 222448 568778 235056 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 33136 131778 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 418832 189002 421104 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 444944 223778 461360 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 310742 489552 311362 499984 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 663808 382938 679504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 417278 632624 417898 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 67408 451754 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 286816 567858 297616 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 67408 131778 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 422096 189002 424368 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 506960 223778 524464 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 530352 318722 538064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 33136 387906 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 87536 447338 92528 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 568158 347568 568778 360720 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 579750 652752 580370 674608 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 87536 127362 92528 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 477584 189002 479856 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 568976 223778 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 552112 318722 563088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382318 410672 382938 428176 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 33136 451754 50640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 538144 567858 548944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 130512 131778 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 480848 189002 483120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 633168 223778 636528 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 592912 318722 600624 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 67408 387906 85456 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 150096 447338 155088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 412480 567858 423280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 150096 127362 155088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 484112 189002 486384 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 637520 223778 639792 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 614672 318722 625648 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 87536 383306 92528 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 130512 451754 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 600704 567858 611504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 193072 131778 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 539600 189002 541872 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 640784 223778 643056 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 652752 318722 663728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 130512 387906 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 213200 447338 217648 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 568158 473776 568778 485840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 213200 127362 215840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 542864 189002 545136 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 644048 223778 646320 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318102 677776 318722 688208 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 150096 383306 155088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 193072 451754 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 567238 663808 567858 674608 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 130790 255632 131410 257904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 546128 189002 548400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 647312 223778 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 105120 319090 119008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 193072 387906 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 275760 447338 280752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 257984 131778 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 601616 189002 603888 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 161152 319090 175040 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 213200 383306 215840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 318736 451754 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 275760 127362 280752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 159494 256176 160114 258992 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 604880 189002 607152 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 223712 319090 238144 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 318736 387906 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 445246 334512 445866 336784 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 318736 131778 334512 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 608144 189002 610416 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 286816 319090 300704 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 256176 387906 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 338864 447338 343312 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 125270 334512 125890 336784 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 611408 189002 613680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 349376 319090 363808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 275760 383306 280752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 256176 451754 273680 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 338864 127362 343312 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 159494 333424 160114 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 666896 189002 669168 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 412480 319090 426368 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 381296 387906 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 401424 447338 406416 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 381296 131778 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 670160 189002 672432 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 475040 319090 491280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 381214 334512 381834 336784 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 444400 451754 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 401424 127362 406416 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188382 673424 189002 675696 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 538144 319090 552032 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 338864 383306 343312 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 415622 333424 416242 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 381296 451754 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 444400 131778 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 33680 193786 48912 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 600704 319090 614592 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 401424 383306 406416 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 464528 447338 468976 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 479654 333424 480274 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 464528 127362 468976 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 203654 48912 204274 51184 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318470 663808 319090 677696 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 444400 387906 461904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 506960 451754 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 506960 131778 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 67408 193786 84912 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 223158 47824 223778 50096 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 87536 319274 90720 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 464528 383306 468976 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 527088 447338 532080 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 527088 127362 532080 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 88080 189370 92528 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 150096 319274 153280 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 506960 387906 525008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 568976 451754 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 130790 568432 131410 570704 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 130512 193786 148016 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 213200 319274 215840 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 527088 383306 532080 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 446718 590192 447338 594640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 570784 131778 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 150096 189370 154544 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 275760 319274 278944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382686 590192 383306 594640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 451134 632624 451754 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 130790 589648 131410 591920 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 193616 193786 211120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 338864 319274 341504 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 386734 568432 387354 570704 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126742 592000 127362 594640 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 159494 568976 160114 571792 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 213200 189370 217648 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 401424 319274 404608 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 632624 387906 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 131158 632624 131778 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 203654 255632 204274 257904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 464528 319274 467168 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 387286 570784 387906 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 257808 193786 273136 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 527088 319274 530272 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 415622 568976 416242 571792 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 276304 189370 280752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 222054 256720 222674 258992 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 318654 590192 319274 592832 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 318736 193786 336240 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 339408 189370 342768 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 381840 193786 399344 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 401424 189370 405872 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 444944 193786 461360 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 464528 189370 468976 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 506960 193786 524464 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 527632 189370 532080 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 568976 193786 586480 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188750 590736 189370 594096 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 193166 633168 193786 650672 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 118690694
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/user_project_wrapper/runs/24_04_02_10_01/results/signoff/user_project_wrapper.magic.gds
string GDS_START 12030138
<< end >>

