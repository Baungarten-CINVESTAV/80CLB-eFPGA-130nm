magic
tech sky130A
magscale 1 2
timestamp 1708041631
<< obsli1 >>
rect 1104 2159 14812 17425
<< obsm1 >>
rect 934 2128 15074 17456
<< metal2 >>
rect 2134 0 2190 800
rect 3422 0 3478 800
rect 4710 0 4766 800
rect 5998 0 6054 800
rect 7286 0 7342 800
rect 8574 0 8630 800
rect 9862 0 9918 800
rect 11150 0 11206 800
rect 12438 0 12494 800
rect 13726 0 13782 800
rect 15014 0 15070 800
<< obsm2 >>
rect 938 856 15068 18601
rect 938 734 2078 856
rect 2246 734 3366 856
rect 3534 734 4654 856
rect 4822 734 5942 856
rect 6110 734 7230 856
rect 7398 734 8518 856
rect 8686 734 9806 856
rect 9974 734 11094 856
rect 11262 734 12382 856
rect 12550 734 13670 856
rect 13838 734 14958 856
<< metal3 >>
rect 0 18504 800 18624
rect 15200 17960 16000 18080
rect 0 17688 800 17808
rect 0 16872 800 16992
rect 15200 16328 16000 16448
rect 0 16056 800 16176
rect 0 15240 800 15360
rect 15200 14696 16000 14816
rect 0 14424 800 14544
rect 0 13608 800 13728
rect 15200 13064 16000 13184
rect 0 12792 800 12912
rect 0 11976 800 12096
rect 15200 11432 16000 11552
rect 0 11160 800 11280
rect 0 10344 800 10464
rect 15200 9800 16000 9920
rect 0 9528 800 9648
rect 0 8712 800 8832
rect 15200 8168 16000 8288
rect 0 7896 800 8016
rect 0 7080 800 7200
rect 15200 6536 16000 6656
rect 0 6264 800 6384
rect 0 5448 800 5568
rect 15200 4904 16000 5024
rect 0 4632 800 4752
rect 0 3816 800 3936
rect 15200 3272 16000 3392
rect 0 3000 800 3120
rect 0 2184 800 2304
rect 15200 1640 16000 1760
<< obsm3 >>
rect 880 18424 15210 18597
rect 798 18160 15210 18424
rect 798 17888 15120 18160
rect 880 17880 15120 17888
rect 880 17608 15210 17880
rect 798 17072 15210 17608
rect 880 16792 15210 17072
rect 798 16528 15210 16792
rect 798 16256 15120 16528
rect 880 16248 15120 16256
rect 880 15976 15210 16248
rect 798 15440 15210 15976
rect 880 15160 15210 15440
rect 798 14896 15210 15160
rect 798 14624 15120 14896
rect 880 14616 15120 14624
rect 880 14344 15210 14616
rect 798 13808 15210 14344
rect 880 13528 15210 13808
rect 798 13264 15210 13528
rect 798 12992 15120 13264
rect 880 12984 15120 12992
rect 880 12712 15210 12984
rect 798 12176 15210 12712
rect 880 11896 15210 12176
rect 798 11632 15210 11896
rect 798 11360 15120 11632
rect 880 11352 15120 11360
rect 880 11080 15210 11352
rect 798 10544 15210 11080
rect 880 10264 15210 10544
rect 798 10000 15210 10264
rect 798 9728 15120 10000
rect 880 9720 15120 9728
rect 880 9448 15210 9720
rect 798 8912 15210 9448
rect 880 8632 15210 8912
rect 798 8368 15210 8632
rect 798 8096 15120 8368
rect 880 8088 15120 8096
rect 880 7816 15210 8088
rect 798 7280 15210 7816
rect 880 7000 15210 7280
rect 798 6736 15210 7000
rect 798 6464 15120 6736
rect 880 6456 15120 6464
rect 880 6184 15210 6456
rect 798 5648 15210 6184
rect 880 5368 15210 5648
rect 798 5104 15210 5368
rect 798 4832 15120 5104
rect 880 4824 15120 4832
rect 880 4552 15210 4824
rect 798 4016 15210 4552
rect 880 3736 15210 4016
rect 798 3472 15210 3736
rect 798 3200 15120 3472
rect 880 3192 15120 3200
rect 880 2920 15210 3192
rect 798 2384 15210 2920
rect 880 2104 15210 2384
rect 798 1840 15210 2104
rect 798 1667 15120 1840
<< metal4 >>
rect 2657 2128 2977 17456
rect 4370 2128 4690 17456
rect 6084 2128 6404 17456
rect 7797 2128 8117 17456
rect 9511 2128 9831 17456
rect 11224 2128 11544 17456
rect 12938 2128 13258 17456
rect 14651 2128 14971 17456
<< labels >>
rlabel metal2 s 13726 0 13782 800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 1 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
rlabel metal3 s 15200 1640 16000 1760 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 15200 3272 16000 3392 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[0]
port 5 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[1]
port 6 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[2]
port 7 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[3]
port 8 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 chanx_left_in[4]
port 9 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 chanx_left_in[5]
port 10 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 chanx_left_in[6]
port 11 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 chanx_left_in[7]
port 12 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 chanx_left_in[8]
port 13 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[0]
port 14 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[1]
port 15 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[2]
port 16 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[3]
port 17 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 chanx_left_out[4]
port 18 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 chanx_left_out[5]
port 19 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 chanx_left_out[6]
port 20 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 chanx_left_out[7]
port 21 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 chanx_left_out[8]
port 22 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_in[0]
port 23 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[1]
port 24 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[2]
port 25 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[3]
port 26 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[4]
port 27 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[5]
port 28 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[6]
port 29 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[7]
port 30 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_in[8]
port 31 nsew signal input
rlabel metal3 s 15200 4904 16000 5024 6 chany_bottom_out[0]
port 32 nsew signal output
rlabel metal3 s 15200 6536 16000 6656 6 chany_bottom_out[1]
port 33 nsew signal output
rlabel metal3 s 15200 8168 16000 8288 6 chany_bottom_out[2]
port 34 nsew signal output
rlabel metal3 s 15200 9800 16000 9920 6 chany_bottom_out[3]
port 35 nsew signal output
rlabel metal3 s 15200 11432 16000 11552 6 chany_bottom_out[4]
port 36 nsew signal output
rlabel metal3 s 15200 13064 16000 13184 6 chany_bottom_out[5]
port 37 nsew signal output
rlabel metal3 s 15200 14696 16000 14816 6 chany_bottom_out[6]
port 38 nsew signal output
rlabel metal3 s 15200 16328 16000 16448 6 chany_bottom_out[7]
port 39 nsew signal output
rlabel metal3 s 15200 17960 16000 18080 6 chany_bottom_out[8]
port 40 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 41 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 42 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 prog_clk
port 43 nsew signal input
rlabel metal4 s 2657 2128 2977 17456 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 17456 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 17456 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 17456 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 17456 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 17456 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 17456 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 17456 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 429044
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_8__10_/runs/24_02_15_17_59/results/signoff/sb_8__10_.magic.gds
string GDS_START 89996
<< end >>

