* NGSPICE file created from sb_8__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

.subckt sb_8__1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
+ prog_clk top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ vdd vss
XFILLER_0_27_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_294_ mem_bottom_track_1.DFF_2_.Q vss vss vdd vdd _039_ sky130_fd_sc_hd__clkbuf_1
X_363_ mux_left_track_1.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net36 sky130_fd_sc_hd__inv_2
X_501_ mux_bottom_track_1.INVTX1_4_.out _105_ vss vss vdd vdd mux_top_track_16.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_108 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_3_28 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_1_130 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_346_ net26 vss vss vdd vdd mux_bottom_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_415_ clknet_2_0__leaf_prog_clk net98 vss vss vdd vdd mem_left_track_11.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_277_ _033_ vss vss vdd vdd _090_ sky130_fd_sc_hd__clkbuf_1
X_200_ mem_left_track_11.DFF_0_.D vss vss vdd vdd _144_ sky130_fd_sc_hd__inv_2
X_329_ _050_ vss vss vdd vdd _056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_136 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_21_95 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold30 mem_top_track_8.DFF_1_.Q vss vss vdd vdd net107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_8 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_6_39 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput53 net53 vss vss vdd vdd chany_bottom_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 vss vss vdd vdd chanx_left_out[6] sky130_fd_sc_hd__clkbuf_4
XTAP_123 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ net10 vss vss vdd vdd mux_bottom_track_17.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_293_ _038_ vss vss vdd vdd _082_ sky130_fd_sc_hd__clkbuf_1
X_500_ mux_top_track_16.mux_l1_in_1_.TGATE_0_.out _104_ vss vss vdd vdd mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_142 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_276_ mem_bottom_track_17.DFF_0_.D vss vss vdd vdd _033_ sky130_fd_sc_hd__clkbuf_1
X_345_ net2 vss vss vdd vdd mux_bottom_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_414_ clknet_2_0__leaf_prog_clk net78 vss vss vdd vdd mem_left_track_9.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_259_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _027_ sky130_fd_sc_hd__clkbuf_1
X_328_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _050_ sky130_fd_sc_hd__clkbuf_1
Xhold31 mem_bottom_track_9.DFF_1_.Q vss vss vdd vdd net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 mem_left_track_13.DFF_1_.Q vss vss vdd vdd net97 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_62 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_21_132 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput43 net43 vss vss vdd vdd chanx_left_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 vss vss vdd vdd chany_top_out[0] sky130_fd_sc_hd__buf_2
XTAP_124 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ net24 vss vss vdd vdd mux_bottom_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_292_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_20 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_275_ _032_ vss vss vdd vdd _094_ sky130_fd_sc_hd__clkbuf_1
X_344_ net5 vss vss vdd vdd mux_bottom_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_413_ clknet_2_0__leaf_prog_clk net92 vss vss vdd vdd mem_left_track_11.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
X_258_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _110_ sky130_fd_sc_hd__inv_2
X_189_ mem_left_track_13.DFF_0_.Q vss vss vdd vdd _153_ sky130_fd_sc_hd__inv_2
X_327_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _064_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_74 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xhold32 mem_top_track_0.DFF_1_.Q vss vss vdd vdd net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 mem_top_track_16.DFF_0_.D vss vss vdd vdd net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 mem_left_track_11.DFF_0_.Q vss vss vdd vdd net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_111 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput44 net44 vss vss vdd vdd chanx_left_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 vss vss vdd vdd chany_top_out[1] sky130_fd_sc_hd__buf_2
XTAP_125 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_27_63 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_27_52 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XTAP_114 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_7 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_360_ net28 vss vss vdd vdd mux_bottom_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_291_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _088_ sky130_fd_sc_hd__inv_2
X_489_ mux_bottom_track_9.INVTX1_5_.out _093_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_13_98 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_65 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_343_ net8 vss vss vdd vdd mux_bottom_track_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_274_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _032_ sky130_fd_sc_hd__clkbuf_1
X_412_ clknet_2_0__leaf_prog_clk net93 vss vss vdd vdd mem_left_track_7.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_519__69 vss vss vdd vdd net69 _519__69/LO sky130_fd_sc_hd__conb_1
XFILLER_0_19_97 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_188_ mem_left_track_13.DFF_1_.Q vss vss vdd vdd _152_ sky130_fd_sc_hd__inv_2
X_326_ _049_ vss vss vdd vdd _058_ sky130_fd_sc_hd__clkbuf_1
X_257_ _026_ vss vss vdd vdd _104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_88 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_309_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _076_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_97 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xhold11 mem_bottom_track_17.DFF_0_.D vss vss vdd vdd net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 mem_left_track_1.DFF_0_.Q vss vss vdd vdd net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 mem_bottom_track_1.DFF_1_.Q vss vss vdd vdd net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput45 net45 vss vss vdd vdd chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vss vss vdd vdd chany_top_out[2] sky130_fd_sc_hd__clkbuf_4
XTAP_126 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_557_ mux_bottom_track_9.INVTX1_0_.out _161_ vss vss vdd vdd mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_488_ mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out _092_ vss vss vdd vdd mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_290_ _037_ vss vss vdd vdd _080_ sky130_fd_sc_hd__clkbuf_1
X_273_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _100_ sky130_fd_sc_hd__inv_2
X_342_ mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net45 sky130_fd_sc_hd__inv_2
X_411_ clknet_2_1__leaf_prog_clk net82 vss vss vdd vdd mem_left_track_7.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_187_ _003_ vss vss vdd vdd _154_ sky130_fd_sc_hd__clkbuf_1
X_325_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_12 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_256_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _026_ sky130_fd_sc_hd__clkbuf_1
X_239_ mem_bottom_track_17.DFF_0_.Q vss vss vdd vdd _020_ sky130_fd_sc_hd__clkbuf_1
X_308_ _043_ vss vss vdd vdd _068_ sky130_fd_sc_hd__clkbuf_1
Xhold34 mem_bottom_track_17.DFF_0_.Q vss vss vdd vdd net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 mem_left_track_11.DFF_1_.Q vss vss vdd vdd net89 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_3__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_135 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput46 net46 vss vss vdd vdd chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__buf_2
Xoutput57 net57 vss vss vdd vdd chany_top_out[3] sky130_fd_sc_hd__buf_2
XTAP_127 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_487_ net66 _091_ vss vss vdd vdd mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_556_ mux_left_track_17.mux_l1_in_0_.TGATE_0_.out _160_ vss vss vdd vdd mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_341_ net34 vss vss vdd vdd mux_top_track_8.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_272_ _031_ vss vss vdd vdd _092_ sky130_fd_sc_hd__clkbuf_1
X_410_ clknet_2_0__leaf_prog_clk net86 vss vss vdd vdd mem_left_track_5.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_99 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_44 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_539_ mux_left_track_9.INVTX1_1_.out _143_ vss vss vdd vdd mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_4_65 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_186_ mem_left_track_15.DFF_1_.Q vss vss vdd vdd _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_22 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_11 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_324_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _065_ sky130_fd_sc_hd__inv_2
X_542__74 vss vss vdd vdd net74 _542__74/LO sky130_fd_sc_hd__conb_1
XFILLER_0_10_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_255_ _025_ vss vss vdd vdd _106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_238_ mem_bottom_track_17.DFF_0_.Q vss vss vdd vdd _121_ sky130_fd_sc_hd__inv_2
X_307_ mem_top_track_8.DFF_1_.Q vss vss vdd vdd _043_ sky130_fd_sc_hd__clkbuf_1
Xhold13 mem_bottom_track_1.DFF_0_.D vss vss vdd vdd net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 mem_top_track_16.DFF_0_.Q vss vss vdd vdd net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 mem_top_track_0.DFF_0_.Q vss vss vdd vdd net112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_136 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_23 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_119 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput47 net47 vss vss vdd vdd chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vss vss vdd vdd chanx_left_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 vss vss vdd vdd chany_top_out[4] sky130_fd_sc_hd__buf_2
XTAP_128 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_117 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_4_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_555_ mux_left_track_17.INVTX1_1_.out _159_ vss vss vdd vdd mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_486_ mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out _090_ vss vss vdd vdd mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_13_46 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_103 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_271_ mem_bottom_track_9.DFF_1_.Q vss vss vdd vdd _031_ sky130_fd_sc_hd__clkbuf_1
X_538_ net73 _142_ vss vss vdd vdd mux_left_track_9.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_340_ mux_top_track_8.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net58 sky130_fd_sc_hd__inv_2
X_469_ mux_top_track_8.mux_l1_in_2_.TGATE_0_.out _073_ vss vss vdd vdd mux_top_track_8.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_185_ _002_ vss vss vdd vdd _155_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_323_ _048_ vss vss vdd vdd _054_ sky130_fd_sc_hd__clkbuf_1
X_254_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_69 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_237_ mem_bottom_track_17.DFF_1_.Q vss vss vdd vdd _119_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_112 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_21_24 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_306_ _042_ vss vss vdd vdd _071_ sky130_fd_sc_hd__clkbuf_1
Xhold14 mem_bottom_track_17.DFF_2_.Q vss vss vdd vdd net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 mem_top_track_16.DFF_1_.Q vss vss vdd vdd net102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_78 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_57 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput48 net48 vss vss vdd vdd chany_bottom_out[3] sky130_fd_sc_hd__clkbuf_4
Xoutput37 net37 vss vss vdd vdd chanx_left_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput59 net59 vss vss vdd vdd chany_top_out[5] sky130_fd_sc_hd__clkbuf_4
XTAP_129 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_89 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_78 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XTAP_118 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_88 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_485_ mux_bottom_track_1.INVTX1_0_.out _089_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_554_ net77 _158_ vss vss vdd vdd mux_left_track_17.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
Xclkbuf_2_0__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_270_ _030_ vss vss vdd vdd _095_ sky130_fd_sc_hd__clkbuf_1
X_399_ clknet_2_3__leaf_prog_clk net102 vss vss vdd vdd mem_bottom_track_1.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
X_537_ mux_left_track_7.INVTX1_0_.out _141_ vss vss vdd vdd mux_left_track_7.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_4_23 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_468_ mux_top_track_8.mux_l2_in_0_.TGATE_0_.out _072_ vss vss vdd vdd mux_top_track_8.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_322_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _048_ sky130_fd_sc_hd__clkbuf_1
X_184_ mem_left_track_15.DFF_0_.Q vss vss vdd vdd _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_46 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_253_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _111_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_24_124 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_236_ mem_bottom_track_17.DFF_2_.Q vss vss vdd vdd _117_ sky130_fd_sc_hd__inv_2
X_305_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_124 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_102 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold26 mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 mem_left_track_9.DFF_0_.Q vss vss vdd vdd net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_69 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_127 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_219_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _133_ sky130_fd_sc_hd__inv_2
Xoutput49 net49 vss vss vdd vdd chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xoutput38 net38 vss vss vdd vdd chanx_left_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_57 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_119 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_553_ mux_bottom_track_17.INVTX1_0_.out _157_ vss vss vdd vdd mux_left_track_15.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_484_ mux_bottom_track_1.INVTX1_2_.out _088_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_398_ clknet_2_3__leaf_prog_clk net83 vss vss vdd vdd mem_bottom_track_9.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_536_ mux_left_track_7.mux_l1_in_0_.TGATE_0_.out _140_ vss vss vdd vdd mux_left_track_7.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_467_ mux_left_track_5.INVTX1_0_.out _071_ vss vss vdd vdd mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_183_ mem_left_track_15.DFF_0_.Q vss vss vdd vdd _157_ sky130_fd_sc_hd__inv_2
X_252_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _109_ sky130_fd_sc_hd__inv_2
X_321_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _061_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_133 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_90 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_519_ net69 _123_ vss vss vdd vdd mux_left_track_1.mux_l1_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_18_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_24_136 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_235_ _019_ vss vss vdd vdd _123_ sky130_fd_sc_hd__clkbuf_1
X_304_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _077_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_136 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_1_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold16 mem_left_track_5.DFF_1_.Q vss vss vdd vdd net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 mem_left_track_3.DFF_0_.Q vss vss vdd vdd net104 sky130_fd_sc_hd__dlygate4sd3_1
X_218_ mem_left_track_3.DFF_1_.Q vss vss vdd vdd _131_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_6 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xoutput39 net39 vss vss vdd vdd chanx_left_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_109 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_80 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_552_ mux_left_track_15.mux_l1_in_0_.TGATE_0_.out _156_ vss vss vdd vdd mux_left_track_15.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_483_ mux_bottom_track_1.INVTX1_4_.out _087_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_397_ clknet_2_3__leaf_prog_clk net103 vss vss vdd vdd mem_bottom_track_9.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_535_ mux_left_track_7.INVTX1_1_.out _139_ vss vss vdd vdd mux_left_track_7.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_466_ mux_bottom_track_9.INVTX1_3_.out _070_ vss vss vdd vdd mux_top_track_8.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_182_ mem_left_track_15.DFF_1_.Q vss vss vdd vdd _156_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_26 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_251_ mem_bottom_track_1.DFF_0_.D vss vss vdd vdd _107_ sky130_fd_sc_hd__inv_2
X_320_ mem_top_track_0.DFF_2_.Q vss vss vdd vdd _063_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_123 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_518_ mux_left_track_1.mux_l1_in_1_.TGATE_0_.out _122_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_449_ net13 vss vss vdd vdd net55 sky130_fd_sc_hd__buf_1
X_234_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _019_ sky130_fd_sc_hd__clkbuf_1
X_303_ mem_top_track_8.DFF_1_.Q vss vss vdd vdd _074_ sky130_fd_sc_hd__inv_2
Xhold28 mem_bottom_track_17.DFF_1_.Q vss vss vdd vdd net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 mem_left_track_1.DFF_1_.Q vss vss vdd vdd net94 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_217_ _013_ vss vss vdd vdd _134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_48 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_37 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_551_ mux_left_track_15.INVTX1_1_.out _155_ vss vss vdd vdd mux_left_track_15.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_92 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_482_ mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out _086_ vss vss vdd vdd mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_107 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_396_ clknet_2_3__leaf_prog_clk net108 vss vss vdd vdd mem_bottom_track_17.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
X_465_ mux_bottom_track_9.INVTX1_5_.out _069_ vss vss vdd vdd mux_top_track_8.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_534_ net72 _138_ vss vss vdd vdd mux_left_track_7.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
XFILLER_0_4_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_250_ _024_ vss vss vdd vdd _113_ sky130_fd_sc_hd__clkbuf_1
X_181_ _001_ vss vss vdd vdd _158_ sky130_fd_sc_hd__clkbuf_1
X_463__64 vss vss vdd vdd net64 _463__64/LO sky130_fd_sc_hd__conb_1
XFILLER_0_27_113 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_517_ mux_bottom_track_17.INVTX1_0_.out _121_ vss vss vdd vdd mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_448_ net14 vss vss vdd vdd net56 sky130_fd_sc_hd__clkbuf_1
X_379_ net18 vss vss vdd vdd mux_left_track_11.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_233_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _126_ sky130_fd_sc_hd__inv_2
X_302_ mem_top_track_16.DFF_0_.D vss vss vdd vdd _072_ sky130_fd_sc_hd__inv_2
Xhold18 mem_left_track_5.DFF_0_.Q vss vss vdd vdd net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 mem_top_track_8.DFF_0_.Q vss vss vdd vdd net106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_216_ mem_left_track_5.DFF_1_.Q vss vss vdd vdd _013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_550_ net76 _154_ vss vss vdd vdd mux_left_track_15.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_481_ mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.out _085_ vss vss vdd vdd mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_21_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_554__77 vss vss vdd vdd net77 _554__77/LO sky130_fd_sc_hd__conb_1
X_533_ mux_left_track_5.INVTX1_0_.out _137_ vss vss vdd vdd mux_left_track_5.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_464_ mux_top_track_8.mux_l1_in_1_.TGATE_0_.out _068_ vss vss vdd vdd mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_395_ clknet_2_3__leaf_prog_clk net90 vss vss vdd vdd mem_bottom_track_1.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_180_ net35 vss vss vdd vdd _001_ sky130_fd_sc_hd__clkbuf_1
X_516_ mux_bottom_track_17.INVTX1_2_.out _120_ vss vss vdd vdd mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_447_ net15 vss vss vdd vdd net57 sky130_fd_sc_hd__clkbuf_1
X_378_ mux_left_track_11.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net41 sky130_fd_sc_hd__inv_2
X_301_ _041_ vss vss vdd vdd _079_ sky130_fd_sc_hd__clkbuf_1
X_232_ _018_ vss vss vdd vdd _122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_70 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold19 mem_left_track_17.DFF_0_.Q vss vss vdd vdd net96 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_17 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_215_ _012_ vss vss vdd vdd _135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_480_ mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out _084_ vss vss vdd vdd mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_24_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_394_ clknet_2_2__leaf_prog_clk net100 vss vss vdd vdd mem_bottom_track_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_463_ net64 _067_ vss vss vdd vdd mux_top_track_8.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_532_ mux_left_track_5.mux_l1_in_0_.TGATE_0_.out _136_ vss vss vdd vdd mux_left_track_5.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_515_ mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out _119_ vss vss vdd vdd mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_377_ net17 vss vss vdd vdd mux_left_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_446_ net17 vss vss vdd vdd net59 sky130_fd_sc_hd__clkbuf_1
X_300_ mem_bottom_track_1.DFF_1_.Q vss vss vdd vdd _041_ sky130_fd_sc_hd__clkbuf_1
X_231_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _018_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XTAP_90 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ vss vss vdd vdd
+ net1 sky130_fd_sc_hd__buf_1
X_214_ mem_left_track_5.DFF_0_.Q vss vss vdd vdd _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_137 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_27_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_18 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_71 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_393_ clknet_2_3__leaf_prog_clk net99 vss vss vdd vdd mem_bottom_track_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_531_ mux_left_track_5.INVTX1_1_.out _135_ vss vss vdd vdd mux_left_track_5.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_462_ mux_top_track_8.mux_l2_in_1_.TGATE_0_.out _066_ vss vss vdd vdd mux_top_track_8.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_514_ mux_bottom_track_17.INVTX1_4_.out _118_ vss vss vdd vdd mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_509__68 vss vss vdd vdd net68 _509__68/LO sky130_fd_sc_hd__conb_1
X_376_ mux_left_track_9.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net40 sky130_fd_sc_hd__inv_2
X_445_ net18 vss vss vdd vdd net60 sky130_fd_sc_hd__clkbuf_1
X_230_ _017_ vss vss vdd vdd _124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_108 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_359_ net4 vss vss vdd vdd mux_bottom_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_0_11_75 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XTAP_91 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net2 sky130_fd_sc_hd__buf_1
XTAP_80 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ mem_left_track_5.DFF_0_.Q vss vss vdd vdd _137_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_7_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_11_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_2_73 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_16_8 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_18 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_3_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_475__65 vss vss vdd vdd net65 _475__65/LO sky130_fd_sc_hd__conb_1
XFILLER_0_0_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_530_ net71 _134_ vss vss vdd vdd mux_left_track_5.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_392_ clknet_2_1__leaf_prog_clk net84 vss vss vdd vdd mem_top_track_8.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
X_461_ mux_top_track_0.INVTX1_0_.out _065_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_513_ mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out _117_ vss vss vdd vdd mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_444_ net19 vss vss vdd vdd net61 sky130_fd_sc_hd__clkbuf_1
X_375_ net21 vss vss vdd vdd mux_left_track_7.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_18_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_358_ net7 vss vss vdd vdd mux_bottom_track_17.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_289_ mem_bottom_track_1.DFF_1_.Q vss vss vdd vdd _037_ sky130_fd_sc_hd__clkbuf_1
XTAP_92 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 ccff_head vss vss vdd vdd net3 sky130_fd_sc_hd__clkbuf_1
XTAP_70 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ mem_left_track_5.DFF_1_.Q vss vss vdd vdd _136_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_96 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_17_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_5_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_460_ mux_left_track_9.INVTX1_1_.out _064_ vss vss vdd vdd mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_391_ clknet_2_1__leaf_prog_clk net106 vss vss vdd vdd mem_top_track_8.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_129 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_512_ mux_bottom_track_17.INVTX1_1_.out _116_ vss vss vdd vdd mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_443_ net22 vss vss vdd vdd net46 sky130_fd_sc_hd__buf_1
X_374_ net15 vss vss vdd vdd mux_left_track_7.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_25_20 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_357_ mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net53 sky130_fd_sc_hd__inv_2
X_288_ _036_ vss vss vdd vdd _083_ sky130_fd_sc_hd__clkbuf_1
Xinput4 chanx_left_in[0] vss vss vdd vdd net4 sky130_fd_sc_hd__clkbuf_1
XTAP_93 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_211_ _011_ vss vss vdd vdd _138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_21 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_409_ clknet_2_0__leaf_prog_clk net95 vss vss vdd vdd mem_left_track_5.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_135 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_390_ clknet_2_1__leaf_prog_clk net107 vss vss vdd vdd mem_top_track_16.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_119 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_108 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_442_ net23 vss vss vdd vdd net47 sky130_fd_sc_hd__clkbuf_1
X_511_ mux_bottom_track_17.INVTX1_3_.out _115_ vss vss vdd vdd mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_373_ mux_left_track_7.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net39 sky130_fd_sc_hd__inv_2
XFILLER_0_26_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_133 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_23_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_287_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _036_ sky130_fd_sc_hd__clkbuf_1
Xinput5 chanx_left_in[1] vss vss vdd vdd net5 sky130_fd_sc_hd__clkbuf_1
X_356_ mux_top_track_16.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net62 sky130_fd_sc_hd__inv_2
XFILLER_0_14_133 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_94 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ clknet_2_2__leaf_prog_clk net94 vss vss vdd vdd mem_left_track_3.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_210_ mem_left_track_7.DFF_1_.Q vss vss vdd vdd _011_ sky130_fd_sc_hd__clkbuf_1
X_339_ net33 vss vss vdd vdd mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
Xinput30 chany_top_in[8] vss vss vdd vdd net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_99 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_510_ mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.out _114_ vss vss vdd vdd mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_441_ net24 vss vss vdd vdd net48 sky130_fd_sc_hd__clkbuf_1
X_372_ net20 vss vss vdd vdd mux_left_track_5.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_26_131 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_44 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_355_ net12 vss vss vdd vdd mux_bottom_track_9.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_286_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _089_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_24 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput6 chanx_left_in[2] vss vss vdd vdd net6 sky130_fd_sc_hd__clkbuf_1
XTAP_95 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_62 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_89 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_407_ clknet_2_0__leaf_prog_clk net104 vss vss vdd vdd mem_left_track_3.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_338_ mux_top_track_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net54 sky130_fd_sc_hd__inv_2
Xinput31 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ vss vss vdd vdd
+ net31 sky130_fd_sc_hd__clkbuf_1
X_487__66 vss vss vdd vdd net66 _487__66/LO sky130_fd_sc_hd__conb_1
XFILLER_0_17_67 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xinput20 chany_bottom_in[7] vss vss vdd vdd net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_550__76 vss vss vdd vdd net76 _550__76/LO sky130_fd_sc_hd__conb_1
X_440_ net26 vss vss vdd vdd net50 sky130_fd_sc_hd__clkbuf_1
X_371_ net14 vss vss vdd vdd mux_left_track_5.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_3_9 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_66 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_354_ net23 vss vss vdd vdd mux_bottom_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_285_ mem_bottom_track_1.DFF_1_.Q vss vss vdd vdd _086_ sky130_fd_sc_hd__inv_2
Xinput7 chanx_left_in[3] vss vss vdd vdd net7 sky130_fd_sc_hd__clkbuf_1
XTAP_96 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_268_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _101_ sky130_fd_sc_hd__inv_2
X_406_ clknet_2_2__leaf_prog_clk net91 vss vss vdd vdd mem_left_track_1.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_337_ _053_ vss vss vdd vdd _059_ sky130_fd_sc_hd__clkbuf_1
X_199_ _007_ vss vss vdd vdd _146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput32 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_ vss vss vdd vdd
+ net32 sky130_fd_sc_hd__clkbuf_1
Xinput10 chanx_left_in[6] vss vss vdd vdd net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 chany_bottom_in[8] vss vss vdd vdd net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_0_127 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_0_116 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_25_79 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_370_ mux_left_track_5.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net38 sky130_fd_sc_hd__inv_2
X_499_ net67 _103_ vss vss vdd vdd mux_top_track_16.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_353_ net27 vss vss vdd vdd mux_bottom_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_422_ clknet_2_3__leaf_prog_clk net80 vss vss vdd vdd mem_left_track_17.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_284_ mem_bottom_track_1.DFF_2_.Q vss vss vdd vdd _084_ sky130_fd_sc_hd__inv_2
Xinput8 chanx_left_in[4] vss vss vdd vdd net8 sky130_fd_sc_hd__clkbuf_1
XTAP_97 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ mem_bottom_track_9.DFF_1_.Q vss vss vdd vdd _098_ sky130_fd_sc_hd__inv_2
X_405_ clknet_2_2__leaf_prog_clk net110 vss vss vdd vdd mem_left_track_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_336_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _053_ sky130_fd_sc_hd__clkbuf_1
X_198_ mem_left_track_11.DFF_1_.Q vss vss vdd vdd _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput33 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ vss vss vdd vdd
+ net33 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[7] vss vss vdd vdd net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 chany_top_in[0] vss vss vdd vdd net22 sky130_fd_sc_hd__buf_1
X_319_ _047_ vss vss vdd vdd _067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_56 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_498_ mux_top_track_16.mux_l2_in_1_.TGATE_0_.out _102_ vss vss vdd vdd mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_421_ clknet_2_3__leaf_prog_clk net96 vss vss vdd vdd net35 sky130_fd_sc_hd__dfxtp_1
Xinput9 chanx_left_in[5] vss vss vdd vdd net9 sky130_fd_sc_hd__clkbuf_1
X_283_ _035_ vss vss vdd vdd _091_ sky130_fd_sc_hd__clkbuf_1
XTAP_98 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ net1 vss vss vdd vdd mux_bottom_track_9.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XTAP_65 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ mem_bottom_track_17.DFF_0_.D vss vss vdd vdd _096_ sky130_fd_sc_hd__inv_2
X_404_ clknet_2_2__leaf_prog_clk net88 vss vss vdd vdd mem_bottom_track_17.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_129 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_20_107 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_335_ _052_ vss vss vdd vdd _057_ sky130_fd_sc_hd__clkbuf_1
X_197_ _006_ vss vss vdd vdd _147_ sky130_fd_sc_hd__clkbuf_1
Xinput34 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 chany_top_in[1] vss vss vdd vdd net23 sky130_fd_sc_hd__buf_1
Xinput12 chanx_left_in[8] vss vss vdd vdd net12 sky130_fd_sc_hd__buf_1
X_249_ mem_bottom_track_17.DFF_1_.Q vss vss vdd vdd _024_ sky130_fd_sc_hd__clkbuf_1
X_318_ mem_top_track_8.DFF_1_.Q vss vss vdd vdd _047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_104 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_3_137 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_538__73 vss vss vdd vdd net73 _538__73/LO sky130_fd_sc_hd__conb_1
XFILLER_0_12_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold1 mem_left_track_7.DFF_1_.Q vss vss vdd vdd net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_497_ mux_bottom_track_9.INVTX1_0_.out _101_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_420_ clknet_2_3__leaf_prog_clk net97 vss vss vdd vdd mem_left_track_15.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_282_ mem_bottom_track_9.DFF_1_.Q vss vss vdd vdd _035_ sky130_fd_sc_hd__clkbuf_1
X_351_ net6 vss vss vdd vdd mux_bottom_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XTAP_99 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ mux_bottom_track_1.INVTX1_1_.out _153_ vss vss vdd vdd mux_left_track_13.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_88 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_403_ clknet_2_2__leaf_prog_clk net111 vss vss vdd vdd mem_bottom_track_17.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_334_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _052_ sky130_fd_sc_hd__clkbuf_1
X_499__67 vss vss vdd vdd net67 _499__67/LO sky130_fd_sc_hd__conb_1
X_265_ _029_ vss vss vdd vdd _103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_102 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_196_ mem_left_track_11.DFF_0_.Q vss vss vdd vdd _006_ sky130_fd_sc_hd__clkbuf_1
Xinput24 chany_top_in[2] vss vss vdd vdd net24 sky130_fd_sc_hd__buf_1
X_248_ mem_bottom_track_17.DFF_1_.Q vss vss vdd vdd _118_ sky130_fd_sc_hd__inv_2
X_179_ _000_ vss vss vdd vdd _159_ sky130_fd_sc_hd__clkbuf_1
X_317_ _046_ vss vss vdd vdd _069_ sky130_fd_sc_hd__clkbuf_1
Xinput13 chany_bottom_in[0] vss vss vdd vdd net13 sky130_fd_sc_hd__buf_1
XFILLER_0_19_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold2 mem_left_track_15.DFF_0_.Q vss vss vdd vdd net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_136 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_125 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_496_ mux_bottom_track_9.INVTX1_2_.out _100_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_8_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_136 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_281_ _034_ vss vss vdd vdd _093_ sky130_fd_sc_hd__clkbuf_1
X_350_ net9 vss vss vdd vdd mux_bottom_track_9.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_479_ mux_bottom_track_1.INVTX1_1_.out _083_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_89 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ mux_left_track_13.mux_l1_in_0_.TGATE_0_.out _152_ vss vss vdd vdd mux_left_track_13.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XTAP_56 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_51 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_402_ clknet_2_2__leaf_prog_clk net105 vss vss vdd vdd mem_bottom_track_17.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_40 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_333_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _060_ sky130_fd_sc_hd__inv_2
X_264_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _029_ sky130_fd_sc_hd__clkbuf_1
X_195_ mem_left_track_11.DFF_0_.Q vss vss vdd vdd _149_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_114 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput25 chany_top_in[3] vss vss vdd vdd net25 sky130_fd_sc_hd__clkbuf_1
X_247_ _023_ vss vss vdd vdd _112_ sky130_fd_sc_hd__clkbuf_1
X_316_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _046_ sky130_fd_sc_hd__clkbuf_1
Xinput14 chany_bottom_in[1] vss vss vdd vdd net14 sky130_fd_sc_hd__buf_1
X_178_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _000_ sky130_fd_sc_hd__clkbuf_1
Xhold3 mem_left_track_15.DFF_1_.Q vss vss vdd vdd net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_94 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_60 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_495_ mux_bottom_track_9.INVTX1_4_.out _099_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_71 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_280_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _034_ sky130_fd_sc_hd__clkbuf_1
X_478_ mux_bottom_track_1.INVTX1_3_.out _082_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_547_ mux_left_track_13.INVTX1_1_.out _151_ vss vss vdd vdd mux_left_track_13.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_57 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_26_60 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_52 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_263_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _108_ sky130_fd_sc_hd__inv_2
XPHY_30 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_194_ mem_left_track_11.DFF_1_.Q vss vss vdd vdd _148_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_39 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_332_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _062_ sky130_fd_sc_hd__inv_2
X_401_ clknet_2_1__leaf_prog_clk net87 vss vss vdd vdd mem_top_track_16.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_126 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xinput26 chany_top_in[4] vss vss vdd vdd net26 sky130_fd_sc_hd__buf_1
X_246_ mem_bottom_track_17.DFF_2_.Q vss vss vdd vdd _023_ sky130_fd_sc_hd__clkbuf_1
X_177_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _161_ sky130_fd_sc_hd__inv_2
X_315_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _075_ sky130_fd_sc_hd__inv_2
Xinput15 chany_bottom_in[2] vss vss vdd vdd net15 sky130_fd_sc_hd__buf_1
X_229_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold4 mem_left_track_13.DFF_0_.Q vss vss vdd vdd net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_494_ mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out _098_ vss vss vdd vdd mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_116 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_477_ mux_bottom_track_1.INVTX1_5_.out _081_ vss vss vdd vdd mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_58 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ net75 _150_ vss vss vdd vdd mux_left_track_13.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
XFILLER_0_26_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_50 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_42 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_31 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_262_ _028_ vss vss vdd vdd _102_ sky130_fd_sc_hd__clkbuf_1
X_400_ clknet_2_0__leaf_prog_clk net101 vss vss vdd vdd mem_top_track_16.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_331_ _051_ vss vss vdd vdd _055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_71 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_193_ _005_ vss vss vdd vdd _150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_12_74 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_529_ mux_left_track_3.INVTX1_0_.out _133_ vss vss vdd vdd mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput27 chany_top_in[5] vss vss vdd vdd net27 sky130_fd_sc_hd__buf_1
X_245_ _022_ vss vss vdd vdd _115_ sky130_fd_sc_hd__clkbuf_1
Xinput16 chany_bottom_in[3] vss vss vdd vdd net16 sky130_fd_sc_hd__clkbuf_1
X_314_ mem_top_track_8.DFF_1_.Q vss vss vdd vdd _073_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_228_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _127_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_74 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold5 mem_left_track_7.DFF_0_.Q vss vss vdd vdd net82 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_117 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_26_106 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_493_ mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.out _097_ vss vss vdd vdd mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_128 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_476_ mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out _080_ vss vss vdd vdd mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_59 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_545_ mux_bottom_track_9.INVTX1_1_.out _149_ vss vss vdd vdd mux_left_track_11.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_54 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_43 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_32 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_261_ mem_bottom_track_1.DFF_0_.D vss vss vdd vdd _028_ sky130_fd_sc_hd__clkbuf_1
X_330_ mem_top_track_0.DFF_2_.Q vss vss vdd vdd _051_ sky130_fd_sc_hd__clkbuf_1
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_192_ mem_left_track_13.DFF_1_.Q vss vss vdd vdd _005_ sky130_fd_sc_hd__clkbuf_1
X_459_ mux_top_track_0.mux_l2_in_0_.TGATE_0_.out _063_ vss vss vdd vdd mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_528_ mux_left_track_3.INVTX1_2_.out _132_ vss vss vdd vdd mux_left_track_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput28 chany_top_in[6] vss vss vdd vdd net28 sky130_fd_sc_hd__buf_1
X_244_ mem_bottom_track_17.DFF_0_.Q vss vss vdd vdd _022_ sky130_fd_sc_hd__clkbuf_1
Xinput17 chany_bottom_in[4] vss vss vdd vdd net17 sky130_fd_sc_hd__buf_1
X_313_ _045_ vss vss vdd vdd _066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_40 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_95 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_227_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _125_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold6 mem_bottom_track_1.DFF_2_.Q vss vss vdd vdd net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_42 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_492_ mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out _096_ vss vss vdd vdd mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_525__70 vss vss vdd vdd net70 _525__70/LO sky130_fd_sc_hd__conb_1
XFILLER_0_26_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_475_ net65 _079_ vss vss vdd vdd mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_544_ mux_left_track_11.mux_l1_in_0_.TGATE_0_.out _148_ vss vss vdd vdd mux_left_track_11.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_55 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_44 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_33 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_260_ _027_ vss vss vdd vdd _105_ sky130_fd_sc_hd__clkbuf_1
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_389_ clknet_2_1__leaf_prog_clk net3 vss vss vdd vdd mem_top_track_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
X_527_ mux_left_track_3.mux_l1_in_0_.TGATE_0_.out _131_ vss vss vdd vdd mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_191_ _004_ vss vss vdd vdd _151_ sky130_fd_sc_hd__clkbuf_1
X_458_ mux_top_track_0.mux_l1_in_2_.TGATE_0_.out _062_ vss vss vdd vdd mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput29 chany_top_in[7] vss vss vdd vdd net29 sky130_fd_sc_hd__clkbuf_1
X_243_ mem_bottom_track_17.DFF_0_.Q vss vss vdd vdd _120_ sky130_fd_sc_hd__inv_2
Xinput18 chany_bottom_in[5] vss vss vdd vdd net18 sky130_fd_sc_hd__buf_1
X_312_ mem_top_track_16.DFF_0_.D vss vss vdd vdd _045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_226_ _016_ vss vss vdd vdd _129_ sky130_fd_sc_hd__clkbuf_1
Xhold7 mem_top_track_0.DFF_2_.Q vss vss vdd vdd net84 sky130_fd_sc_hd__dlygate4sd3_1
X_209_ _010_ vss vss vdd vdd _139_ sky130_fd_sc_hd__clkbuf_1
X_491_ mux_bottom_track_9.INVTX1_1_.out _095_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_108 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_22_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_22_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_474_ mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out _078_ vss vss vdd vdd mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_543_ mux_left_track_11.INVTX1_1_.out _147_ vss vss vdd vdd mux_left_track_11.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_26_75 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_13_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_63 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_45 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_34 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_190_ mem_left_track_13.DFF_0_.Q vss vss vdd vdd _004_ sky130_fd_sc_hd__clkbuf_1
X_526_ mux_left_track_3.INVTX1_1_.out _130_ vss vss vdd vdd mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_388_ clknet_2_1__leaf_prog_clk net112 vss vss vdd vdd mem_top_track_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_457_ mux_top_track_0.mux_l1_in_0_.TGATE_0_.out _061_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_114 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_242_ _021_ vss vss vdd vdd _114_ sky130_fd_sc_hd__clkbuf_1
Xinput19 chany_bottom_in[6] vss vss vdd vdd net19 sky130_fd_sc_hd__buf_1
XFILLER_0_5_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_311_ _044_ vss vss vdd vdd _070_ sky130_fd_sc_hd__clkbuf_1
X_509_ net68 _113_ vss vss vdd vdd mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_225_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _016_ sky130_fd_sc_hd__clkbuf_1
Xhold8 mem_left_track_11.DFF_0_.D vss vss vdd vdd net85 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_208_ mem_left_track_7.DFF_0_.Q vss vss vdd vdd _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_43 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_32 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_534__72 vss vss vdd vdd net72 _534__72/LO sky130_fd_sc_hd__conb_1
X_490_ mux_bottom_track_9.INVTX1_3_.out _094_ vss vss vdd vdd mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_11 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_473_ mux_top_track_8.INVTX1_0_.out _077_ vss vss vdd vdd mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_542_ net74 _146_ vss vss vdd vdd mux_left_track_11.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_26_98 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_46 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_456_ mux_bottom_track_17.INVTX1_3_.out _060_ vss vss vdd vdd mux_top_track_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_387_ clknet_2_1__leaf_prog_clk net109 vss vss vdd vdd mem_top_track_0.DFF_2_.Q sky130_fd_sc_hd__dfxtp_1
X_525_ net70 _129_ vss vss vdd vdd mux_left_track_3.mux_l1_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_310_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _044_ sky130_fd_sc_hd__clkbuf_1
X_439_ net27 vss vss vdd vdd net51 sky130_fd_sc_hd__clkbuf_1
X_508_ mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out _112_ vss vss vdd vdd mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_241_ mem_bottom_track_17.DFF_1_.Q vss vss vdd vdd _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_224_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _132_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_77 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xhold9 mem_left_track_3.DFF_1_.Q vss vss vdd vdd net86 sky130_fd_sc_hd__dlygate4sd3_1
X_207_ mem_left_track_7.DFF_0_.Q vss vss vdd vdd _141_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_99 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_0_88 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_0_11 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_23 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_541_ mux_bottom_track_17.INVTX1_1_.out _145_ vss vss vdd vdd mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_472_ mux_left_track_11.INVTX1_1_.out _076_ vss vss vdd vdd mux_top_track_8.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_26_11 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_13_124 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_9_129 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_47 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_386_ net35 vss vss vdd vdd _160_ sky130_fd_sc_hd__inv_2
X_524_ mux_left_track_3.mux_l1_in_1_.TGATE_0_.out _128_ vss vss vdd vdd mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_455_ net63 _059_ vss vss vdd vdd mux_top_track_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_240_ _020_ vss vss vdd vdd _116_ sky130_fd_sc_hd__clkbuf_1
X_438_ net28 vss vss vdd vdd net52 sky130_fd_sc_hd__clkbuf_1
X_369_ net31 vss vss vdd vdd mux_left_track_3.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_0_3_44 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_507_ mux_left_track_7.INVTX1_0_.out _111_ vss vss vdd vdd mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_223_ _015_ vss vss vdd vdd _128_ sky130_fd_sc_hd__clkbuf_1
X_206_ mem_left_track_7.DFF_1_.Q vss vss vdd vdd _140_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_35 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_471_ mux_bottom_track_9.INVTX1_4_.out _075_ vss vss vdd vdd mux_top_track_8.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_540_ mux_left_track_9.mux_l1_in_0_.TGATE_0_.out _144_ vss vss vdd vdd mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_26_89 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_48 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_37 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_136 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_385_ net29 vss vss vdd vdd mux_left_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_523_ mux_bottom_track_1.INVTX1_0_.out _127_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_454_ mux_top_track_0.mux_l1_in_1_.TGATE_0_.out _058_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_5_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_299_ _040_ vss vss vdd vdd _081_ sky130_fd_sc_hd__clkbuf_1
X_506_ mux_bottom_track_1.INVTX1_3_.out _110_ vss vss vdd vdd mux_top_track_16.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_368_ net13 vss vss vdd vdd mux_left_track_3.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_222_ mem_left_track_3.DFF_1_.Q vss vss vdd vdd _015_ sky130_fd_sc_hd__clkbuf_1
X_205_ _009_ vss vss vdd vdd _142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_88 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_16_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_470_ mux_top_track_8.mux_l1_in_0_.TGATE_0_.out _074_ vss vss vdd vdd mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_49 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_38 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_12 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_23 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_522_ mux_left_track_1.INVTX1_2_.out _126_ vss vss vdd vdd mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_453_ mux_bottom_track_17.INVTX1_4_.out _057_ vss vss vdd vdd mux_top_track_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_384_ mux_left_track_17.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net44 sky130_fd_sc_hd__inv_2
X_298_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _040_ sky130_fd_sc_hd__clkbuf_1
X_367_ net16 vss vss vdd vdd mux_left_track_3.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_505_ mux_top_track_16.mux_l1_in_0_.TGATE_0_.out _109_ vss vss vdd vdd mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_221_ _014_ vss vss vdd vdd _130_ sky130_fd_sc_hd__clkbuf_1
X_419_ clknet_2_2__leaf_prog_clk net79 vss vss vdd vdd mem_left_track_15.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_204_ mem_left_track_11.DFF_0_.D vss vss vdd vdd _009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_124 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_90 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_28 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_383_ net30 vss vss vdd vdd mux_left_track_15.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XPHY_39 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_521_ mux_left_track_1.mux_l1_in_0_.TGATE_0_.out _125_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_452_ mux_bottom_track_17.INVTX1_2_.out _056_ vss vss vdd vdd mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xoutput60 net60 vss vss vdd vdd chany_top_out[6] sky130_fd_sc_hd__buf_2
XTAP_130 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_297_ mem_bottom_track_1.DFF_0_.Q vss vss vdd vdd _087_ sky130_fd_sc_hd__inv_2
X_504_ mux_bottom_track_1.INVTX1_5_.out _108_ vss vss vdd vdd mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_116 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_366_ mux_left_track_3.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net37 sky130_fd_sc_hd__inv_2
XFILLER_0_18_37 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_220_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _014_ sky130_fd_sc_hd__clkbuf_1
X_349_ mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net49 sky130_fd_sc_hd__inv_2
X_418_ clknet_2_0__leaf_prog_clk net89 vss vss vdd vdd mem_left_track_13.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_203_ _008_ vss vss vdd vdd _143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_24 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_136 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_26_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_520_ mux_left_track_1.INVTX1_1_.out _124_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_81 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput50 net50 vss vss vdd vdd chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vss vss vdd vdd chany_top_out[7] sky130_fd_sc_hd__clkbuf_4
X_382_ mux_left_track_15.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net43 sky130_fd_sc_hd__inv_2
X_451_ mux_top_track_0.mux_l2_in_1_.TGATE_0_.out _055_ vss vss vdd vdd mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XTAP_120 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_365_ net32 vss vss vdd vdd mux_left_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_296_ mem_bottom_track_1.DFF_1_.Q vss vss vdd vdd _085_ sky130_fd_sc_hd__inv_2
X_503_ mux_top_track_16.mux_l2_in_0_.TGATE_0_.out _107_ vss vss vdd vdd mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_2_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_348_ net11 vss vss vdd vdd mux_bottom_track_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_279_ mem_bottom_track_9.DFF_0_.Q vss vss vdd vdd _099_ sky130_fd_sc_hd__inv_2
X_417_ clknet_2_2__leaf_prog_clk net81 vss vss vdd vdd mem_left_track_13.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_546__75 vss vss vdd vdd net75 _546__75/LO sky130_fd_sc_hd__conb_1
X_202_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_455__63 vss vss vdd vdd net63 _455__63/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_137 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_22_107 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_59 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput51 net51 vss vss vdd vdd chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vss vss vdd vdd chany_top_out[8] sky130_fd_sc_hd__buf_2
X_381_ net19 vss vss vdd vdd mux_left_track_13.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xoutput40 net40 vss vss vdd vdd chanx_left_out[4] sky130_fd_sc_hd__clkbuf_4
X_450_ mux_left_track_3.INVTX1_0_.out _054_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_121 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_23_17 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_502_ mux_left_track_13.INVTX1_1_.out _106_ vss vss vdd vdd mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_3 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_364_ net25 vss vss vdd vdd mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_295_ _039_ vss vss vdd vdd _078_ sky130_fd_sc_hd__clkbuf_1
X_278_ mem_bottom_track_9.DFF_1_.Q vss vss vdd vdd _097_ sky130_fd_sc_hd__inv_2
X_347_ net22 vss vss vdd vdd mux_bottom_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_0_3 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_416_ clknet_2_0__leaf_prog_clk net85 vss vss vdd vdd mem_left_track_11.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_71 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_201_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _145_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_60 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_37 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_19_124 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_21_83 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_530__71 vss vss vdd vdd net71 _530__71/LO sky130_fd_sc_hd__conb_1
XFILLER_0_26_17 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput52 net52 vss vss vdd vdd chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_12_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput41 net41 vss vss vdd vdd chanx_left_out[5] sky130_fd_sc_hd__clkbuf_4
X_380_ mux_left_track_13.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net42 sky130_fd_sc_hd__inv_2
XTAP_122 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

