magic
tech sky130A
magscale 1 2
timestamp 1708041394
<< obsli1 >>
rect 1104 2159 14812 21777
<< obsm1 >>
rect 566 1980 15350 22160
<< metal2 >>
rect 938 23200 994 24000
rect 1674 23200 1730 24000
rect 2410 23200 2466 24000
rect 3146 23200 3202 24000
rect 3882 23200 3938 24000
rect 4618 23200 4674 24000
rect 5354 23200 5410 24000
rect 6090 23200 6146 24000
rect 6826 23200 6882 24000
rect 7562 23200 7618 24000
rect 8298 23200 8354 24000
rect 9034 23200 9090 24000
rect 9770 23200 9826 24000
rect 10506 23200 10562 24000
rect 11242 23200 11298 24000
rect 11978 23200 12034 24000
rect 12714 23200 12770 24000
rect 13450 23200 13506 24000
rect 14186 23200 14242 24000
rect 14922 23200 14978 24000
rect 570 0 626 800
rect 1306 0 1362 800
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
<< obsm2 >>
rect 572 23144 882 23338
rect 1050 23144 1618 23338
rect 1786 23144 2354 23338
rect 2522 23144 3090 23338
rect 3258 23144 3826 23338
rect 3994 23144 4562 23338
rect 4730 23144 5298 23338
rect 5466 23144 6034 23338
rect 6202 23144 6770 23338
rect 6938 23144 7506 23338
rect 7674 23144 8242 23338
rect 8410 23144 8978 23338
rect 9146 23144 9714 23338
rect 9882 23144 10450 23338
rect 10618 23144 11186 23338
rect 11354 23144 11922 23338
rect 12090 23144 12658 23338
rect 12826 23144 13394 23338
rect 13562 23144 14130 23338
rect 14298 23144 14866 23338
rect 15034 23144 15344 23338
rect 572 856 15344 23144
rect 682 303 1250 856
rect 1418 303 1986 856
rect 2154 303 2722 856
rect 2890 303 3458 856
rect 3626 303 4194 856
rect 4362 303 4930 856
rect 5098 303 5666 856
rect 5834 303 6402 856
rect 6570 303 7138 856
rect 7306 303 7874 856
rect 8042 303 8610 856
rect 8778 303 9346 856
rect 9514 303 10082 856
rect 10250 303 10818 856
rect 10986 303 11554 856
rect 11722 303 12290 856
rect 12458 303 13026 856
rect 13194 303 13762 856
rect 13930 303 14498 856
rect 14666 303 15344 856
<< metal3 >>
rect 0 23128 800 23248
rect 15200 23128 16000 23248
rect 0 22040 800 22160
rect 15200 22040 16000 22160
rect 0 20952 800 21072
rect 15200 20952 16000 21072
rect 0 19864 800 19984
rect 15200 19864 16000 19984
rect 0 18776 800 18896
rect 15200 18776 16000 18896
rect 0 17688 800 17808
rect 15200 17688 16000 17808
rect 0 16600 800 16720
rect 15200 16600 16000 16720
rect 0 15512 800 15632
rect 15200 15512 16000 15632
rect 0 14424 800 14544
rect 15200 14424 16000 14544
rect 0 13336 800 13456
rect 15200 13336 16000 13456
rect 0 12248 800 12368
rect 15200 12248 16000 12368
rect 0 11160 800 11280
rect 15200 11160 16000 11280
rect 0 10072 800 10192
rect 15200 10072 16000 10192
rect 0 8984 800 9104
rect 15200 8984 16000 9104
rect 0 7896 800 8016
rect 15200 7896 16000 8016
rect 0 6808 800 6928
rect 15200 6808 16000 6928
rect 0 5720 800 5840
rect 15200 5720 16000 5840
rect 0 4632 800 4752
rect 15200 4632 16000 4752
rect 0 3544 800 3664
rect 15200 3544 16000 3664
rect 0 2456 800 2576
rect 15200 2456 16000 2576
rect 0 1368 800 1488
rect 15200 1368 16000 1488
rect 15200 280 16000 400
<< obsm3 >>
rect 880 23048 15120 23221
rect 798 22240 15200 23048
rect 880 21960 15120 22240
rect 798 21152 15200 21960
rect 880 20872 15120 21152
rect 798 20064 15200 20872
rect 880 19784 15120 20064
rect 798 18976 15200 19784
rect 880 18696 15120 18976
rect 798 17888 15200 18696
rect 880 17608 15120 17888
rect 798 16800 15200 17608
rect 880 16520 15120 16800
rect 798 15712 15200 16520
rect 880 15432 15120 15712
rect 798 14624 15200 15432
rect 880 14344 15120 14624
rect 798 13536 15200 14344
rect 880 13256 15120 13536
rect 798 12448 15200 13256
rect 880 12168 15120 12448
rect 798 11360 15200 12168
rect 880 11080 15120 11360
rect 798 10272 15200 11080
rect 880 9992 15120 10272
rect 798 9184 15200 9992
rect 880 8904 15120 9184
rect 798 8096 15200 8904
rect 880 7816 15120 8096
rect 798 7008 15200 7816
rect 880 6728 15120 7008
rect 798 5920 15200 6728
rect 880 5640 15120 5920
rect 798 4832 15200 5640
rect 880 4552 15120 4832
rect 798 3744 15200 4552
rect 880 3464 15120 3744
rect 798 2656 15200 3464
rect 880 2376 15120 2656
rect 798 1568 15200 2376
rect 880 1288 15120 1568
rect 798 480 15200 1288
rect 798 307 15120 480
<< metal4 >>
rect 2657 2128 2977 21808
rect 4370 2128 4690 21808
rect 6084 2128 6404 21808
rect 7797 2128 8117 21808
rect 9511 2128 9831 21808
rect 11224 2128 11544 21808
rect 12938 2128 13258 21808
rect 14651 2128 14971 21808
<< obsm4 >>
rect 1899 2048 2577 20773
rect 3057 2048 4290 20773
rect 4770 2048 6004 20773
rect 6484 2048 7717 20773
rect 8197 2048 9431 20773
rect 9911 2048 11144 20773
rect 11624 2048 11901 20773
rect 1899 1803 11901 2048
<< labels >>
rlabel metal2 s 7930 0 7986 800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 1 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 2 nsew signal input
rlabel metal3 s 15200 22040 16000 22160 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 15200 23128 16000 23248 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 chanx_left_in[0]
port 5 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[1]
port 6 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 chanx_left_in[2]
port 7 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 8 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[4]
port 9 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 chanx_left_in[5]
port 10 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[6]
port 11 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[7]
port 12 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[8]
port 13 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[0]
port 14 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[1]
port 15 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 chanx_left_out[2]
port 16 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 chanx_left_out[3]
port 17 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[4]
port 18 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 chanx_left_out[5]
port 19 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 chanx_left_out[6]
port 20 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[7]
port 21 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 chanx_left_out[8]
port 22 nsew signal output
rlabel metal3 s 15200 280 16000 400 6 chanx_right_in[0]
port 23 nsew signal input
rlabel metal3 s 15200 1368 16000 1488 6 chanx_right_in[1]
port 24 nsew signal input
rlabel metal3 s 15200 2456 16000 2576 6 chanx_right_in[2]
port 25 nsew signal input
rlabel metal3 s 15200 3544 16000 3664 6 chanx_right_in[3]
port 26 nsew signal input
rlabel metal3 s 15200 4632 16000 4752 6 chanx_right_in[4]
port 27 nsew signal input
rlabel metal3 s 15200 5720 16000 5840 6 chanx_right_in[5]
port 28 nsew signal input
rlabel metal3 s 15200 6808 16000 6928 6 chanx_right_in[6]
port 29 nsew signal input
rlabel metal3 s 15200 7896 16000 8016 6 chanx_right_in[7]
port 30 nsew signal input
rlabel metal3 s 15200 8984 16000 9104 6 chanx_right_in[8]
port 31 nsew signal input
rlabel metal3 s 15200 10072 16000 10192 6 chanx_right_out[0]
port 32 nsew signal output
rlabel metal3 s 15200 11160 16000 11280 6 chanx_right_out[1]
port 33 nsew signal output
rlabel metal3 s 15200 12248 16000 12368 6 chanx_right_out[2]
port 34 nsew signal output
rlabel metal3 s 15200 13336 16000 13456 6 chanx_right_out[3]
port 35 nsew signal output
rlabel metal3 s 15200 14424 16000 14544 6 chanx_right_out[4]
port 36 nsew signal output
rlabel metal3 s 15200 15512 16000 15632 6 chanx_right_out[5]
port 37 nsew signal output
rlabel metal3 s 15200 16600 16000 16720 6 chanx_right_out[6]
port 38 nsew signal output
rlabel metal3 s 15200 17688 16000 17808 6 chanx_right_out[7]
port 39 nsew signal output
rlabel metal3 s 15200 18776 16000 18896 6 chanx_right_out[8]
port 40 nsew signal output
rlabel metal2 s 570 0 626 800 6 chany_bottom_in[0]
port 41 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 chany_bottom_in[1]
port 42 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 chany_bottom_in[2]
port 43 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_in[3]
port 44 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_in[4]
port 45 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[5]
port 46 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[6]
port 47 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[7]
port 48 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[8]
port 49 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_out[0]
port 50 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_out[1]
port 51 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_out[2]
port 52 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_out[3]
port 53 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_out[4]
port 54 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_out[5]
port 55 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[6]
port 56 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[7]
port 57 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[8]
port 58 nsew signal output
rlabel metal2 s 938 23200 994 24000 6 chany_top_in[0]
port 59 nsew signal input
rlabel metal2 s 1674 23200 1730 24000 6 chany_top_in[1]
port 60 nsew signal input
rlabel metal2 s 2410 23200 2466 24000 6 chany_top_in[2]
port 61 nsew signal input
rlabel metal2 s 3146 23200 3202 24000 6 chany_top_in[3]
port 62 nsew signal input
rlabel metal2 s 3882 23200 3938 24000 6 chany_top_in[4]
port 63 nsew signal input
rlabel metal2 s 4618 23200 4674 24000 6 chany_top_in[5]
port 64 nsew signal input
rlabel metal2 s 5354 23200 5410 24000 6 chany_top_in[6]
port 65 nsew signal input
rlabel metal2 s 6090 23200 6146 24000 6 chany_top_in[7]
port 66 nsew signal input
rlabel metal2 s 6826 23200 6882 24000 6 chany_top_in[8]
port 67 nsew signal input
rlabel metal2 s 7562 23200 7618 24000 6 chany_top_out[0]
port 68 nsew signal output
rlabel metal2 s 8298 23200 8354 24000 6 chany_top_out[1]
port 69 nsew signal output
rlabel metal2 s 9034 23200 9090 24000 6 chany_top_out[2]
port 70 nsew signal output
rlabel metal2 s 9770 23200 9826 24000 6 chany_top_out[3]
port 71 nsew signal output
rlabel metal2 s 10506 23200 10562 24000 6 chany_top_out[4]
port 72 nsew signal output
rlabel metal2 s 11242 23200 11298 24000 6 chany_top_out[5]
port 73 nsew signal output
rlabel metal2 s 11978 23200 12034 24000 6 chany_top_out[6]
port 74 nsew signal output
rlabel metal2 s 12714 23200 12770 24000 6 chany_top_out[7]
port 75 nsew signal output
rlabel metal2 s 13450 23200 13506 24000 6 chany_top_out[8]
port 76 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 77 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 78 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 prog_clk
port 79 nsew signal input
rlabel metal3 s 15200 19864 16000 19984 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 80 nsew signal input
rlabel metal3 s 15200 20952 16000 21072 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 81 nsew signal input
rlabel metal2 s 14186 23200 14242 24000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 82 nsew signal input
rlabel metal2 s 14922 23200 14978 24000 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 83 nsew signal input
rlabel metal4 s 2657 2128 2977 21808 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 21808 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 21808 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 21808 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 21808 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 21808 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 21808 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 21808 6 vss
port 85 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1506748
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_1__1_/runs/24_02_15_17_55/results/signoff/sb_1__1_.magic.gds
string GDS_START 111472
<< end >>

