magic
tech sky130A
magscale 1 2
timestamp 1708041521
<< obsli1 >>
rect 1104 2159 14812 13617
<< obsm1 >>
rect 934 1924 15074 13648
<< metal2 >>
rect 1030 15200 1086 16000
rect 2410 15200 2466 16000
rect 3790 15200 3846 16000
rect 5170 15200 5226 16000
rect 6550 15200 6606 16000
rect 7930 15200 7986 16000
rect 9310 15200 9366 16000
rect 10690 15200 10746 16000
rect 12070 15200 12126 16000
rect 13450 15200 13506 16000
rect 14830 15200 14886 16000
rect 2502 0 2558 800
rect 4066 0 4122 800
rect 5630 0 5686 800
rect 7194 0 7250 800
rect 8758 0 8814 800
rect 10322 0 10378 800
rect 11886 0 11942 800
rect 13450 0 13506 800
rect 15014 0 15070 800
<< obsm2 >>
rect 938 15144 974 15314
rect 1142 15144 2354 15314
rect 2522 15144 3734 15314
rect 3902 15144 5114 15314
rect 5282 15144 6494 15314
rect 6662 15144 7874 15314
rect 8042 15144 9254 15314
rect 9422 15144 10634 15314
rect 10802 15144 12014 15314
rect 12182 15144 13394 15314
rect 13562 15144 14774 15314
rect 14942 15144 15068 15314
rect 938 856 15068 15144
rect 938 734 2446 856
rect 2614 734 4010 856
rect 4178 734 5574 856
rect 5742 734 7138 856
rect 7306 734 8702 856
rect 8870 734 10266 856
rect 10434 734 11830 856
rect 11998 734 13394 856
rect 13562 734 14958 856
<< metal3 >>
rect 15200 14696 16000 14816
rect 0 14424 800 14544
rect 0 13336 800 13456
rect 15200 13336 16000 13456
rect 0 12248 800 12368
rect 15200 11976 16000 12096
rect 0 11160 800 11280
rect 15200 10616 16000 10736
rect 0 10072 800 10192
rect 15200 9256 16000 9376
rect 0 8984 800 9104
rect 0 7896 800 8016
rect 15200 7896 16000 8016
rect 0 6808 800 6928
rect 15200 6536 16000 6656
rect 0 5720 800 5840
rect 15200 5176 16000 5296
rect 0 4632 800 4752
rect 15200 3816 16000 3936
rect 0 3544 800 3664
rect 0 2456 800 2576
rect 15200 2456 16000 2576
rect 15200 1096 16000 1216
<< obsm3 >>
rect 798 14624 15120 14789
rect 880 14616 15120 14624
rect 880 14344 15210 14616
rect 798 13536 15210 14344
rect 880 13256 15120 13536
rect 798 12448 15210 13256
rect 880 12176 15210 12448
rect 880 12168 15120 12176
rect 798 11896 15120 12168
rect 798 11360 15210 11896
rect 880 11080 15210 11360
rect 798 10816 15210 11080
rect 798 10536 15120 10816
rect 798 10272 15210 10536
rect 880 9992 15210 10272
rect 798 9456 15210 9992
rect 798 9184 15120 9456
rect 880 9176 15120 9184
rect 880 8904 15210 9176
rect 798 8096 15210 8904
rect 880 7816 15120 8096
rect 798 7008 15210 7816
rect 880 6736 15210 7008
rect 880 6728 15120 6736
rect 798 6456 15120 6728
rect 798 5920 15210 6456
rect 880 5640 15210 5920
rect 798 5376 15210 5640
rect 798 5096 15120 5376
rect 798 4832 15210 5096
rect 880 4552 15210 4832
rect 798 4016 15210 4552
rect 798 3744 15120 4016
rect 880 3736 15120 3744
rect 880 3464 15210 3736
rect 798 2656 15210 3464
rect 880 2376 15120 2656
rect 798 1296 15210 2376
rect 798 1123 15120 1296
<< metal4 >>
rect 2657 2128 2977 13648
rect 4370 2128 4690 13648
rect 6084 2128 6404 13648
rect 7797 2128 8117 13648
rect 9511 2128 9831 13648
rect 11224 2128 11544 13648
rect 12938 2128 13258 13648
rect 14651 2128 14971 13648
<< labels >>
rlabel metal3 s 15200 13336 16000 13456 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 15200 14696 16000 14816 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 15200 1096 16000 1216 6 chanx_left_in[0]
port 3 nsew signal input
rlabel metal3 s 15200 2456 16000 2576 6 chanx_left_in[1]
port 4 nsew signal input
rlabel metal3 s 15200 3816 16000 3936 6 chanx_left_in[2]
port 5 nsew signal input
rlabel metal3 s 15200 5176 16000 5296 6 chanx_left_in[3]
port 6 nsew signal input
rlabel metal3 s 15200 6536 16000 6656 6 chanx_left_in[4]
port 7 nsew signal input
rlabel metal3 s 15200 7896 16000 8016 6 chanx_left_in[5]
port 8 nsew signal input
rlabel metal3 s 15200 9256 16000 9376 6 chanx_left_in[6]
port 9 nsew signal input
rlabel metal3 s 15200 10616 16000 10736 6 chanx_left_in[7]
port 10 nsew signal input
rlabel metal3 s 15200 11976 16000 12096 6 chanx_left_in[8]
port 11 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 chanx_left_out[0]
port 12 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 chanx_left_out[1]
port 13 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 chanx_left_out[2]
port 14 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 chanx_left_out[3]
port 15 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 chanx_left_out[4]
port 16 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 chanx_left_out[5]
port 17 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 chanx_left_out[6]
port 18 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 chanx_left_out[7]
port 19 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 chanx_left_out[8]
port 20 nsew signal output
rlabel metal2 s 1030 15200 1086 16000 6 chany_top_in[0]
port 21 nsew signal input
rlabel metal2 s 2410 15200 2466 16000 6 chany_top_in[1]
port 22 nsew signal input
rlabel metal2 s 3790 15200 3846 16000 6 chany_top_in[2]
port 23 nsew signal input
rlabel metal2 s 5170 15200 5226 16000 6 chany_top_in[3]
port 24 nsew signal input
rlabel metal2 s 6550 15200 6606 16000 6 chany_top_in[4]
port 25 nsew signal input
rlabel metal2 s 7930 15200 7986 16000 6 chany_top_in[5]
port 26 nsew signal input
rlabel metal2 s 9310 15200 9366 16000 6 chany_top_in[6]
port 27 nsew signal input
rlabel metal2 s 10690 15200 10746 16000 6 chany_top_in[7]
port 28 nsew signal input
rlabel metal2 s 12070 15200 12126 16000 6 chany_top_in[8]
port 29 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 chany_top_out[0]
port 30 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 chany_top_out[1]
port 31 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 chany_top_out[2]
port 32 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 chany_top_out[3]
port 33 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 chany_top_out[4]
port 34 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 chany_top_out[5]
port 35 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 chany_top_out[6]
port 36 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 chany_top_out[7]
port 37 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 chany_top_out[8]
port 38 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 39 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 40 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 prog_clk
port 41 nsew signal input
rlabel metal2 s 13450 15200 13506 16000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 42 nsew signal input
rlabel metal2 s 14830 15200 14886 16000 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 43 nsew signal input
rlabel metal4 s 2657 2128 2977 13648 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 13648 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 13648 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 13648 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 13648 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 13648 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 13648 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 13648 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 16000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 382174
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_8__0_/runs/24_02_15_17_58/results/signoff/sb_8__0_.magic.gds
string GDS_START 85502
<< end >>

