magic
tech sky130A
magscale 1 2
timestamp 1708041323
<< viali >>
rect 6561 17289 6595 17323
rect 7481 17289 7515 17323
rect 7849 17289 7883 17323
rect 9321 17289 9355 17323
rect 9965 17289 9999 17323
rect 10701 17289 10735 17323
rect 11621 17289 11655 17323
rect 12265 17289 12299 17323
rect 13001 17289 13035 17323
rect 13829 17289 13863 17323
rect 10241 17221 10275 17255
rect 1501 17153 1535 17187
rect 1777 17153 1811 17187
rect 2053 17153 2087 17187
rect 2605 17153 2639 17187
rect 2881 17153 2915 17187
rect 3341 17153 3375 17187
rect 3617 17153 3651 17187
rect 5457 17153 5491 17187
rect 5733 17153 5767 17187
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 6653 17153 6687 17187
rect 6929 17153 6963 17187
rect 7389 17153 7423 17187
rect 7665 17153 7699 17187
rect 7765 17153 7799 17187
rect 8217 17153 8251 17187
rect 9229 17153 9263 17187
rect 10977 17153 11011 17187
rect 11897 17153 11931 17187
rect 12173 17153 12207 17187
rect 12909 17153 12943 17187
rect 13553 17153 13587 17187
rect 14105 17153 14139 17187
rect 2513 17085 2547 17119
rect 3249 17085 3283 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4721 17085 4755 17119
rect 8033 17085 8067 17119
rect 3433 17017 3467 17051
rect 5641 17017 5675 17051
rect 7297 17017 7331 17051
rect 1685 16949 1719 16983
rect 1961 16949 1995 16983
rect 2237 16949 2271 16983
rect 2789 16949 2823 16983
rect 3065 16949 3099 16983
rect 4537 16949 4571 16983
rect 5273 16949 5307 16983
rect 5825 16949 5859 16983
rect 6009 16949 6043 16983
rect 6745 16949 6779 16983
rect 7113 16949 7147 16983
rect 8493 16949 8527 16983
rect 14197 16949 14231 16983
rect 3341 16745 3375 16779
rect 4537 16745 4571 16779
rect 8677 16745 8711 16779
rect 11713 16745 11747 16779
rect 11897 16745 11931 16779
rect 12633 16745 12667 16779
rect 12909 16745 12943 16779
rect 13369 16745 13403 16779
rect 13829 16745 13863 16779
rect 2789 16677 2823 16711
rect 7297 16677 7331 16711
rect 3893 16609 3927 16643
rect 4077 16609 4111 16643
rect 5641 16609 5675 16643
rect 6377 16609 6411 16643
rect 9689 16609 9723 16643
rect 10149 16609 10183 16643
rect 1409 16541 1443 16575
rect 1685 16541 1719 16575
rect 1961 16541 1995 16575
rect 2237 16541 2271 16575
rect 2605 16541 2639 16575
rect 2881 16541 2915 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 7113 16541 7147 16575
rect 7397 16541 7431 16575
rect 7665 16541 7699 16575
rect 8585 16541 8619 16575
rect 10609 16541 10643 16575
rect 10793 16541 10827 16575
rect 11345 16541 11379 16575
rect 11621 16541 11655 16575
rect 12081 16541 12115 16575
rect 12357 16541 12391 16575
rect 12449 16541 12483 16575
rect 12725 16541 12759 16575
rect 13185 16541 13219 16575
rect 14105 16541 14139 16575
rect 5733 16473 5767 16507
rect 6285 16473 6319 16507
rect 9045 16473 9079 16507
rect 9137 16473 9171 16507
rect 9873 16473 9907 16507
rect 9965 16473 9999 16507
rect 11437 16473 11471 16507
rect 13553 16473 13587 16507
rect 1593 16405 1627 16439
rect 1777 16405 1811 16439
rect 2053 16405 2087 16439
rect 2421 16405 2455 16439
rect 2973 16405 3007 16439
rect 3525 16405 3559 16439
rect 5457 16405 5491 16439
rect 7021 16405 7055 16439
rect 7573 16405 7607 16439
rect 8309 16405 8343 16439
rect 11253 16405 11287 16439
rect 12265 16405 12299 16439
rect 14197 16405 14231 16439
rect 2881 16201 2915 16235
rect 4445 16201 4479 16235
rect 6009 16201 6043 16235
rect 9045 16201 9079 16235
rect 9413 16201 9447 16235
rect 10885 16201 10919 16235
rect 11713 16201 11747 16235
rect 13645 16201 13679 16235
rect 14381 16201 14415 16235
rect 4016 16133 4050 16167
rect 4896 16133 4930 16167
rect 6561 16133 6595 16167
rect 8410 16133 8444 16167
rect 9689 16133 9723 16167
rect 14105 16133 14139 16167
rect 1777 16065 1811 16099
rect 2053 16065 2087 16099
rect 2145 16065 2179 16099
rect 4377 16065 4411 16099
rect 8861 16065 8895 16099
rect 9229 16065 9263 16099
rect 10149 16065 10183 16099
rect 10333 16065 10367 16099
rect 10425 16065 10459 16099
rect 10701 16065 10735 16099
rect 11621 16065 11655 16099
rect 13277 16065 13311 16099
rect 13553 16065 13587 16099
rect 2329 15997 2363 16031
rect 4261 15997 4295 16031
rect 4629 15997 4663 16031
rect 6469 15997 6503 16031
rect 6745 15997 6779 16031
rect 8677 15997 8711 16031
rect 11161 15997 11195 16031
rect 12817 15997 12851 16031
rect 1869 15929 1903 15963
rect 2789 15929 2823 15963
rect 7297 15929 7331 15963
rect 1685 15861 1719 15895
rect 10609 15861 10643 15895
rect 13461 15861 13495 15895
rect 2697 15657 2731 15691
rect 4169 15657 4203 15691
rect 5917 15657 5951 15691
rect 8493 15657 8527 15691
rect 9781 15657 9815 15691
rect 10149 15657 10183 15691
rect 13093 15657 13127 15691
rect 4629 15589 4663 15623
rect 5089 15589 5123 15623
rect 12357 15589 12391 15623
rect 3525 15521 3559 15555
rect 5549 15521 5583 15555
rect 8033 15521 8067 15555
rect 8953 15521 8987 15555
rect 10425 15521 10459 15555
rect 11253 15521 11287 15555
rect 12633 15521 12667 15555
rect 2789 15453 2823 15487
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 4261 15453 4295 15487
rect 4813 15453 4847 15487
rect 4905 15453 4939 15487
rect 5273 15453 5307 15487
rect 5733 15453 5767 15487
rect 6285 15453 6319 15487
rect 6552 15453 6586 15487
rect 7849 15453 7883 15487
rect 8585 15453 8619 15487
rect 9689 15453 9723 15487
rect 9965 15453 9999 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 11437 15453 11471 15487
rect 12173 15453 12207 15487
rect 12449 15453 12483 15487
rect 14105 15453 14139 15487
rect 8677 15385 8711 15419
rect 11161 15385 11195 15419
rect 11897 15385 11931 15419
rect 13185 15385 13219 15419
rect 13737 15385 13771 15419
rect 13829 15385 13863 15419
rect 5457 15317 5491 15351
rect 7665 15317 7699 15351
rect 9597 15317 9631 15351
rect 14197 15317 14231 15351
rect 2973 15113 3007 15147
rect 8033 15113 8067 15147
rect 10425 15113 10459 15147
rect 11529 15113 11563 15147
rect 11989 15113 12023 15147
rect 13461 15113 13495 15147
rect 14381 15113 14415 15147
rect 2789 14977 2823 15011
rect 3249 14977 3283 15011
rect 3433 14977 3467 15011
rect 3525 14977 3559 15011
rect 3709 14977 3743 15011
rect 5181 14977 5215 15011
rect 6561 14977 6595 15011
rect 7757 14977 7791 15011
rect 8677 14977 8711 15011
rect 9413 14977 9447 15011
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 14105 14977 14139 15011
rect 14289 14977 14323 15011
rect 3893 14909 3927 14943
rect 6837 14909 6871 14943
rect 7021 14909 7055 14943
rect 9229 14909 9263 14943
rect 10057 14909 10091 14943
rect 12081 14909 12115 14943
rect 12817 14909 12851 14943
rect 13001 14909 13035 14943
rect 3065 14841 3099 14875
rect 7941 14841 7975 14875
rect 4169 14773 4203 14807
rect 5273 14773 5307 14807
rect 6745 14773 6779 14807
rect 7481 14773 7515 14807
rect 8769 14773 8803 14807
rect 9505 14773 9539 14807
rect 11253 14773 11287 14807
rect 12725 14773 12759 14807
rect 13553 14773 13587 14807
rect 4997 14569 5031 14603
rect 6009 14569 6043 14603
rect 8309 14569 8343 14603
rect 10425 14569 10459 14603
rect 13369 14569 13403 14603
rect 13553 14569 13587 14603
rect 14289 14569 14323 14603
rect 3617 14501 3651 14535
rect 5089 14501 5123 14535
rect 7389 14501 7423 14535
rect 4353 14433 4387 14467
rect 5365 14433 5399 14467
rect 5549 14433 5583 14467
rect 6561 14433 6595 14467
rect 6929 14433 6963 14467
rect 7665 14433 7699 14467
rect 8125 14433 8159 14467
rect 9045 14433 9079 14467
rect 1409 14365 1443 14399
rect 3433 14365 3467 14399
rect 4537 14365 4571 14399
rect 4813 14365 4847 14399
rect 5273 14365 5307 14399
rect 6285 14365 6319 14399
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 7481 14365 7515 14399
rect 8493 14365 8527 14399
rect 8769 14365 8803 14399
rect 11630 14365 11664 14399
rect 11897 14365 11931 14399
rect 11989 14365 12023 14399
rect 12256 14365 12290 14399
rect 13645 14365 13679 14399
rect 14473 14365 14507 14399
rect 9312 14297 9346 14331
rect 1593 14229 1627 14263
rect 3893 14229 3927 14263
rect 6193 14229 6227 14263
rect 8677 14229 8711 14263
rect 10517 14229 10551 14263
rect 1685 14025 1719 14059
rect 3249 14025 3283 14059
rect 5825 14025 5859 14059
rect 6101 14025 6135 14059
rect 7849 14025 7883 14059
rect 8217 14025 8251 14059
rect 10333 14025 10367 14059
rect 10609 14025 10643 14059
rect 11345 14025 11379 14059
rect 4445 13957 4479 13991
rect 9330 13957 9364 13991
rect 12072 13957 12106 13991
rect 1409 13889 1443 13923
rect 1869 13889 1903 13923
rect 1961 13889 1995 13923
rect 3065 13889 3099 13923
rect 3341 13889 3375 13923
rect 3433 13889 3467 13923
rect 4077 13889 4111 13923
rect 4353 13889 4387 13923
rect 4905 13889 4939 13923
rect 5181 13889 5215 13923
rect 5365 13889 5399 13923
rect 6017 13889 6051 13923
rect 6644 13889 6678 13923
rect 8033 13889 8067 13923
rect 10149 13889 10183 13923
rect 10425 13889 10459 13923
rect 11713 13889 11747 13923
rect 14473 13889 14507 13923
rect 2145 13821 2179 13855
rect 4261 13821 4295 13855
rect 6377 13821 6411 13855
rect 9597 13821 9631 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 11621 13821 11655 13855
rect 11805 13821 11839 13855
rect 14197 13821 14231 13855
rect 1593 13753 1627 13787
rect 2513 13685 2547 13719
rect 3617 13685 3651 13719
rect 4721 13685 4755 13719
rect 7757 13685 7791 13719
rect 13185 13685 13219 13719
rect 1777 13481 1811 13515
rect 3617 13481 3651 13515
rect 8953 13481 8987 13515
rect 10333 13481 10367 13515
rect 10793 13481 10827 13515
rect 11713 13481 11747 13515
rect 13461 13481 13495 13515
rect 2329 13413 2363 13447
rect 2605 13413 2639 13447
rect 6653 13413 6687 13447
rect 3157 13345 3191 13379
rect 4997 13345 5031 13379
rect 5549 13345 5583 13379
rect 7573 13345 7607 13379
rect 7849 13345 7883 13379
rect 8309 13345 8343 13379
rect 9873 13345 9907 13379
rect 11345 13345 11379 13379
rect 12081 13345 12115 13379
rect 1409 13277 1443 13311
rect 1685 13277 1719 13311
rect 2145 13277 2179 13311
rect 2421 13277 2455 13311
rect 2881 13277 2915 13311
rect 2973 13277 3007 13311
rect 3985 13277 4019 13311
rect 4261 13277 4295 13311
rect 4353 13277 4387 13311
rect 4629 13277 4663 13311
rect 4905 13277 4939 13311
rect 5365 13277 5399 13311
rect 6193 13277 6227 13311
rect 6469 13277 6503 13311
rect 8769 13277 8803 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 11161 13277 11195 13311
rect 6929 13209 6963 13243
rect 7941 13209 7975 13243
rect 8677 13209 8711 13243
rect 12348 13209 12382 13243
rect 1593 13141 1627 13175
rect 2789 13141 2823 13175
rect 3801 13141 3835 13175
rect 4077 13141 4111 13175
rect 4537 13141 4571 13175
rect 4813 13141 4847 13175
rect 6009 13141 6043 13175
rect 6285 13141 6319 13175
rect 7021 13141 7055 13175
rect 13645 13141 13679 13175
rect 2513 12937 2547 12971
rect 9137 12937 9171 12971
rect 9781 12937 9815 12971
rect 10425 12937 10459 12971
rect 4353 12869 4387 12903
rect 5365 12869 5399 12903
rect 7849 12869 7883 12903
rect 1777 12801 1811 12835
rect 1869 12801 1903 12835
rect 4445 12801 4479 12835
rect 6009 12801 6043 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 7297 12801 7331 12835
rect 9873 12801 9907 12835
rect 9965 12801 9999 12835
rect 10241 12801 10275 12835
rect 11345 12801 11379 12835
rect 12541 12801 12575 12835
rect 13185 12801 13219 12835
rect 13369 12801 13403 12835
rect 2053 12733 2087 12767
rect 4629 12733 4663 12767
rect 5273 12733 5307 12767
rect 5549 12733 5583 12767
rect 7113 12733 7147 12767
rect 11161 12733 11195 12767
rect 11529 12733 11563 12767
rect 14197 12733 14231 12767
rect 14473 12733 14507 12767
rect 1685 12665 1719 12699
rect 3065 12665 3099 12699
rect 6193 12665 6227 12699
rect 10149 12665 10183 12699
rect 4813 12597 4847 12631
rect 7021 12597 7055 12631
rect 7481 12597 7515 12631
rect 10977 12597 11011 12631
rect 11897 12597 11931 12631
rect 12633 12597 12667 12631
rect 13461 12597 13495 12631
rect 4445 12393 4479 12427
rect 6009 12393 6043 12427
rect 10885 12393 10919 12427
rect 14105 12393 14139 12427
rect 3525 12325 3559 12359
rect 9137 12325 9171 12359
rect 13277 12325 13311 12359
rect 2605 12257 2639 12291
rect 3801 12257 3835 12291
rect 3985 12257 4019 12291
rect 6377 12257 6411 12291
rect 7941 12257 7975 12291
rect 8309 12257 8343 12291
rect 10057 12257 10091 12291
rect 12265 12257 12299 12291
rect 12541 12257 12575 12291
rect 13829 12257 13863 12291
rect 1593 12189 1627 12223
rect 2789 12189 2823 12223
rect 3433 12189 3467 12223
rect 4721 12189 4755 12223
rect 4997 12189 5031 12223
rect 5273 12189 5307 12223
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 6644 12189 6678 12223
rect 8953 12189 8987 12223
rect 9413 12189 9447 12223
rect 9781 12189 9815 12223
rect 10241 12189 10275 12223
rect 12357 12189 12391 12223
rect 14289 12189 14323 12223
rect 8033 12121 8067 12155
rect 12020 12121 12054 12155
rect 13737 12121 13771 12155
rect 1685 12053 1719 12087
rect 2421 12053 2455 12087
rect 3249 12053 3283 12087
rect 4905 12053 4939 12087
rect 5181 12053 5215 12087
rect 7757 12053 7791 12087
rect 9229 12053 9263 12087
rect 9965 12053 9999 12087
rect 10701 12053 10735 12087
rect 13001 12053 13035 12087
rect 1869 11849 1903 11883
rect 4169 11849 4203 11883
rect 10333 11849 10367 11883
rect 10609 11849 10643 11883
rect 11529 11849 11563 11883
rect 13185 11849 13219 11883
rect 14289 11849 14323 11883
rect 2697 11781 2731 11815
rect 3034 11781 3068 11815
rect 6929 11781 6963 11815
rect 14013 11781 14047 11815
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 2145 11713 2179 11747
rect 4905 11713 4939 11747
rect 5273 11713 5307 11747
rect 8769 11713 8803 11747
rect 9025 11713 9059 11747
rect 10425 11713 10459 11747
rect 11069 11713 11103 11747
rect 11253 11713 11287 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 12072 11713 12106 11747
rect 13461 11713 13495 11747
rect 14473 11713 14507 11747
rect 2789 11645 2823 11679
rect 14105 11645 14139 11679
rect 5089 11577 5123 11611
rect 10149 11577 10183 11611
rect 1593 11509 1627 11543
rect 4353 11509 4387 11543
rect 8217 11509 8251 11543
rect 1409 11305 1443 11339
rect 5641 11305 5675 11339
rect 12357 11305 12391 11339
rect 12633 11305 12667 11339
rect 13553 11305 13587 11339
rect 13829 11305 13863 11339
rect 6469 11237 6503 11271
rect 6929 11237 6963 11271
rect 8769 11237 8803 11271
rect 12173 11237 12207 11271
rect 14197 11237 14231 11271
rect 2789 11169 2823 11203
rect 6745 11169 6779 11203
rect 7571 11169 7605 11203
rect 8401 11169 8435 11203
rect 9137 11169 9171 11203
rect 10149 11169 10183 11203
rect 11345 11169 11379 11203
rect 11621 11169 11655 11203
rect 3985 11101 4019 11135
rect 5089 11101 5123 11135
rect 5457 11101 5491 11135
rect 5549 11101 5583 11135
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 6561 11101 6595 11135
rect 7297 11101 7331 11135
rect 7757 11101 7791 11135
rect 8309 11101 8343 11135
rect 8585 11101 8619 11135
rect 8953 11101 8987 11135
rect 10333 11101 10367 11135
rect 10977 11101 11011 11135
rect 12081 11101 12115 11135
rect 12541 11101 12575 11135
rect 13277 11101 13311 11135
rect 13369 11101 13403 11135
rect 13645 11101 13679 11135
rect 14105 11101 14139 11135
rect 2522 11033 2556 11067
rect 2973 11033 3007 11067
rect 3065 11033 3099 11067
rect 3617 11033 3651 11067
rect 4077 11033 4111 11067
rect 4629 11033 4663 11067
rect 4721 11033 4755 11067
rect 4997 11033 5031 11067
rect 9597 11033 9631 11067
rect 9689 11033 9723 11067
rect 10425 11033 10459 11067
rect 11437 11033 11471 11067
rect 3801 10965 3835 10999
rect 5273 10965 5307 10999
rect 7481 10965 7515 10999
rect 8217 10965 8251 10999
rect 2513 10761 2547 10795
rect 3249 10761 3283 10795
rect 11529 10761 11563 10795
rect 13185 10761 13219 10795
rect 4414 10693 4448 10727
rect 12050 10693 12084 10727
rect 2605 10625 2639 10659
rect 3341 10625 3375 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 6561 10625 6595 10659
rect 6653 10625 6687 10659
rect 7021 10625 7055 10659
rect 7481 10625 7515 10659
rect 8309 10625 8343 10659
rect 9045 10625 9079 10659
rect 11713 10625 11747 10659
rect 13277 10625 13311 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 1961 10557 1995 10591
rect 2789 10557 2823 10591
rect 4169 10557 4203 10591
rect 6837 10557 6871 10591
rect 8125 10557 8159 10591
rect 8493 10557 8527 10591
rect 9229 10557 9263 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 11805 10557 11839 10591
rect 5549 10489 5583 10523
rect 3433 10421 3467 10455
rect 5733 10421 5767 10455
rect 6101 10421 6135 10455
rect 7573 10421 7607 10455
rect 8953 10421 8987 10455
rect 9689 10421 9723 10455
rect 10517 10421 10551 10455
rect 10977 10421 11011 10455
rect 13461 10421 13495 10455
rect 2513 10217 2547 10251
rect 5273 10217 5307 10251
rect 8401 10217 8435 10251
rect 9045 10217 9079 10251
rect 10149 10217 10183 10251
rect 10793 10217 10827 10251
rect 12173 10217 12207 10251
rect 13093 10217 13127 10251
rect 13461 10217 13495 10251
rect 2605 10149 2639 10183
rect 6745 10149 6779 10183
rect 10517 10149 10551 10183
rect 12081 10149 12115 10183
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 6285 10081 6319 10115
rect 11161 10081 11195 10115
rect 11529 10081 11563 10115
rect 2329 10013 2363 10047
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 5089 10013 5123 10047
rect 6101 10013 6135 10047
rect 6837 10013 6871 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 10241 10013 10275 10047
rect 10333 10013 10367 10047
rect 10609 10013 10643 10047
rect 11897 10013 11931 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13645 10013 13679 10047
rect 13829 10013 13863 10047
rect 14473 10013 14507 10047
rect 1501 9945 1535 9979
rect 1685 9945 1719 9979
rect 6009 9945 6043 9979
rect 7104 9945 7138 9979
rect 11253 9945 11287 9979
rect 2973 9877 3007 9911
rect 8217 9877 8251 9911
rect 14289 9877 14323 9911
rect 5917 9673 5951 9707
rect 7021 9673 7055 9707
rect 12357 9673 12391 9707
rect 8217 9605 8251 9639
rect 13277 9605 13311 9639
rect 1409 9537 1443 9571
rect 1869 9537 1903 9571
rect 3902 9537 3936 9571
rect 4445 9537 4479 9571
rect 5733 9537 5767 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 8861 9537 8895 9571
rect 9781 9537 9815 9571
rect 10048 9537 10082 9571
rect 12265 9537 12299 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 14197 9537 14231 9571
rect 14289 9537 14323 9571
rect 1777 9469 1811 9503
rect 2421 9469 2455 9503
rect 2605 9469 2639 9503
rect 4169 9469 4203 9503
rect 7573 9469 7607 9503
rect 9505 9469 9539 9503
rect 9689 9469 9723 9503
rect 12081 9469 12115 9503
rect 13737 9469 13771 9503
rect 13921 9469 13955 9503
rect 14381 9469 14415 9503
rect 2789 9401 2823 9435
rect 7297 9401 7331 9435
rect 11161 9401 11195 9435
rect 13001 9401 13035 9435
rect 14013 9401 14047 9435
rect 1593 9333 1627 9367
rect 2237 9333 2271 9367
rect 4629 9333 4663 9367
rect 8309 9333 8343 9367
rect 9321 9333 9355 9367
rect 11529 9333 11563 9367
rect 12725 9333 12759 9367
rect 2329 9129 2363 9163
rect 2881 9129 2915 9163
rect 8309 9129 8343 9163
rect 8493 9129 8527 9163
rect 9413 9129 9447 9163
rect 13093 9129 13127 9163
rect 13461 9129 13495 9163
rect 3985 9061 4019 9095
rect 4261 9061 4295 9095
rect 5549 9061 5583 9095
rect 13001 9061 13035 9095
rect 2145 8993 2179 9027
rect 4537 8993 4571 9027
rect 5825 8993 5859 9027
rect 1961 8925 1995 8959
rect 2973 8925 3007 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4353 8925 4387 8959
rect 5273 8925 5307 8959
rect 5365 8925 5399 8959
rect 5641 8925 5675 8959
rect 6561 8925 6595 8959
rect 6929 8925 6963 8959
rect 8677 8925 8711 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 11630 8925 11664 8959
rect 11897 8925 11931 8959
rect 12357 8925 12391 8959
rect 12541 8925 12575 8959
rect 13277 8925 13311 8959
rect 13369 8925 13403 8959
rect 13645 8925 13679 8959
rect 14289 8925 14323 8959
rect 1501 8857 1535 8891
rect 7196 8857 7230 8891
rect 9689 8857 9723 8891
rect 13737 8857 13771 8891
rect 1593 8789 1627 8823
rect 4997 8789 5031 8823
rect 5181 8789 5215 8823
rect 6285 8789 6319 8823
rect 6469 8789 6503 8823
rect 9045 8789 9079 8823
rect 10517 8789 10551 8823
rect 14105 8789 14139 8823
rect 1961 8585 1995 8619
rect 3801 8585 3835 8619
rect 4537 8585 4571 8619
rect 5457 8585 5491 8619
rect 6193 8585 6227 8619
rect 8033 8585 8067 8619
rect 1593 8517 1627 8551
rect 9781 8517 9815 8551
rect 10517 8517 10551 8551
rect 10609 8517 10643 8551
rect 1501 8449 1535 8483
rect 1777 8449 1811 8483
rect 2053 8449 2087 8483
rect 2145 8449 2179 8483
rect 2513 8449 2547 8483
rect 3709 8449 3743 8483
rect 4997 8449 5031 8483
rect 5273 8449 5307 8483
rect 5733 8449 5767 8483
rect 6561 8447 6595 8481
rect 6837 8449 6871 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8392 8449 8426 8483
rect 14105 8449 14139 8483
rect 2329 8381 2363 8415
rect 3525 8381 3559 8415
rect 4353 8381 4387 8415
rect 5181 8381 5215 8415
rect 5549 8381 5583 8415
rect 7021 8381 7055 8415
rect 7665 8381 7699 8415
rect 9689 8381 9723 8415
rect 10793 8381 10827 8415
rect 12081 8381 12115 8415
rect 12265 8381 12299 8415
rect 2973 8313 3007 8347
rect 3341 8313 3375 8347
rect 6653 8313 6687 8347
rect 7205 8313 7239 8347
rect 9505 8313 9539 8347
rect 10241 8313 10275 8347
rect 14197 8313 14231 8347
rect 11621 8245 11655 8279
rect 1593 8041 1627 8075
rect 3985 8041 4019 8075
rect 8493 8041 8527 8075
rect 9873 8041 9907 8075
rect 10241 8041 10275 8075
rect 11621 8041 11655 8075
rect 4353 7973 4387 8007
rect 9689 7973 9723 8007
rect 10333 7973 10367 8007
rect 11345 7973 11379 8007
rect 5733 7905 5767 7939
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 9045 7905 9079 7939
rect 9229 7905 9263 7939
rect 1777 7837 1811 7871
rect 2145 7837 2179 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 5917 7837 5951 7871
rect 6561 7837 6595 7871
rect 7665 7837 7699 7871
rect 8677 7837 8711 7871
rect 9957 7839 9991 7873
rect 10081 7837 10115 7871
rect 10517 7837 10551 7871
rect 11161 7837 11195 7871
rect 11437 7837 11471 7871
rect 2412 7769 2446 7803
rect 4445 7769 4479 7803
rect 4997 7769 5031 7803
rect 5089 7769 5123 7803
rect 5273 7769 5307 7803
rect 7389 7769 7423 7803
rect 2053 7701 2087 7735
rect 3525 7701 3559 7735
rect 6009 7701 6043 7735
rect 7481 7701 7515 7735
rect 2513 7497 2547 7531
rect 4721 7497 4755 7531
rect 9321 7497 9355 7531
rect 4353 7429 4387 7463
rect 7849 7429 7883 7463
rect 1593 7361 1627 7395
rect 4629 7361 4663 7395
rect 5181 7361 5215 7395
rect 7113 7361 7147 7395
rect 14473 7361 14507 7395
rect 1961 7293 1995 7327
rect 6929 7293 6963 7327
rect 7297 7293 7331 7327
rect 1777 7157 1811 7191
rect 3065 7157 3099 7191
rect 4997 7157 5031 7191
rect 6377 7157 6411 7191
rect 7481 7157 7515 7191
rect 14289 7157 14323 7191
rect 1409 6953 1443 6987
rect 4629 6953 4663 6987
rect 7021 6953 7055 6987
rect 2789 6817 2823 6851
rect 5457 6817 5491 6851
rect 8769 6817 8803 6851
rect 9689 6817 9723 6851
rect 2533 6749 2567 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 3525 6749 3559 6783
rect 4813 6749 4847 6783
rect 5724 6749 5758 6783
rect 6929 6749 6963 6783
rect 9781 6749 9815 6783
rect 3893 6681 3927 6715
rect 3985 6681 4019 6715
rect 4537 6681 4571 6715
rect 8502 6681 8536 6715
rect 9045 6681 9079 6715
rect 9137 6681 9171 6715
rect 6837 6613 6871 6647
rect 7389 6613 7423 6647
rect 9965 6613 9999 6647
rect 1777 6409 1811 6443
rect 2053 6409 2087 6443
rect 8493 6409 8527 6443
rect 10425 6409 10459 6443
rect 10977 6409 11011 6443
rect 11989 6409 12023 6443
rect 9413 6341 9447 6375
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7196 6273 7230 6307
rect 10241 6273 10275 6307
rect 10333 6273 10367 6307
rect 10885 6273 10919 6307
rect 12081 6273 12115 6307
rect 14473 6273 14507 6307
rect 9045 6205 9079 6239
rect 9321 6205 9355 6239
rect 10609 6205 10643 6239
rect 2697 6137 2731 6171
rect 6561 6137 6595 6171
rect 8309 6137 8343 6171
rect 9873 6137 9907 6171
rect 10057 6137 10091 6171
rect 14289 6137 14323 6171
rect 2513 6069 2547 6103
rect 2881 6069 2915 6103
rect 6745 6069 6779 6103
rect 1593 5865 1627 5899
rect 7665 5865 7699 5899
rect 8769 5865 8803 5899
rect 9229 5865 9263 5899
rect 6837 5797 6871 5831
rect 7941 5797 7975 5831
rect 9413 5729 9447 5763
rect 9597 5729 9631 5763
rect 1409 5661 1443 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 7021 5661 7055 5695
rect 7757 5661 7791 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 10057 5661 10091 5695
rect 12357 5661 12391 5695
rect 6561 5525 6595 5559
rect 10241 5525 10275 5559
rect 12173 5525 12207 5559
rect 7113 5321 7147 5355
rect 8217 5321 8251 5355
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 7205 5185 7239 5219
rect 7389 5185 7423 5219
rect 8953 5185 8987 5219
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 8677 5117 8711 5151
rect 8861 5117 8895 5151
rect 5917 5049 5951 5083
rect 6193 5049 6227 5083
rect 7573 5049 7607 5083
rect 9045 5049 9079 5083
rect 7021 4777 7055 4811
rect 8125 4777 8159 4811
rect 8677 4777 8711 4811
rect 14381 4777 14415 4811
rect 7389 4709 7423 4743
rect 7665 4641 7699 4675
rect 1409 4573 1443 4607
rect 7113 4573 7147 4607
rect 7205 4573 7239 4607
rect 7481 4573 7515 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 8585 4575 8619 4609
rect 14197 4573 14231 4607
rect 1593 4437 1627 4471
rect 8953 4097 8987 4131
rect 9137 3893 9171 3927
rect 5273 3689 5307 3723
rect 14289 3689 14323 3723
rect 1593 3621 1627 3655
rect 1409 3485 1443 3519
rect 5365 3485 5399 3519
rect 14473 3485 14507 3519
rect 13645 3077 13679 3111
rect 13921 3077 13955 3111
rect 1777 3009 1811 3043
rect 2053 3009 2087 3043
rect 2145 3009 2179 3043
rect 4077 3009 4111 3043
rect 5273 3009 5307 3043
rect 6745 3009 6779 3043
rect 8309 3009 8343 3043
rect 9597 3009 9631 3043
rect 10517 3009 10551 3043
rect 11897 3009 11931 3043
rect 12449 3009 12483 3043
rect 1501 2805 1535 2839
rect 4169 2805 4203 2839
rect 5457 2805 5491 2839
rect 6561 2805 6595 2839
rect 8217 2805 8251 2839
rect 9505 2805 9539 2839
rect 10609 2805 10643 2839
rect 12081 2805 12115 2839
rect 12633 2805 12667 2839
rect 13553 2805 13587 2839
rect 14013 2805 14047 2839
rect 14289 2601 14323 2635
rect 2605 2397 2639 2431
rect 3433 2397 3467 2431
rect 4261 2397 4295 2431
rect 4813 2397 4847 2431
rect 5641 2397 5675 2431
rect 6745 2397 6779 2431
rect 8401 2397 8435 2431
rect 9045 2397 9079 2431
rect 9781 2397 9815 2431
rect 10609 2397 10643 2431
rect 11621 2397 11655 2431
rect 12265 2397 12299 2431
rect 13093 2397 13127 2431
rect 14473 2397 14507 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 2237 2329 2271 2363
rect 3065 2329 3099 2363
rect 3893 2329 3927 2363
rect 6377 2329 6411 2363
rect 7205 2329 7239 2363
rect 7573 2329 7607 2363
rect 4905 2261 4939 2295
rect 5733 2261 5767 2295
rect 8125 2261 8159 2295
rect 9137 2261 9171 2295
rect 9873 2261 9907 2295
rect 10701 2261 10735 2295
rect 11713 2261 11747 2295
rect 12541 2261 12575 2295
rect 13185 2261 13219 2295
<< metal1 >>
rect 7650 17756 7656 17808
rect 7708 17796 7714 17808
rect 8294 17796 8300 17808
rect 7708 17768 8300 17796
rect 7708 17756 7714 17768
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 4614 17592 4620 17604
rect 3108 17564 4620 17592
rect 3108 17552 3114 17564
rect 4614 17552 4620 17564
rect 4672 17552 4678 17604
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 6638 17524 6644 17536
rect 3292 17496 6644 17524
rect 3292 17484 3298 17496
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 934 17280 940 17332
rect 992 17280 998 17332
rect 2406 17280 2412 17332
rect 2464 17280 2470 17332
rect 3142 17320 3148 17332
rect 2516 17292 3148 17320
rect 952 17184 980 17280
rect 2424 17252 2452 17280
rect 1780 17224 2452 17252
rect 1780 17193 1808 17224
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 952 17156 1501 17184
rect 1489 17153 1501 17156
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17184 2099 17187
rect 2516 17184 2544 17292
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 5350 17320 5356 17332
rect 3252 17292 5356 17320
rect 3050 17252 3056 17264
rect 2608 17224 3056 17252
rect 2608 17193 2636 17224
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 2087 17156 2544 17184
rect 2593 17187 2651 17193
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 2593 17153 2605 17187
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17184 2927 17187
rect 3252 17184 3280 17292
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 6086 17320 6092 17332
rect 5460 17292 6092 17320
rect 5460 17252 5488 17292
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6549 17323 6607 17329
rect 6549 17289 6561 17323
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17289 7527 17323
rect 7469 17283 7527 17289
rect 4816 17224 5488 17252
rect 2915 17156 3280 17184
rect 3329 17187 3387 17193
rect 2915 17153 2927 17156
rect 2869 17147 2927 17153
rect 3329 17153 3341 17187
rect 3375 17184 3387 17187
rect 3605 17187 3663 17193
rect 3375 17156 3464 17184
rect 3375 17153 3387 17156
rect 3329 17147 3387 17153
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17085 2559 17119
rect 2501 17079 2559 17085
rect 2516 17048 2544 17079
rect 3234 17076 3240 17128
rect 3292 17076 3298 17128
rect 3436 17057 3464 17156
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 4816 17184 4844 17224
rect 3651 17156 4844 17184
rect 5445 17187 5503 17193
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5718 17184 5724 17196
rect 5491 17156 5724 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6564 17184 6592 17283
rect 6641 17187 6699 17193
rect 6641 17184 6653 17187
rect 6564 17156 6653 17184
rect 6365 17147 6423 17153
rect 6641 17153 6653 17156
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 7484 17184 7512 17283
rect 7650 17280 7656 17332
rect 7708 17280 7714 17332
rect 7837 17323 7895 17329
rect 7837 17289 7849 17323
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 7668 17193 7696 17280
rect 7852 17252 7880 17283
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 9088 17292 9321 17320
rect 9088 17280 9094 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9824 17292 9965 17320
rect 9824 17280 9830 17292
rect 9953 17289 9965 17292
rect 9999 17289 10011 17323
rect 9953 17283 10011 17289
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10560 17292 10701 17320
rect 10560 17280 10566 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11204 17292 11621 17320
rect 11204 17280 11210 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12253 17323 12311 17329
rect 12253 17320 12265 17323
rect 12032 17292 12265 17320
rect 12032 17280 12038 17292
rect 12253 17289 12265 17292
rect 12299 17289 12311 17323
rect 12253 17283 12311 17289
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12768 17292 13001 17320
rect 12768 17280 12774 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13504 17292 13829 17320
rect 13504 17280 13510 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 10229 17255 10287 17261
rect 7852 17224 8248 17252
rect 7423 17156 7512 17184
rect 7653 17187 7711 17193
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7653 17153 7665 17187
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 3421 17051 3479 17057
rect 2516 17020 3372 17048
rect 1670 16940 1676 16992
rect 1728 16940 1734 16992
rect 1946 16940 1952 16992
rect 2004 16940 2010 16992
rect 2222 16940 2228 16992
rect 2280 16940 2286 16992
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 2958 16980 2964 16992
rect 2823 16952 2964 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16980 3111 16983
rect 3234 16980 3240 16992
rect 3099 16952 3240 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3344 16980 3372 17020
rect 3421 17017 3433 17051
rect 3467 17017 3479 17051
rect 3421 17011 3479 17017
rect 3896 16980 3924 17079
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 6196 17116 6224 17147
rect 4709 17079 4767 17085
rect 5644 17088 6224 17116
rect 6380 17116 6408 17147
rect 6822 17116 6828 17128
rect 6380 17088 6828 17116
rect 4724 16992 4752 17079
rect 5644 17057 5672 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6932 17116 6960 17147
rect 7750 17144 7756 17196
rect 7808 17144 7814 17196
rect 8220 17193 8248 17224
rect 10229 17221 10241 17255
rect 10275 17252 10287 17255
rect 11698 17252 11704 17264
rect 10275 17224 11704 17252
rect 10275 17221 10287 17224
rect 10229 17215 10287 17221
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 9214 17144 9220 17196
rect 9272 17144 9278 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 7558 17116 7564 17128
rect 6932 17088 7564 17116
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 10980 17116 11008 17147
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12676 17156 12909 17184
rect 12676 17144 12682 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13320 17156 13553 17184
rect 13320 17144 13326 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13780 17156 14105 17184
rect 13780 17144 13786 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 12066 17116 12072 17128
rect 10980 17088 12072 17116
rect 8021 17079 8079 17085
rect 5629 17051 5687 17057
rect 5629 17017 5641 17051
rect 5675 17017 5687 17051
rect 5629 17011 5687 17017
rect 7285 17051 7343 17057
rect 7285 17017 7297 17051
rect 7331 17048 7343 17051
rect 8036 17048 8064 17079
rect 12066 17076 12072 17088
rect 12124 17076 12130 17128
rect 7331 17020 8064 17048
rect 7331 17017 7343 17020
rect 7285 17011 7343 17017
rect 3344 16952 3924 16980
rect 4522 16940 4528 16992
rect 4580 16940 4586 16992
rect 4706 16940 4712 16992
rect 4764 16940 4770 16992
rect 5258 16940 5264 16992
rect 5316 16940 5322 16992
rect 5810 16940 5816 16992
rect 5868 16940 5874 16992
rect 5994 16940 6000 16992
rect 6052 16940 6058 16992
rect 6730 16940 6736 16992
rect 6788 16940 6794 16992
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 8386 16980 8392 16992
rect 7147 16952 8392 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 14185 16983 14243 16989
rect 14185 16980 14197 16983
rect 11112 16952 14197 16980
rect 11112 16940 11118 16952
rect 14185 16949 14197 16952
rect 14231 16949 14243 16983
rect 14185 16943 14243 16949
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 1670 16736 1676 16788
rect 1728 16736 1734 16788
rect 3050 16736 3056 16788
rect 3108 16736 3114 16788
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 4062 16776 4068 16788
rect 3375 16748 4068 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4522 16736 4528 16788
rect 4580 16736 4586 16788
rect 8665 16779 8723 16785
rect 6564 16748 7788 16776
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 1688 16581 1716 16736
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16677 2835 16711
rect 2777 16671 2835 16677
rect 1872 16612 2084 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 1762 16532 1768 16584
rect 1820 16572 1826 16584
rect 1872 16572 1900 16612
rect 1820 16544 1900 16572
rect 1949 16575 2007 16581
rect 1820 16532 1826 16544
rect 1949 16541 1961 16575
rect 1995 16541 2007 16575
rect 2056 16572 2084 16612
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 2056 16544 2237 16572
rect 1949 16535 2007 16541
rect 2225 16541 2237 16544
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16541 2651 16575
rect 2792 16572 2820 16671
rect 3068 16640 3096 16736
rect 3068 16612 3464 16640
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 2792 16544 2881 16572
rect 2593 16535 2651 16541
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 1964 16504 1992 16535
rect 1596 16476 1992 16504
rect 2608 16504 2636 16535
rect 3142 16532 3148 16584
rect 3200 16532 3206 16584
rect 3436 16581 3464 16612
rect 3878 16600 3884 16652
rect 3936 16600 3942 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4154 16640 4160 16652
rect 4111 16612 4160 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4540 16640 4568 16736
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 4540 16612 5641 16640
rect 5629 16609 5641 16612
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 5776 16612 6377 16640
rect 5776 16600 5782 16612
rect 6365 16609 6377 16612
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 3568 16544 4752 16572
rect 3568 16532 3574 16544
rect 3786 16504 3792 16516
rect 2608 16476 3792 16504
rect 1596 16445 1624 16476
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 4724 16504 4752 16544
rect 4798 16532 4804 16584
rect 4856 16532 4862 16584
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 6564 16516 6592 16748
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 7331 16680 7512 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7385 16575 7443 16581
rect 7385 16541 7397 16575
rect 7431 16572 7443 16575
rect 7484 16572 7512 16680
rect 7431 16544 7512 16572
rect 7431 16541 7443 16544
rect 7385 16535 7443 16541
rect 4890 16504 4896 16516
rect 4724 16476 4896 16504
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 5721 16507 5779 16513
rect 5721 16473 5733 16507
rect 5767 16504 5779 16507
rect 5994 16504 6000 16516
rect 5767 16476 6000 16504
rect 5767 16473 5779 16476
rect 5721 16467 5779 16473
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 6273 16507 6331 16513
rect 6273 16473 6285 16507
rect 6319 16504 6331 16507
rect 6546 16504 6552 16516
rect 6319 16476 6552 16504
rect 6319 16473 6331 16476
rect 6273 16467 6331 16473
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 7116 16504 7144 16535
rect 7650 16532 7656 16584
rect 7708 16532 7714 16584
rect 7760 16572 7788 16748
rect 8665 16745 8677 16779
rect 8711 16776 8723 16779
rect 9214 16776 9220 16788
rect 8711 16748 9220 16776
rect 8711 16745 8723 16748
rect 8665 16739 8723 16745
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 11698 16736 11704 16788
rect 11756 16736 11762 16788
rect 11882 16736 11888 16788
rect 11940 16736 11946 16788
rect 12618 16736 12624 16788
rect 12676 16736 12682 16788
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 13262 16776 13268 16788
rect 12943 16748 13268 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 13357 16779 13415 16785
rect 13357 16745 13369 16779
rect 13403 16776 13415 16779
rect 13722 16776 13728 16788
rect 13403 16748 13728 16776
rect 13403 16745 13415 16748
rect 13357 16739 13415 16745
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 14182 16776 14188 16788
rect 13863 16748 14188 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 12526 16708 12532 16720
rect 12360 16680 12532 16708
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9723 16612 10149 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10137 16609 10149 16612
rect 10183 16640 10195 16643
rect 10183 16612 11652 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 7760 16544 8585 16572
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 10594 16532 10600 16584
rect 10652 16532 10658 16584
rect 10778 16532 10784 16584
rect 10836 16532 10842 16584
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11624 16581 11652 16612
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 11204 16544 11345 16572
rect 11204 16532 11210 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12360 16581 12388 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 13170 16708 13176 16720
rect 13096 16680 13176 16708
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 12032 16544 12081 16572
rect 12032 16532 12038 16544
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 7668 16504 7696 16532
rect 7116 16476 7696 16504
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8536 16476 9045 16504
rect 8536 16464 8542 16476
rect 9033 16473 9045 16476
rect 9079 16473 9091 16507
rect 9033 16467 9091 16473
rect 9122 16464 9128 16516
rect 9180 16464 9186 16516
rect 9861 16507 9919 16513
rect 9861 16504 9873 16507
rect 9784 16476 9873 16504
rect 9784 16448 9812 16476
rect 9861 16473 9873 16476
rect 9907 16473 9919 16507
rect 9861 16467 9919 16473
rect 9950 16464 9956 16516
rect 10008 16464 10014 16516
rect 10686 16464 10692 16516
rect 10744 16504 10750 16516
rect 11425 16507 11483 16513
rect 11425 16504 11437 16507
rect 10744 16476 11437 16504
rect 10744 16464 10750 16476
rect 11425 16473 11437 16476
rect 11471 16473 11483 16507
rect 12452 16504 12480 16535
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 12584 16544 12725 16572
rect 12584 16532 12590 16544
rect 12713 16541 12725 16544
rect 12759 16541 12771 16575
rect 13096 16572 13124 16680
rect 13170 16668 13176 16680
rect 13228 16668 13234 16720
rect 13173 16575 13231 16581
rect 13173 16572 13185 16575
rect 13096 16544 13185 16572
rect 12713 16535 12771 16541
rect 13173 16541 13185 16544
rect 13219 16541 13231 16575
rect 13173 16535 13231 16541
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13688 16544 14105 16572
rect 13688 16532 13694 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 13262 16504 13268 16516
rect 12452 16476 13268 16504
rect 11425 16467 11483 16473
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 13538 16464 13544 16516
rect 13596 16464 13602 16516
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 1762 16396 1768 16448
rect 1820 16396 1826 16448
rect 2038 16396 2044 16448
rect 2096 16396 2102 16448
rect 2409 16439 2467 16445
rect 2409 16405 2421 16439
rect 2455 16436 2467 16439
rect 2866 16436 2872 16448
rect 2455 16408 2872 16436
rect 2455 16405 2467 16408
rect 2409 16399 2467 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 2961 16439 3019 16445
rect 2961 16405 2973 16439
rect 3007 16436 3019 16439
rect 3418 16436 3424 16448
rect 3007 16408 3424 16436
rect 3007 16405 3019 16408
rect 2961 16399 3019 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 3513 16439 3571 16445
rect 3513 16405 3525 16439
rect 3559 16436 3571 16439
rect 5074 16436 5080 16448
rect 3559 16408 5080 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5442 16396 5448 16448
rect 5500 16396 5506 16448
rect 7006 16396 7012 16448
rect 7064 16396 7070 16448
rect 7558 16396 7564 16448
rect 7616 16396 7622 16448
rect 8294 16396 8300 16448
rect 8352 16396 8358 16448
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 11241 16439 11299 16445
rect 11241 16436 11253 16439
rect 9824 16408 11253 16436
rect 9824 16396 9830 16408
rect 11241 16405 11253 16408
rect 11287 16405 11299 16439
rect 11241 16399 11299 16405
rect 12250 16396 12256 16448
rect 12308 16396 12314 16448
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 14185 16439 14243 16445
rect 14185 16436 14197 16439
rect 13780 16408 14197 16436
rect 13780 16396 13786 16408
rect 14185 16405 14197 16408
rect 14231 16405 14243 16439
rect 14185 16399 14243 16405
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 1762 16192 1768 16244
rect 1820 16192 1826 16244
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 3418 16232 3424 16244
rect 2915 16204 3424 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 4433 16235 4491 16241
rect 4433 16201 4445 16235
rect 4479 16232 4491 16235
rect 4982 16232 4988 16244
rect 4479 16204 4988 16232
rect 4479 16201 4491 16204
rect 4433 16195 4491 16201
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5776 16204 6009 16232
rect 5776 16192 5782 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 8294 16192 8300 16244
rect 8352 16192 8358 16244
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16201 9091 16235
rect 9033 16195 9091 16201
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9950 16232 9956 16244
rect 9447 16204 9956 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 1780 16164 1808 16192
rect 4004 16167 4062 16173
rect 1780 16136 2176 16164
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1811 16068 1900 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1872 15969 1900 16068
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2148 16105 2176 16136
rect 4004 16133 4016 16167
rect 4050 16164 4062 16167
rect 4246 16164 4252 16176
rect 4050 16136 4252 16164
rect 4050 16133 4062 16136
rect 4004 16127 4062 16133
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 4706 16164 4712 16176
rect 4417 16136 4712 16164
rect 4417 16105 4445 16136
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 4884 16167 4942 16173
rect 4884 16133 4896 16167
rect 4930 16164 4942 16167
rect 5258 16164 5264 16176
rect 4930 16136 5264 16164
rect 4930 16133 4942 16136
rect 4884 16127 4942 16133
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 5868 16136 6561 16164
rect 5868 16124 5874 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 8312 16164 8340 16192
rect 8398 16167 8456 16173
rect 8398 16164 8410 16167
rect 8312 16136 8410 16164
rect 6549 16127 6607 16133
rect 8398 16133 8410 16136
rect 8444 16133 8456 16167
rect 8398 16127 8456 16133
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 4365 16099 4445 16105
rect 4365 16065 4377 16099
rect 4411 16068 4445 16099
rect 4411 16065 4423 16068
rect 4365 16059 4423 16065
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 8846 16096 8852 16108
rect 5500 16068 6040 16096
rect 5500 16056 5506 16068
rect 2314 15988 2320 16040
rect 2372 15988 2378 16040
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 16028 4307 16031
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4295 16000 4629 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 6012 16028 6040 16068
rect 7300 16068 8852 16096
rect 6457 16031 6515 16037
rect 6457 16028 6469 16031
rect 6012 16000 6469 16028
rect 4617 15991 4675 15997
rect 6457 15997 6469 16000
rect 6503 15997 6515 16031
rect 6457 15991 6515 15997
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15929 1915 15963
rect 1857 15923 1915 15929
rect 2777 15963 2835 15969
rect 2777 15929 2789 15963
rect 2823 15960 2835 15963
rect 2823 15932 3372 15960
rect 2823 15929 2835 15932
rect 2777 15923 2835 15929
rect 1670 15852 1676 15904
rect 1728 15852 1734 15904
rect 3344 15892 3372 15932
rect 3510 15892 3516 15904
rect 3344 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 4632 15892 4660 15991
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 6604 16000 6745 16028
rect 6604 15988 6610 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 7300 15969 7328 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9048 16096 9076 16195
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10686 16192 10692 16244
rect 10744 16192 10750 16244
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10836 16204 10885 16232
rect 10836 16192 10842 16204
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11701 16235 11759 16241
rect 11701 16201 11713 16235
rect 11747 16232 11759 16235
rect 12158 16232 12164 16244
rect 11747 16204 12164 16232
rect 11747 16201 11759 16204
rect 11701 16195 11759 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12250 16192 12256 16244
rect 12308 16232 12314 16244
rect 12308 16204 12434 16232
rect 12308 16192 12314 16204
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 9766 16164 9772 16176
rect 9723 16136 9772 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 9766 16124 9772 16136
rect 9824 16124 9830 16176
rect 10704 16164 10732 16192
rect 10152 16136 10732 16164
rect 12406 16164 12434 16204
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13596 16204 13645 16232
rect 13596 16192 13602 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 13633 16195 13691 16201
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 15010 16232 15016 16244
rect 14415 16204 15016 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 12406 16136 14105 16164
rect 10152 16105 10180 16136
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 14093 16127 14151 16133
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 9048 16068 9229 16096
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9030 16028 9036 16040
rect 8711 16000 9036 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 10336 16028 10364 16059
rect 10410 16056 10416 16108
rect 10468 16056 10474 16108
rect 10686 16056 10692 16108
rect 10744 16056 10750 16108
rect 11609 16099 11667 16105
rect 11609 16065 11621 16099
rect 11655 16096 11667 16099
rect 11655 16068 11744 16096
rect 11655 16065 11667 16068
rect 11609 16059 11667 16065
rect 11054 16028 11060 16040
rect 10336 16000 11060 16028
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11146 15988 11152 16040
rect 11204 15988 11210 16040
rect 7285 15963 7343 15969
rect 7285 15929 7297 15963
rect 7331 15929 7343 15963
rect 7285 15923 7343 15929
rect 11716 15904 11744 16068
rect 12342 16056 12348 16108
rect 12400 16096 12406 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 12400 16068 13277 16096
rect 12400 16056 12406 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13412 16068 13553 16096
rect 13412 16056 13418 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 12802 15988 12808 16040
rect 12860 15988 12866 16040
rect 6454 15892 6460 15904
rect 4632 15864 6460 15892
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 10597 15895 10655 15901
rect 10597 15861 10609 15895
rect 10643 15892 10655 15895
rect 11054 15892 11060 15904
rect 10643 15864 11060 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11698 15852 11704 15904
rect 11756 15852 11762 15904
rect 13446 15852 13452 15904
rect 13504 15852 13510 15904
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2372 15660 2697 15688
rect 2372 15648 2378 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 4154 15648 4160 15700
rect 4212 15648 4218 15700
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 5905 15691 5963 15697
rect 5905 15688 5917 15691
rect 5500 15660 5917 15688
rect 5500 15648 5506 15660
rect 5905 15657 5917 15660
rect 5951 15657 5963 15691
rect 5905 15651 5963 15657
rect 6012 15660 7236 15688
rect 3160 15620 3188 15648
rect 4617 15623 4675 15629
rect 4617 15620 4629 15623
rect 3160 15592 4629 15620
rect 4617 15589 4629 15592
rect 4663 15589 4675 15623
rect 4617 15583 4675 15589
rect 3418 15512 3424 15564
rect 3476 15512 3482 15564
rect 3510 15512 3516 15564
rect 3568 15552 3574 15564
rect 4816 15552 4844 15648
rect 5077 15623 5135 15629
rect 5077 15589 5089 15623
rect 5123 15589 5135 15623
rect 6012 15620 6040 15660
rect 5077 15583 5135 15589
rect 5552 15592 6040 15620
rect 7208 15620 7236 15660
rect 8478 15648 8484 15700
rect 8536 15648 8542 15700
rect 9122 15648 9128 15700
rect 9180 15688 9186 15700
rect 9769 15691 9827 15697
rect 9769 15688 9781 15691
rect 9180 15660 9781 15688
rect 9180 15648 9186 15660
rect 9769 15657 9781 15660
rect 9815 15657 9827 15691
rect 9769 15651 9827 15657
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10686 15688 10692 15700
rect 10183 15660 10692 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11146 15648 11152 15700
rect 11204 15648 11210 15700
rect 12802 15648 12808 15700
rect 12860 15648 12866 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13354 15688 13360 15700
rect 13127 15660 13360 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13446 15648 13452 15700
rect 13504 15648 13510 15700
rect 7208 15592 10824 15620
rect 3568 15524 4844 15552
rect 3568 15512 3574 15524
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15453 2835 15487
rect 2777 15447 2835 15453
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 2958 15484 2964 15496
rect 2915 15456 2964 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 2792 15416 2820 15447
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3050 15444 3056 15496
rect 3108 15444 3114 15496
rect 3436 15484 3464 15512
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 3436 15456 4261 15484
rect 4249 15453 4261 15456
rect 4295 15484 4307 15487
rect 4706 15484 4712 15496
rect 4295 15456 4712 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4706 15444 4712 15456
rect 4764 15484 4770 15496
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4764 15456 4813 15484
rect 4764 15444 4770 15456
rect 4801 15453 4813 15456
rect 4847 15484 4859 15487
rect 4893 15487 4951 15493
rect 4893 15484 4905 15487
rect 4847 15456 4905 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 4893 15453 4905 15456
rect 4939 15453 4951 15487
rect 5092 15484 5120 15583
rect 5552 15564 5580 15592
rect 5534 15512 5540 15564
rect 5592 15512 5598 15564
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7616 15524 8033 15552
rect 7616 15512 7622 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8846 15512 8852 15564
rect 8904 15552 8910 15564
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8904 15524 8953 15552
rect 8904 15512 8910 15524
rect 8941 15521 8953 15524
rect 8987 15552 8999 15555
rect 10413 15555 10471 15561
rect 8987 15524 9720 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 5092 15456 5273 15484
rect 4893 15447 4951 15453
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5500 15456 5733 15484
rect 5500 15444 5506 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6540 15487 6598 15493
rect 6319 15456 6500 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6472 15428 6500 15456
rect 6540 15453 6552 15487
rect 6586 15484 6598 15487
rect 7006 15484 7012 15496
rect 6586 15456 7012 15484
rect 6586 15453 6598 15456
rect 6540 15447 6598 15453
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7524 15456 7849 15484
rect 7524 15444 7530 15456
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 9692 15493 9720 15524
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 10594 15552 10600 15564
rect 10459 15524 10600 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8444 15456 8585 15484
rect 8444 15444 8450 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 2792 15388 3372 15416
rect 3344 15360 3372 15388
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 4120 15388 5672 15416
rect 4120 15376 4126 15388
rect 3326 15308 3332 15360
rect 3384 15308 3390 15360
rect 5442 15308 5448 15360
rect 5500 15308 5506 15360
rect 5644 15348 5672 15388
rect 6454 15376 6460 15428
rect 6512 15376 6518 15428
rect 7098 15376 7104 15428
rect 7156 15416 7162 15428
rect 8665 15419 8723 15425
rect 8665 15416 8677 15419
rect 7156 15388 8677 15416
rect 7156 15376 7162 15388
rect 8665 15385 8677 15388
rect 8711 15385 8723 15419
rect 9968 15416 9996 15447
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10686 15444 10692 15496
rect 10744 15444 10750 15496
rect 10796 15484 10824 15592
rect 11164 15552 11192 15648
rect 12345 15623 12403 15629
rect 12345 15589 12357 15623
rect 12391 15589 12403 15623
rect 12345 15583 12403 15589
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11164 15524 11253 15552
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 12360 15552 12388 15583
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 11241 15515 11299 15521
rect 11348 15524 12020 15552
rect 12360 15524 12633 15552
rect 11348 15484 11376 15524
rect 10796 15456 11376 15484
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 11606 15484 11612 15496
rect 11471 15456 11612 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 8665 15379 8723 15385
rect 8772 15388 9996 15416
rect 6914 15348 6920 15360
rect 5644 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8772 15348 8800 15388
rect 7708 15320 8800 15348
rect 7708 15308 7714 15320
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9585 15351 9643 15357
rect 9585 15348 9597 15351
rect 9364 15320 9597 15348
rect 9364 15308 9370 15320
rect 9585 15317 9597 15320
rect 9631 15317 9643 15351
rect 9968 15348 9996 15388
rect 11149 15419 11207 15425
rect 11149 15385 11161 15419
rect 11195 15416 11207 15419
rect 11698 15416 11704 15428
rect 11195 15388 11704 15416
rect 11195 15385 11207 15388
rect 11149 15379 11207 15385
rect 11698 15376 11704 15388
rect 11756 15416 11762 15428
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11756 15388 11897 15416
rect 11756 15376 11762 15388
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11992 15416 12020 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 12158 15444 12164 15496
rect 12216 15444 12222 15496
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15484 12495 15487
rect 12820 15484 12848 15648
rect 13464 15552 13492 15648
rect 13464 15524 14136 15552
rect 14108 15493 14136 15524
rect 12483 15456 12848 15484
rect 14093 15487 14151 15493
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 13173 15419 13231 15425
rect 13173 15416 13185 15419
rect 11992 15388 13185 15416
rect 11885 15379 11943 15385
rect 13173 15385 13185 15388
rect 13219 15385 13231 15419
rect 13173 15379 13231 15385
rect 13722 15376 13728 15428
rect 13780 15376 13786 15428
rect 13814 15376 13820 15428
rect 13872 15376 13878 15428
rect 11238 15348 11244 15360
rect 9968 15320 11244 15348
rect 9585 15311 9643 15317
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3050 15144 3056 15156
rect 3007 15116 3056 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3234 15104 3240 15156
rect 3292 15144 3298 15156
rect 3292 15116 4292 15144
rect 3292 15104 3298 15116
rect 2222 15036 2228 15088
rect 2280 15076 2286 15088
rect 2280 15048 3464 15076
rect 2280 15036 2286 15048
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 3237 15011 3295 15017
rect 2823 14980 3096 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 3068 14881 3096 14980
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3326 15008 3332 15020
rect 3283 14980 3332 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3053 14875 3111 14881
rect 3053 14841 3065 14875
rect 3099 14841 3111 14875
rect 3053 14835 3111 14841
rect 3252 14804 3280 14971
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3436 15017 3464 15048
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 15008 3571 15011
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3559 14980 3709 15008
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 3697 14977 3709 14980
rect 3743 15008 3755 15011
rect 4264 15008 4292 15116
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 4396 15116 8033 15144
rect 4396 15104 4402 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10686 15144 10692 15156
rect 10459 15116 10692 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11606 15144 11612 15156
rect 11563 15116 11612 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12158 15144 12164 15156
rect 12023 15116 12164 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13412 15116 13461 15144
rect 13412 15104 13418 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14369 15147 14427 15153
rect 14369 15144 14381 15147
rect 13872 15116 14381 15144
rect 13872 15104 13878 15116
rect 14369 15113 14381 15116
rect 14415 15113 14427 15147
rect 14369 15107 14427 15113
rect 4798 15036 4804 15088
rect 4856 15076 4862 15088
rect 4856 15048 8708 15076
rect 4856 15036 4862 15048
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 3743 14980 4200 15008
rect 4264 14980 5181 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14909 3939 14943
rect 4172 14940 4200 14980
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 6546 14968 6552 15020
rect 6604 14968 6610 15020
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 8680 15017 8708 15048
rect 9416 15048 14228 15076
rect 9416 15017 9444 15048
rect 14200 15020 14228 15048
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 9401 15011 9459 15017
rect 8711 14980 9352 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 4172 14912 5212 14940
rect 3881 14903 3939 14909
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 3896 14872 3924 14903
rect 4798 14872 4804 14884
rect 3660 14844 3924 14872
rect 3988 14844 4804 14872
rect 3660 14832 3666 14844
rect 3988 14804 4016 14844
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 5184 14816 5212 14912
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 5994 14832 6000 14884
rect 6052 14872 6058 14884
rect 7024 14872 7052 14903
rect 6052 14844 7052 14872
rect 7929 14875 7987 14881
rect 6052 14832 6058 14844
rect 7929 14841 7941 14875
rect 7975 14872 7987 14875
rect 9232 14872 9260 14903
rect 7975 14844 9260 14872
rect 9324 14872 9352 14980
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10468 14980 10517 15008
rect 10468 14968 10474 14980
rect 10505 14977 10517 14980
rect 10551 15008 10563 15011
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 10551 14980 10609 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 10597 14977 10609 14980
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11112 14980 11713 15008
rect 11112 14968 11118 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 13354 15008 13360 15020
rect 11839 14980 13360 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 13354 14968 13360 14980
rect 13412 15008 13418 15020
rect 14093 15011 14151 15017
rect 14093 15008 14105 15011
rect 13412 14980 14105 15008
rect 13412 14968 13418 14980
rect 14093 14977 14105 14980
rect 14139 14977 14151 15011
rect 14093 14971 14151 14977
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11940 14912 12081 14940
rect 11940 14900 11946 14912
rect 12069 14909 12081 14912
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14940 13047 14943
rect 13538 14940 13544 14952
rect 13035 14912 13544 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 9324 14844 11376 14872
rect 7975 14841 7987 14844
rect 7929 14835 7987 14841
rect 3252 14776 4016 14804
rect 4154 14764 4160 14816
rect 4212 14764 4218 14816
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 5258 14764 5264 14816
rect 5316 14764 5322 14816
rect 6733 14807 6791 14813
rect 6733 14773 6745 14807
rect 6779 14804 6791 14807
rect 7190 14804 7196 14816
rect 6779 14776 7196 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7834 14804 7840 14816
rect 7515 14776 7840 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8754 14764 8760 14816
rect 8812 14764 8818 14816
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 9493 14807 9551 14813
rect 9493 14804 9505 14807
rect 9456 14776 9505 14804
rect 9456 14764 9462 14776
rect 9493 14773 9505 14776
rect 9539 14773 9551 14807
rect 9493 14767 9551 14773
rect 11238 14764 11244 14816
rect 11296 14764 11302 14816
rect 11348 14804 11376 14844
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 12820 14872 12848 14903
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 11756 14844 12848 14872
rect 11756 14832 11762 14844
rect 12434 14804 12440 14816
rect 11348 14776 12440 14804
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12710 14764 12716 14816
rect 12768 14764 12774 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13541 14807 13599 14813
rect 13541 14804 13553 14807
rect 12860 14776 13553 14804
rect 12860 14764 12866 14776
rect 13541 14773 13553 14776
rect 13587 14773 13599 14807
rect 13541 14767 13599 14773
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 4985 14603 5043 14609
rect 4985 14569 4997 14603
rect 5031 14600 5043 14603
rect 5031 14572 5580 14600
rect 5031 14569 5043 14572
rect 4985 14563 5043 14569
rect 3605 14535 3663 14541
rect 3605 14501 3617 14535
rect 3651 14532 3663 14535
rect 5077 14535 5135 14541
rect 3651 14504 4384 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 4356 14473 4384 14504
rect 5077 14501 5089 14535
rect 5123 14501 5135 14535
rect 5077 14495 5135 14501
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 3418 14356 3424 14408
rect 3476 14356 3482 14408
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14396 4859 14399
rect 5092 14396 5120 14495
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 5316 14504 5396 14532
rect 5316 14492 5322 14504
rect 5368 14473 5396 14504
rect 5552 14473 5580 14572
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5868 14572 6009 14600
rect 5868 14560 5874 14572
rect 5997 14569 6009 14572
rect 6043 14600 6055 14603
rect 6822 14600 6828 14612
rect 6043 14572 6828 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7190 14560 7196 14612
rect 7248 14560 7254 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 7800 14572 8309 14600
rect 7800 14560 7806 14572
rect 8297 14569 8309 14572
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 8754 14560 8760 14612
rect 8812 14560 8818 14612
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 13354 14560 13360 14612
rect 13412 14560 13418 14612
rect 13538 14560 13544 14612
rect 13596 14560 13602 14612
rect 14274 14560 14280 14612
rect 14332 14560 14338 14612
rect 5902 14492 5908 14544
rect 5960 14532 5966 14544
rect 5960 14504 7144 14532
rect 5960 14492 5966 14504
rect 7116 14476 7144 14504
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 4847 14368 5120 14396
rect 5184 14436 5365 14464
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 4540 14328 4568 14359
rect 5184 14328 5212 14436
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6595 14436 6929 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 7098 14424 7104 14476
rect 7156 14424 7162 14476
rect 7208 14464 7236 14560
rect 7377 14535 7435 14541
rect 7377 14501 7389 14535
rect 7423 14532 7435 14535
rect 8772 14532 8800 14560
rect 7423 14504 8800 14532
rect 7423 14501 7435 14504
rect 7377 14495 7435 14501
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7208 14436 7665 14464
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 7653 14427 7711 14433
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 5316 14368 6285 14396
rect 5316 14356 5322 14368
rect 6273 14365 6285 14368
rect 6319 14396 6331 14399
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6319 14368 6469 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7116 14396 7144 14424
rect 6779 14368 7144 14396
rect 7469 14399 7527 14405
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7760 14396 7788 14504
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8113 14467 8171 14473
rect 8113 14464 8125 14467
rect 7892 14436 8125 14464
rect 7892 14424 7898 14436
rect 8113 14433 8125 14436
rect 8159 14433 8171 14467
rect 8113 14427 8171 14433
rect 9030 14424 9036 14476
rect 9088 14424 9094 14476
rect 10042 14424 10048 14476
rect 10100 14424 10106 14476
rect 7515 14368 7788 14396
rect 8481 14399 8539 14405
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 8481 14365 8493 14399
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 4540 14300 5212 14328
rect 1578 14220 1584 14272
rect 1636 14220 1642 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4154 14260 4160 14272
rect 3927 14232 4160 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 6178 14220 6184 14272
rect 6236 14220 6242 14272
rect 6472 14260 6500 14359
rect 8496 14328 8524 14359
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 10060 14396 10088 14424
rect 8812 14368 10088 14396
rect 8812 14356 8818 14368
rect 11238 14356 11244 14408
rect 11296 14396 11302 14408
rect 11618 14399 11676 14405
rect 11618 14396 11630 14399
rect 11296 14368 11630 14396
rect 11296 14356 11302 14368
rect 11618 14365 11630 14368
rect 11664 14365 11676 14399
rect 11618 14359 11676 14365
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11848 14368 11897 14396
rect 11848 14356 11854 14368
rect 11885 14365 11897 14368
rect 11931 14396 11943 14399
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11931 14368 11989 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12244 14399 12302 14405
rect 12244 14365 12256 14399
rect 12290 14396 12302 14399
rect 12710 14396 12716 14408
rect 12290 14368 12716 14396
rect 12290 14365 12302 14368
rect 12244 14359 12302 14365
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 13372 14396 13400 14560
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13372 14368 13645 14396
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14550 14396 14556 14408
rect 14507 14368 14556 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 8846 14328 8852 14340
rect 8496 14300 8852 14328
rect 8496 14260 8524 14300
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 9300 14331 9358 14337
rect 9300 14297 9312 14331
rect 9346 14328 9358 14331
rect 9398 14328 9404 14340
rect 9346 14300 9404 14328
rect 9346 14297 9358 14300
rect 9300 14291 9358 14297
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 6472 14232 8524 14260
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 9858 14260 9864 14272
rect 8711 14232 9864 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14260 10563 14263
rect 11882 14260 11888 14272
rect 10551 14232 11888 14260
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 13630 14260 13636 14272
rect 12492 14232 13636 14260
rect 12492 14220 12498 14232
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14025 1731 14059
rect 1673 14019 1731 14025
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13920 1455 13923
rect 1688 13920 1716 14019
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 3418 14056 3424 14068
rect 3283 14028 3424 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3602 14016 3608 14068
rect 3660 14016 3666 14068
rect 4798 14016 4804 14068
rect 4856 14016 4862 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6089 14059 6147 14065
rect 6089 14056 6101 14059
rect 6052 14028 6101 14056
rect 6052 14016 6058 14028
rect 6089 14025 6101 14028
rect 6135 14025 6147 14059
rect 6089 14019 6147 14025
rect 6178 14016 6184 14068
rect 6236 14016 6242 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 6604 14028 7849 14056
rect 6604 14016 6610 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 8205 14059 8263 14065
rect 8205 14025 8217 14059
rect 8251 14056 8263 14059
rect 8754 14056 8760 14068
rect 8251 14028 8760 14056
rect 8251 14025 8263 14028
rect 8205 14019 8263 14025
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14025 10379 14059
rect 10321 14019 10379 14025
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 11054 14056 11060 14068
rect 10643 14028 11060 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 1964 13988 1992 14016
rect 1872 13960 2774 13988
rect 1872 13929 1900 13960
rect 1443 13892 1716 13920
rect 1857 13923 1915 13929
rect 1443 13889 1455 13892
rect 1397 13883 1455 13889
rect 1857 13889 1869 13923
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2038 13920 2044 13932
rect 1995 13892 2044 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2746 13920 2774 13960
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2746 13892 3065 13920
rect 3053 13889 3065 13892
rect 3099 13920 3111 13923
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 3099 13892 3341 13920
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3620 13920 3648 14016
rect 4433 13991 4491 13997
rect 4433 13988 4445 13991
rect 4080 13960 4445 13988
rect 4080 13929 4108 13960
rect 4433 13957 4445 13960
rect 4479 13957 4491 13991
rect 4433 13951 4491 13957
rect 3467 13892 3648 13920
rect 4065 13923 4123 13929
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4065 13883 4123 13889
rect 4172 13892 4353 13920
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 1596 13824 2145 13852
rect 1596 13793 1624 13824
rect 2133 13821 2145 13824
rect 2179 13821 2191 13855
rect 3344 13852 3372 13883
rect 4172 13852 4200 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 4816 13920 4844 14016
rect 6196 13988 6224 14016
rect 5368 13960 6224 13988
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4816 13892 4905 13920
rect 4341 13883 4399 13889
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5166 13880 5172 13932
rect 5224 13880 5230 13932
rect 5368 13929 5396 13960
rect 9306 13948 9312 14000
rect 9364 13997 9370 14000
rect 9364 13988 9376 13997
rect 9364 13960 9409 13988
rect 9364 13951 9376 13960
rect 9364 13948 9370 13951
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5902 13880 5908 13932
rect 5960 13880 5966 13932
rect 6005 13923 6063 13929
rect 6005 13889 6017 13923
rect 6051 13920 6063 13923
rect 6454 13920 6460 13932
rect 6051 13892 6132 13920
rect 6051 13889 6063 13892
rect 6005 13883 6063 13889
rect 3344 13824 4200 13852
rect 4249 13855 4307 13861
rect 2133 13815 2191 13821
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 5920 13852 5948 13880
rect 6104 13852 6132 13892
rect 6380 13892 6460 13920
rect 6380 13861 6408 13892
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 6632 13923 6690 13929
rect 6632 13889 6644 13923
rect 6678 13920 6690 13923
rect 7742 13920 7748 13932
rect 6678 13892 7748 13920
rect 6678 13889 6690 13892
rect 6632 13883 6690 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 4295 13824 5948 13852
rect 6012 13824 6132 13852
rect 6365 13855 6423 13861
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 6012 13796 6040 13824
rect 6365 13821 6377 13855
rect 6411 13821 6423 13855
rect 8036 13852 8064 13883
rect 9030 13880 9036 13932
rect 9088 13920 9094 13932
rect 10137 13923 10195 13929
rect 9088 13892 9628 13920
rect 9088 13880 9094 13892
rect 9600 13861 9628 13892
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10336 13920 10364 14019
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11698 14056 11704 14068
rect 11379 14028 11704 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 12802 14016 12808 14068
rect 12860 14016 12866 14068
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 10336 13892 10425 13920
rect 10137 13883 10195 13889
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10413 13883 10471 13889
rect 10520 13892 11713 13920
rect 6365 13815 6423 13821
rect 7760 13824 8064 13852
rect 9585 13855 9643 13861
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13753 1639 13787
rect 1581 13747 1639 13753
rect 5626 13744 5632 13796
rect 5684 13744 5690 13796
rect 5994 13744 6000 13796
rect 6052 13744 6058 13796
rect 2498 13676 2504 13728
rect 2556 13676 2562 13728
rect 3602 13676 3608 13728
rect 3660 13676 3666 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4709 13719 4767 13725
rect 4709 13716 4721 13719
rect 4580 13688 4721 13716
rect 4580 13676 4586 13688
rect 4709 13685 4721 13688
rect 4755 13685 4767 13719
rect 5644 13716 5672 13744
rect 6380 13716 6408 13815
rect 5644 13688 6408 13716
rect 4709 13679 4767 13685
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 7760 13725 7788 13824
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 10152 13852 10180 13883
rect 10520 13852 10548 13892
rect 11701 13889 11713 13892
rect 11747 13920 11759 13923
rect 11900 13920 11928 14016
rect 12060 13991 12118 13997
rect 12060 13957 12072 13991
rect 12106 13988 12118 13991
rect 12820 13988 12848 14016
rect 12106 13960 12848 13988
rect 12106 13957 12118 13960
rect 12060 13951 12118 13957
rect 11747 13892 11928 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 14458 13880 14464 13932
rect 14516 13880 14522 13932
rect 10152 13824 10548 13852
rect 9585 13815 9643 13821
rect 9600 13784 9628 13815
rect 10686 13812 10692 13864
rect 10744 13812 10750 13864
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13852 10931 13855
rect 11609 13855 11667 13861
rect 11609 13852 11621 13855
rect 10919 13824 11621 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 11609 13821 11621 13824
rect 11655 13821 11667 13855
rect 11609 13815 11667 13821
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 11808 13784 11836 13812
rect 9600 13756 11836 13784
rect 7745 13719 7803 13725
rect 7745 13716 7757 13719
rect 7616 13688 7757 13716
rect 7616 13676 7622 13688
rect 7745 13685 7757 13688
rect 7791 13685 7803 13719
rect 7745 13679 7803 13685
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 12584 13688 13185 13716
rect 12584 13676 12590 13688
rect 13173 13685 13185 13688
rect 13219 13685 13231 13719
rect 13173 13679 13231 13685
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 1811 13484 3556 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13413 2375 13447
rect 2317 13407 2375 13413
rect 2593 13447 2651 13453
rect 2593 13413 2605 13447
rect 2639 13444 2651 13447
rect 3528 13444 3556 13484
rect 3602 13472 3608 13524
rect 3660 13472 3666 13524
rect 3712 13484 7328 13512
rect 3712 13444 3740 13484
rect 5258 13444 5264 13456
rect 2639 13416 2774 13444
rect 3528 13416 3740 13444
rect 3896 13416 4844 13444
rect 2639 13413 2651 13416
rect 2593 13407 2651 13413
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1636 13280 1685 13308
rect 1636 13268 1642 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1673 13271 1731 13277
rect 1964 13280 2145 13308
rect 1964 13184 1992 13280
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2332 13308 2360 13407
rect 2746 13376 2774 13416
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2746 13348 3157 13376
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2332 13280 2421 13308
rect 2133 13271 2191 13277
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3050 13308 3056 13320
rect 3007 13280 3056 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 2884 13240 2912 13271
rect 3050 13268 3056 13280
rect 3108 13308 3114 13320
rect 3418 13308 3424 13320
rect 3108 13280 3424 13308
rect 3108 13268 3114 13280
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 3896 13240 3924 13416
rect 4816 13388 4844 13416
rect 4908 13416 5264 13444
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4120 13348 4292 13376
rect 4120 13336 4126 13348
rect 4264 13317 4292 13348
rect 4798 13336 4804 13388
rect 4856 13336 4862 13388
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 4522 13308 4528 13320
rect 4387 13280 4528 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 2884 13212 3924 13240
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 1946 13132 1952 13184
rect 2004 13132 2010 13184
rect 2774 13132 2780 13184
rect 2832 13132 2838 13184
rect 3786 13132 3792 13184
rect 3844 13132 3850 13184
rect 3988 13172 4016 13271
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4908 13317 4936 13416
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 6641 13447 6699 13453
rect 6641 13413 6653 13447
rect 6687 13444 6699 13447
rect 7190 13444 7196 13456
rect 6687 13416 7196 13444
rect 6687 13413 6699 13416
rect 6641 13407 6699 13413
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 7300 13444 7328 13484
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 7800 13484 8953 13512
rect 7800 13472 7806 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10502 13512 10508 13524
rect 10367 13484 10508 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10502 13472 10508 13484
rect 10560 13512 10566 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10560 13484 10793 13512
rect 10560 13472 10566 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 10781 13475 10839 13481
rect 11698 13472 11704 13524
rect 11756 13472 11762 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 13630 13512 13636 13524
rect 13495 13484 13636 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 7300 13416 10732 13444
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5537 13379 5595 13385
rect 5537 13376 5549 13379
rect 5031 13348 5549 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 5537 13345 5549 13348
rect 5583 13345 5595 13379
rect 7558 13376 7564 13388
rect 5537 13339 5595 13345
rect 6380 13348 7564 13376
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4663 13280 4905 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6380 13308 6408 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 7837 13379 7895 13385
rect 7837 13376 7849 13379
rect 7708 13348 7849 13376
rect 7708 13336 7714 13348
rect 7837 13345 7849 13348
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 8294 13336 8300 13388
rect 8352 13336 8358 13388
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 6236 13280 6408 13308
rect 6236 13268 6242 13280
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 8754 13268 8760 13320
rect 8812 13268 8818 13320
rect 8846 13268 8852 13320
rect 8904 13308 8910 13320
rect 9306 13308 9312 13320
rect 8904 13280 9312 13308
rect 8904 13268 8910 13280
rect 9306 13268 9312 13280
rect 9364 13308 9370 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9364 13280 9505 13308
rect 9364 13268 9370 13280
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 10410 13268 10416 13320
rect 10468 13268 10474 13320
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 10704 13308 10732 13416
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11112 13348 11345 13376
rect 11112 13336 11118 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11848 13348 12081 13376
rect 11848 13336 11854 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10704 13280 11161 13308
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 14182 13308 14188 13320
rect 11149 13271 11207 13277
rect 11256 13280 14188 13308
rect 6917 13243 6975 13249
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 7098 13240 7104 13252
rect 6963 13212 7104 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 7929 13243 7987 13249
rect 7929 13209 7941 13243
rect 7975 13240 7987 13243
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 7975 13212 8677 13240
rect 7975 13209 7987 13212
rect 7929 13203 7987 13209
rect 8665 13209 8677 13212
rect 8711 13209 8723 13243
rect 8665 13203 8723 13209
rect 10502 13200 10508 13252
rect 10560 13240 10566 13252
rect 11256 13240 11284 13280
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 10560 13212 11284 13240
rect 12336 13243 12394 13249
rect 10560 13200 10566 13212
rect 12336 13209 12348 13243
rect 12382 13240 12394 13243
rect 13998 13240 14004 13252
rect 12382 13212 14004 13240
rect 12382 13209 12394 13212
rect 12336 13203 12394 13209
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 3988 13144 4077 13172
rect 4065 13141 4077 13144
rect 4111 13141 4123 13175
rect 4065 13135 4123 13141
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 4706 13172 4712 13184
rect 4571 13144 4712 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4798 13132 4804 13184
rect 4856 13132 4862 13184
rect 5997 13175 6055 13181
rect 5997 13141 6009 13175
rect 6043 13172 6055 13175
rect 6086 13172 6092 13184
rect 6043 13144 6092 13172
rect 6043 13141 6055 13144
rect 5997 13135 6055 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 7006 13132 7012 13184
rect 7064 13132 7070 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 11940 13144 13645 13172
rect 11940 13132 11946 13144
rect 13633 13141 13645 13144
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 2498 12928 2504 12980
rect 2556 12928 2562 12980
rect 2774 12968 2780 12980
rect 2746 12928 2780 12968
rect 2832 12928 2838 12980
rect 4356 12940 7880 12968
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2746 12832 2774 12928
rect 4356 12909 4384 12940
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12869 4399 12903
rect 4341 12863 4399 12869
rect 4706 12860 4712 12912
rect 4764 12900 4770 12912
rect 5353 12903 5411 12909
rect 5353 12900 5365 12903
rect 4764 12872 5365 12900
rect 4764 12860 4770 12872
rect 5353 12869 5365 12872
rect 5399 12869 5411 12903
rect 6178 12900 6184 12912
rect 5353 12863 5411 12869
rect 6012 12872 6184 12900
rect 1903 12804 2774 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 1780 12764 1808 12795
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 6012 12841 6040 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 6328 12872 6592 12900
rect 6328 12860 6334 12872
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4212 12804 4445 12832
rect 4212 12792 4218 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6144 12804 6377 12832
rect 6144 12792 6150 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6454 12792 6460 12844
rect 6512 12792 6518 12844
rect 6564 12841 6592 12872
rect 7098 12860 7104 12912
rect 7156 12860 7162 12912
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7852 12909 7880 12940
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 9088 12940 9137 12968
rect 9088 12928 9094 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9732 12940 9781 12968
rect 9732 12928 9738 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 10413 12971 10471 12977
rect 9769 12931 9827 12937
rect 9876 12940 10180 12968
rect 7837 12903 7895 12909
rect 7248 12872 7328 12900
rect 7248 12860 7254 12872
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 1946 12764 1952 12776
rect 1780 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12733 2099 12767
rect 2041 12727 2099 12733
rect 1673 12699 1731 12705
rect 1673 12665 1685 12699
rect 1719 12696 1731 12699
rect 2056 12696 2084 12727
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 5442 12764 5448 12776
rect 5307 12736 5448 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5534 12724 5540 12776
rect 5592 12724 5598 12776
rect 1719 12668 2084 12696
rect 3053 12699 3111 12705
rect 1719 12665 1731 12668
rect 1673 12659 1731 12665
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 5626 12696 5632 12708
rect 3099 12668 5632 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 6181 12699 6239 12705
rect 6181 12665 6193 12699
rect 6227 12696 6239 12699
rect 6472 12696 6500 12792
rect 7116 12773 7144 12860
rect 7300 12841 7328 12872
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 8202 12900 8208 12912
rect 7883 12872 8208 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 9876 12900 9904 12940
rect 8312 12872 9904 12900
rect 10152 12900 10180 12940
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 10594 12968 10600 12980
rect 10459 12940 10600 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12032 12940 13308 12968
rect 12032 12928 12038 12940
rect 11992 12900 12020 12928
rect 10152 12872 12020 12900
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 8312 12696 8340 12872
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 6227 12668 6500 12696
rect 6564 12668 8340 12696
rect 6227 12665 6239 12668
rect 6181 12659 6239 12665
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4764 12600 4813 12628
rect 4764 12588 4770 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 6564 12628 6592 12668
rect 4948 12600 6592 12628
rect 7009 12631 7067 12637
rect 4948 12588 4954 12600
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7466 12628 7472 12640
rect 7055 12600 7472 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 9876 12628 9904 12795
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 10152 12804 10241 12832
rect 10152 12705 10180 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11882 12832 11888 12844
rect 11379 12804 11888 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 13096 12804 13185 12832
rect 13096 12776 13124 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 10137 12699 10195 12705
rect 10137 12665 10149 12699
rect 10183 12665 10195 12699
rect 10137 12659 10195 12665
rect 10502 12656 10508 12708
rect 10560 12656 10566 12708
rect 11164 12696 11192 12727
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 13078 12724 13084 12776
rect 13136 12724 13142 12776
rect 13280 12764 13308 12940
rect 13354 12792 13360 12844
rect 13412 12792 13418 12844
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 13280 12736 14197 12764
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14185 12727 14243 12733
rect 14458 12724 14464 12776
rect 14516 12724 14522 12776
rect 14090 12696 14096 12708
rect 11164 12668 13124 12696
rect 10520 12628 10548 12656
rect 9876 12600 10548 12628
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12628 11023 12631
rect 11698 12628 11704 12640
rect 11011 12600 11704 12628
rect 11011 12597 11023 12600
rect 10965 12591 11023 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 11882 12588 11888 12640
rect 11940 12588 11946 12640
rect 12618 12588 12624 12640
rect 12676 12588 12682 12640
rect 13096 12628 13124 12668
rect 13372 12668 14096 12696
rect 13372 12628 13400 12668
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 13096 12600 13400 12628
rect 13446 12588 13452 12640
rect 13504 12588 13510 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4706 12424 4712 12436
rect 4479 12396 4712 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5994 12384 6000 12436
rect 6052 12384 6058 12436
rect 6104 12396 9260 12424
rect 3513 12359 3571 12365
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 4522 12356 4528 12368
rect 3559 12328 4528 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 4522 12316 4528 12328
rect 4580 12316 4586 12368
rect 6104 12356 6132 12396
rect 4816 12328 6132 12356
rect 2498 12248 2504 12300
rect 2556 12288 2562 12300
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 2556 12260 2605 12288
rect 2556 12248 2562 12260
rect 2593 12257 2605 12260
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3660 12260 3801 12288
rect 3660 12248 3666 12260
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 3970 12248 3976 12300
rect 4028 12248 4034 12300
rect 1578 12180 1584 12232
rect 1636 12180 1642 12232
rect 2774 12180 2780 12232
rect 2832 12180 2838 12232
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 3384 12192 3433 12220
rect 3384 12180 3390 12192
rect 3421 12189 3433 12192
rect 3467 12220 3479 12223
rect 4062 12220 4068 12232
rect 3467 12192 4068 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 4816 12152 4844 12328
rect 7558 12316 7564 12368
rect 7616 12356 7622 12368
rect 8754 12356 8760 12368
rect 7616 12328 8760 12356
rect 7616 12316 7622 12328
rect 8754 12316 8760 12328
rect 8812 12356 8818 12368
rect 9125 12359 9183 12365
rect 8812 12328 8984 12356
rect 8812 12316 8818 12328
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 5684 12260 6377 12288
rect 5684 12248 5690 12260
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7524 12260 7941 12288
rect 7524 12248 7530 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8294 12248 8300 12300
rect 8352 12248 8358 12300
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5258 12180 5264 12232
rect 5316 12180 5322 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 5399 12192 5549 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 6632 12223 6690 12229
rect 6632 12189 6644 12223
rect 6678 12220 6690 12223
rect 7006 12220 7012 12232
rect 6678 12192 7012 12220
rect 6678 12189 6690 12192
rect 6632 12183 6690 12189
rect 5736 12152 5764 12183
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 8956 12229 8984 12328
rect 9125 12325 9137 12359
rect 9171 12325 9183 12359
rect 9232 12356 9260 12396
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 9364 12396 10885 12424
rect 9364 12384 9370 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 14090 12384 14096 12436
rect 14148 12384 14154 12436
rect 9232 12328 11284 12356
rect 9125 12319 9183 12325
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12189 8999 12223
rect 9140 12220 9168 12319
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10410 12288 10416 12300
rect 10100 12260 10416 12288
rect 10100 12248 10106 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9140 12192 9413 12220
rect 8941 12183 8999 12189
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 11146 12220 11152 12232
rect 10275 12192 11152 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 1688 12124 4844 12152
rect 4908 12124 5764 12152
rect 8021 12155 8079 12161
rect 1688 12093 1716 12124
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12053 1731 12087
rect 1673 12047 1731 12053
rect 2406 12044 2412 12096
rect 2464 12044 2470 12096
rect 3234 12044 3240 12096
rect 3292 12044 3298 12096
rect 4908 12093 4936 12124
rect 8021 12121 8033 12155
rect 8067 12121 8079 12155
rect 9784 12152 9812 12183
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11256 12220 11284 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13170 12356 13176 12368
rect 12768 12328 13176 12356
rect 12768 12316 12774 12328
rect 13170 12316 13176 12328
rect 13228 12356 13234 12368
rect 13265 12359 13323 12365
rect 13265 12356 13277 12359
rect 13228 12328 13277 12356
rect 13228 12316 13234 12328
rect 13265 12325 13277 12328
rect 13311 12325 13323 12359
rect 13265 12319 13323 12325
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 13446 12288 13452 12300
rect 12575 12260 13452 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 13630 12248 13636 12300
rect 13688 12288 13694 12300
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13688 12260 13829 12288
rect 13688 12248 13694 12260
rect 13817 12257 13829 12260
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 11256 12192 12357 12220
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 10778 12152 10784 12164
rect 9784 12124 10784 12152
rect 8021 12115 8079 12121
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5810 12084 5816 12096
rect 5215 12056 5816 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7616 12056 7757 12084
rect 7616 12044 7622 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 8036 12084 8064 12115
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 12008 12155 12066 12161
rect 12008 12121 12020 12155
rect 12054 12152 12066 12155
rect 12636 12152 12664 12180
rect 12054 12124 12664 12152
rect 12054 12121 12066 12124
rect 12008 12115 12066 12121
rect 13722 12112 13728 12164
rect 13780 12112 13786 12164
rect 14292 12152 14320 12183
rect 13924 12124 14320 12152
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8036 12056 9229 12084
rect 7745 12047 7803 12053
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 9953 12087 10011 12093
rect 9953 12053 9965 12087
rect 9999 12084 10011 12087
rect 10502 12084 10508 12096
rect 9999 12056 10508 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11054 12084 11060 12096
rect 10744 12056 11060 12084
rect 10744 12044 10750 12056
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12342 12084 12348 12096
rect 11756 12056 12348 12084
rect 11756 12044 11762 12056
rect 12342 12044 12348 12056
rect 12400 12084 12406 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12400 12056 13001 12084
rect 12400 12044 12406 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 13924 12084 13952 12124
rect 13596 12056 13952 12084
rect 13596 12044 13602 12056
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 2774 11880 2780 11892
rect 1903 11852 2780 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4203 11852 4936 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 2685 11815 2743 11821
rect 2685 11781 2697 11815
rect 2731 11812 2743 11815
rect 3022 11815 3080 11821
rect 3022 11812 3034 11815
rect 2731 11784 3034 11812
rect 2731 11781 2743 11784
rect 2685 11775 2743 11781
rect 3022 11781 3034 11784
rect 3068 11781 3080 11815
rect 3022 11775 3080 11781
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1544 11716 1777 11744
rect 1544 11704 1550 11716
rect 1765 11713 1777 11716
rect 1811 11744 1823 11747
rect 2133 11747 2191 11753
rect 2133 11744 2145 11747
rect 1811 11716 2145 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2133 11713 2145 11716
rect 2179 11744 2191 11747
rect 3326 11744 3332 11756
rect 2179 11716 3332 11744
rect 2179 11713 2191 11716
rect 2133 11707 2191 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 4908 11753 4936 11852
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 10100 11852 10333 11880
rect 10100 11840 10106 11852
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 10321 11843 10379 11849
rect 10597 11883 10655 11889
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 10686 11880 10692 11892
rect 10643 11852 10692 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 10836 11852 11529 11880
rect 10836 11840 10842 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 13262 11880 13268 11892
rect 13219 11852 13268 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14016 11852 14289 11880
rect 6914 11772 6920 11824
rect 6972 11772 6978 11824
rect 9048 11812 9076 11840
rect 12250 11812 12256 11824
rect 8772 11784 12256 11812
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 5074 11744 5080 11756
rect 4939 11716 5080 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5074 11704 5080 11716
rect 5132 11744 5138 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 5132 11716 5273 11744
rect 5132 11704 5138 11716
rect 5261 11713 5273 11716
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 8478 11744 8484 11756
rect 5408 11716 8484 11744
rect 5408 11704 5414 11716
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 8772 11753 8800 11784
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 9013 11747 9071 11753
rect 9013 11744 9025 11747
rect 8757 11707 8815 11713
rect 8864 11716 9025 11744
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 1578 11500 1584 11552
rect 1636 11500 1642 11552
rect 2792 11540 2820 11639
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 8864 11676 8892 11716
rect 9013 11713 9025 11716
rect 9059 11713 9071 11747
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 9013 11707 9071 11713
rect 9784 11716 10425 11744
rect 7524 11648 8892 11676
rect 7524 11636 7530 11648
rect 3970 11568 3976 11620
rect 4028 11608 4034 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4028 11580 5089 11608
rect 4028 11568 4034 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 7650 11608 7656 11620
rect 7432 11580 7656 11608
rect 7432 11568 7438 11580
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 8128 11580 8800 11608
rect 3050 11540 3056 11552
rect 2792 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4304 11512 4353 11540
rect 4304 11500 4310 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 4982 11500 4988 11552
rect 5040 11540 5046 11552
rect 8128 11540 8156 11580
rect 5040 11512 8156 11540
rect 5040 11500 5046 11512
rect 8202 11500 8208 11552
rect 8260 11500 8266 11552
rect 8772 11540 8800 11580
rect 9784 11540 9812 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10560 11716 11069 11744
rect 10560 11704 10566 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11744 11299 11747
rect 11514 11744 11520 11756
rect 11287 11716 11520 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11808 11753 11836 11784
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 14016 11821 14044 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 14001 11815 14059 11821
rect 12400 11784 12756 11812
rect 12400 11772 12406 11784
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 12060 11747 12118 11753
rect 12060 11713 12072 11747
rect 12106 11744 12118 11747
rect 12618 11744 12624 11756
rect 12106 11716 12624 11744
rect 12106 11713 12118 11716
rect 12060 11707 12118 11713
rect 11716 11676 11744 11707
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12728 11744 12756 11784
rect 14001 11781 14013 11815
rect 14047 11781 14059 11815
rect 14001 11775 14059 11781
rect 12728 11716 12848 11744
rect 10980 11648 11744 11676
rect 12820 11676 12848 11716
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13449 11747 13507 11753
rect 13449 11744 13461 11747
rect 13228 11716 13461 11744
rect 13228 11704 13234 11716
rect 13449 11713 13461 11716
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11744 14519 11747
rect 14507 11716 14872 11744
rect 14507 11713 14519 11716
rect 14461 11707 14519 11713
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 12820 11648 14105 11676
rect 10980 11620 11008 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 10137 11611 10195 11617
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 10318 11608 10324 11620
rect 10183 11580 10324 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10318 11568 10324 11580
rect 10376 11608 10382 11620
rect 10962 11608 10968 11620
rect 10376 11580 10968 11608
rect 10376 11568 10382 11580
rect 10962 11568 10968 11580
rect 11020 11568 11026 11620
rect 12434 11540 12440 11552
rect 8772 11512 12440 11540
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 1486 11336 1492 11348
rect 1443 11308 1492 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 1578 11296 1584 11348
rect 1636 11336 1642 11348
rect 4982 11336 4988 11348
rect 1636 11308 4988 11336
rect 1636 11296 1642 11308
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 5074 11296 5080 11348
rect 5132 11296 5138 11348
rect 5629 11339 5687 11345
rect 5629 11305 5641 11339
rect 5675 11305 5687 11339
rect 8386 11336 8392 11348
rect 5629 11299 5687 11305
rect 6932 11308 8392 11336
rect 4154 11228 4160 11280
rect 4212 11228 4218 11280
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3050 11200 3056 11212
rect 2823 11172 3056 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3050 11160 3056 11172
rect 3108 11200 3114 11212
rect 4172 11200 4200 11228
rect 3108 11172 4200 11200
rect 3108 11160 3114 11172
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 5092 11141 5120 11296
rect 5644 11268 5672 11299
rect 6932 11277 6960 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 11974 11336 11980 11348
rect 8536 11308 10364 11336
rect 8536 11296 8542 11308
rect 6457 11271 6515 11277
rect 5644 11240 6224 11268
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 6196 11200 6224 11240
rect 6457 11237 6469 11271
rect 6503 11268 6515 11271
rect 6917 11271 6975 11277
rect 6917 11268 6929 11271
rect 6503 11240 6929 11268
rect 6503 11237 6515 11240
rect 6457 11231 6515 11237
rect 6917 11237 6929 11240
rect 6963 11237 6975 11271
rect 8757 11271 8815 11277
rect 6917 11231 6975 11237
rect 7392 11240 8340 11268
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 5224 11172 5672 11200
rect 6196 11172 6745 11200
rect 5224 11160 5230 11172
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11134 5503 11135
rect 5534 11134 5540 11144
rect 5491 11106 5540 11134
rect 5491 11101 5503 11106
rect 5445 11095 5503 11101
rect 5534 11092 5540 11106
rect 5592 11092 5598 11144
rect 5644 11132 5672 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 7392 11200 7420 11240
rect 7576 11209 7656 11212
rect 6733 11163 6791 11169
rect 6932 11172 7420 11200
rect 7559 11203 7656 11209
rect 6932 11144 6960 11172
rect 7559 11169 7571 11203
rect 7605 11184 7656 11203
rect 7605 11169 7617 11184
rect 7559 11163 7617 11169
rect 7650 11160 7656 11184
rect 7708 11160 7714 11212
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 5644 11104 5825 11132
rect 5813 11101 5825 11104
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 2498 11024 2504 11076
rect 2556 11073 2562 11076
rect 2556 11027 2568 11073
rect 2961 11067 3019 11073
rect 2961 11033 2973 11067
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 3053 11067 3111 11073
rect 3053 11033 3065 11067
rect 3099 11064 3111 11067
rect 3605 11067 3663 11073
rect 3099 11036 3556 11064
rect 3099 11033 3111 11036
rect 3053 11027 3111 11033
rect 2556 11024 2562 11027
rect 2976 10996 3004 11027
rect 3234 10996 3240 11008
rect 2976 10968 3240 10996
rect 3234 10956 3240 10968
rect 3292 10956 3298 11008
rect 3528 10996 3556 11036
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 4062 11064 4068 11076
rect 3651 11036 4068 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4617 11067 4675 11073
rect 4617 11033 4629 11067
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 3789 10999 3847 11005
rect 3789 10996 3801 10999
rect 3528 10968 3801 10996
rect 3789 10965 3801 10968
rect 3835 10965 3847 10999
rect 4632 10996 4660 11027
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 4985 11067 5043 11073
rect 4985 11064 4997 11067
rect 4816 11036 4997 11064
rect 4816 10996 4844 11036
rect 4985 11033 4997 11036
rect 5031 11033 5043 11067
rect 4985 11027 5043 11033
rect 4632 10968 4844 10996
rect 3789 10959 3847 10965
rect 5258 10956 5264 11008
rect 5316 10956 5322 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 6012 10996 6040 11095
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6512 11104 6561 11132
rect 6512 11092 6518 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 8312 11141 8340 11240
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 10226 11268 10232 11280
rect 8803 11240 10232 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 10336 11268 10364 11308
rect 10796 11308 11980 11336
rect 10796 11268 10824 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 12124 11308 12357 11336
rect 12124 11296 12130 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 12618 11296 12624 11348
rect 12676 11296 12682 11348
rect 13262 11296 13268 11348
rect 13320 11296 13326 11348
rect 13538 11296 13544 11348
rect 13596 11296 13602 11348
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 14844 11336 14872 11716
rect 13863 11308 14872 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 10336 11240 10824 11268
rect 11054 11228 11060 11280
rect 11112 11228 11118 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 11204 11240 12173 11268
rect 11204 11228 11210 11240
rect 12161 11237 12173 11240
rect 12207 11237 12219 11271
rect 12161 11231 12219 11237
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8435 11172 9137 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 11072 11200 11100 11228
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 10183 11172 10640 11200
rect 11072 11172 11345 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7484 11104 7757 11132
rect 7484 11005 7512 11104
rect 7745 11101 7757 11104
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8343 11104 8585 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8720 11104 8953 11132
rect 8720 11092 8726 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10502 11132 10508 11144
rect 10367 11104 10508 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 9585 11067 9643 11073
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 9674 11064 9680 11076
rect 9631 11036 9680 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 10612 11064 10640 11172
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11606 11160 11612 11212
rect 11664 11160 11670 11212
rect 13280 11200 13308 11296
rect 13740 11268 13768 11296
rect 14185 11271 14243 11277
rect 14185 11268 14197 11271
rect 13740 11240 14197 11268
rect 14185 11237 14197 11240
rect 14231 11237 14243 11271
rect 14185 11231 14243 11237
rect 13280 11172 13676 11200
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 12069 11135 12127 11141
rect 11020 11104 11192 11132
rect 11020 11092 11026 11104
rect 11054 11064 11060 11076
rect 10612 11036 11060 11064
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11164 11064 11192 11104
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 13265 11135 13323 11141
rect 12575 11104 12756 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 11425 11067 11483 11073
rect 11164 11036 11376 11064
rect 5684 10968 6040 10996
rect 7469 10999 7527 11005
rect 5684 10956 5690 10968
rect 7469 10965 7481 10999
rect 7515 10965 7527 10999
rect 7469 10959 7527 10965
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 7708 10968 8217 10996
rect 7708 10956 7714 10968
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 11348 10996 11376 11036
rect 11425 11033 11437 11067
rect 11471 11064 11483 11067
rect 11698 11064 11704 11076
rect 11471 11036 11704 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 12084 11064 12112 11095
rect 11808 11036 12112 11064
rect 11808 10996 11836 11036
rect 12728 11008 12756 11104
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13354 11132 13360 11144
rect 13311 11104 13360 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13648 11141 13676 11172
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13679 11104 14105 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 11348 10968 11836 10996
rect 8205 10959 8263 10965
rect 12710 10956 12716 11008
rect 12768 10956 12774 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 2498 10752 2504 10804
rect 2556 10752 2562 10804
rect 3234 10752 3240 10804
rect 3292 10752 3298 10804
rect 10226 10752 10232 10804
rect 10284 10752 10290 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11112 10764 11529 10792
rect 11112 10752 11118 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 13354 10792 13360 10804
rect 13219 10764 13360 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 1854 10684 1860 10736
rect 1912 10724 1918 10736
rect 1912 10696 2774 10724
rect 1912 10684 1918 10696
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 2464 10628 2605 10656
rect 2464 10616 2470 10628
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 2746 10656 2774 10696
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 4402 10727 4460 10733
rect 4402 10724 4414 10727
rect 4304 10696 4414 10724
rect 4304 10684 4310 10696
rect 4402 10693 4414 10696
rect 4448 10693 4460 10727
rect 8662 10724 8668 10736
rect 4402 10687 4460 10693
rect 7392 10696 8668 10724
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2746 10628 3341 10656
rect 2593 10619 2651 10625
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 5902 10616 5908 10668
rect 5960 10616 5966 10668
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6362 10656 6368 10668
rect 6043 10628 6368 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6687 10628 7021 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2777 10591 2835 10597
rect 2777 10588 2789 10591
rect 2556 10560 2789 10588
rect 2556 10548 2562 10560
rect 2777 10557 2789 10560
rect 2823 10557 2835 10591
rect 2777 10551 2835 10557
rect 4154 10548 4160 10600
rect 4212 10548 4218 10600
rect 6564 10532 6592 10619
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7392 10588 7420 10696
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7650 10656 7656 10668
rect 7515 10628 7656 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7650 10616 7656 10628
rect 7708 10656 7714 10668
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 7708 10628 8309 10656
rect 7708 10616 7714 10628
rect 8297 10625 8309 10628
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8444 10628 9045 10656
rect 8444 10616 8450 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10244 10656 10272 10752
rect 11882 10684 11888 10736
rect 11940 10724 11946 10736
rect 12038 10727 12096 10733
rect 12038 10724 12050 10727
rect 11940 10696 12050 10724
rect 11940 10684 11946 10696
rect 12038 10693 12050 10696
rect 12084 10693 12096 10727
rect 12038 10687 12096 10693
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 12768 10696 14228 10724
rect 12768 10684 12774 10696
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 9732 10628 10180 10656
rect 10244 10628 11713 10656
rect 9732 10616 9738 10628
rect 6880 10560 7420 10588
rect 6880 10548 6886 10560
rect 7558 10548 7564 10600
rect 7616 10588 7622 10600
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 7616 10560 8125 10588
rect 7616 10548 7622 10560
rect 8113 10557 8125 10560
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 8478 10548 8484 10600
rect 8536 10548 8542 10600
rect 9214 10548 9220 10600
rect 9272 10548 9278 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6546 10520 6552 10532
rect 5592 10492 6552 10520
rect 5592 10480 5598 10492
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 9876 10520 9904 10551
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 10152 10588 10180 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 14200 10665 14228 10696
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 12492 10628 13277 10656
rect 12492 10616 12498 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10152 10560 10609 10588
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10778 10548 10784 10600
rect 10836 10548 10842 10600
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 6788 10492 9904 10520
rect 10244 10492 11100 10520
rect 6788 10480 6794 10492
rect 10244 10464 10272 10492
rect 3418 10412 3424 10464
rect 3476 10412 3482 10464
rect 5718 10412 5724 10464
rect 5776 10412 5782 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 6052 10424 6101 10452
rect 6052 10412 6058 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6822 10452 6828 10464
rect 6420 10424 6828 10452
rect 6420 10412 6426 10424
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7558 10412 7564 10464
rect 7616 10412 7622 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9677 10455 9735 10461
rect 9677 10452 9689 10455
rect 8987 10424 9689 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9677 10421 9689 10424
rect 9723 10452 9735 10455
rect 9950 10452 9956 10464
rect 9723 10424 9956 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10226 10412 10232 10464
rect 10284 10412 10290 10464
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 10962 10452 10968 10464
rect 10551 10424 10968 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11072 10452 11100 10492
rect 12802 10452 12808 10464
rect 11072 10424 12808 10452
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 13906 10452 13912 10464
rect 13495 10424 13912 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 2498 10208 2504 10260
rect 2556 10208 2562 10260
rect 3418 10208 3424 10260
rect 3476 10208 3482 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5626 10248 5632 10260
rect 5307 10220 5632 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 5718 10208 5724 10260
rect 5776 10208 5782 10260
rect 5994 10208 6000 10260
rect 6052 10208 6058 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8478 10248 8484 10260
rect 8435 10220 8484 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9214 10248 9220 10260
rect 9079 10220 9220 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 10100 10220 10149 10248
rect 10100 10208 10106 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10778 10208 10784 10260
rect 10836 10208 10842 10260
rect 10962 10208 10968 10260
rect 11020 10208 11026 10260
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 11756 10220 12173 10248
rect 11756 10208 11762 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 13127 10220 13461 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13449 10217 13461 10220
rect 13495 10248 13507 10251
rect 13630 10248 13636 10260
rect 13495 10220 13636 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 2593 10183 2651 10189
rect 2593 10149 2605 10183
rect 2639 10149 2651 10183
rect 3436 10180 3464 10208
rect 3436 10152 5488 10180
rect 2593 10143 2651 10149
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2608 10044 2636 10143
rect 3326 10112 3332 10124
rect 2792 10084 3332 10112
rect 2792 10053 2820 10084
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 5224 10084 5365 10112
rect 5224 10072 5230 10084
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 2363 10016 2636 10044
rect 2777 10047 2835 10053
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 3142 10044 3148 10056
rect 2915 10016 3148 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5258 10044 5264 10056
rect 5123 10016 5264 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5460 10044 5488 10152
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10112 5595 10115
rect 5736 10112 5764 10208
rect 5583 10084 5764 10112
rect 6012 10112 6040 10208
rect 6730 10140 6736 10192
rect 6788 10140 6794 10192
rect 10226 10180 10232 10192
rect 8128 10152 10232 10180
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 6012 10084 6285 10112
rect 5583 10081 5595 10084
rect 5537 10075 5595 10081
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5460 10016 6101 10044
rect 6089 10013 6101 10016
rect 6135 10044 6147 10047
rect 6454 10044 6460 10056
rect 6135 10016 6460 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1489 9979 1547 9985
rect 1489 9976 1501 9979
rect 992 9948 1501 9976
rect 992 9936 998 9948
rect 1489 9945 1501 9948
rect 1535 9945 1547 9979
rect 1489 9939 1547 9945
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 5997 9979 6055 9985
rect 1719 9948 5948 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 4798 9908 4804 9920
rect 3007 9880 4804 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5920 9908 5948 9948
rect 5997 9945 6009 9979
rect 6043 9976 6055 9979
rect 6748 9976 6776 10140
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6914 10044 6920 10056
rect 6871 10016 6920 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7098 9985 7104 9988
rect 6043 9948 6776 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 7092 9939 7104 9985
rect 7098 9936 7104 9939
rect 7156 9936 7162 9988
rect 8128 9908 8156 10152
rect 9232 10124 9260 10152
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 10505 10183 10563 10189
rect 10505 10149 10517 10183
rect 10551 10149 10563 10183
rect 10505 10143 10563 10149
rect 9214 10072 9220 10124
rect 9272 10072 9278 10124
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10318 10044 10324 10056
rect 10275 10016 10324 10044
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 8846 9976 8852 9988
rect 8220 9948 8852 9976
rect 8220 9917 8248 9948
rect 8846 9936 8852 9948
rect 8904 9976 8910 9988
rect 8956 9976 8984 10007
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10520 10044 10548 10143
rect 10980 10112 11008 10208
rect 11606 10140 11612 10192
rect 11664 10140 11670 10192
rect 12069 10183 12127 10189
rect 12069 10149 12081 10183
rect 12115 10149 12127 10183
rect 12069 10143 12127 10149
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 10980 10084 11161 10112
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11624 10112 11652 10140
rect 11563 10084 11652 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10520 10016 10609 10044
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 12084 10044 12112 10143
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 12084 10016 12357 10044
rect 11885 10007 11943 10013
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 8904 9948 8984 9976
rect 11241 9979 11299 9985
rect 8904 9936 8910 9948
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 11606 9976 11612 9988
rect 11287 9948 11612 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 11900 9920 11928 10007
rect 12434 10004 12440 10056
rect 12492 10004 12498 10056
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12802 10044 12808 10056
rect 12667 10016 12808 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13630 10004 13636 10056
rect 13688 10004 13694 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13780 10016 13829 10044
rect 13780 10004 13786 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 14918 10044 14924 10056
rect 14507 10016 14924 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 5920 9880 8156 9908
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 11882 9868 11888 9920
rect 11940 9868 11946 9920
rect 14274 9868 14280 9920
rect 14332 9868 14338 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 5902 9664 5908 9716
rect 5960 9664 5966 9716
rect 7009 9707 7067 9713
rect 7009 9673 7021 9707
rect 7055 9704 7067 9707
rect 7098 9704 7104 9716
rect 7055 9676 7104 9704
rect 7055 9673 7067 9676
rect 7009 9667 7067 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 9692 9676 10272 9704
rect 4448 9608 7236 9636
rect 4448 9580 4476 9608
rect 1394 9528 1400 9580
rect 1452 9528 1458 9580
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2130 9568 2136 9580
rect 1903 9540 2136 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 3878 9528 3884 9580
rect 3936 9577 3942 9580
rect 3936 9531 3948 9577
rect 3936 9528 3942 9531
rect 4430 9528 4436 9580
rect 4488 9528 4494 9580
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6546 9568 6552 9580
rect 6503 9540 6552 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 1811 9472 2421 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 2556 9472 2605 9500
rect 2556 9460 2562 9472
rect 2593 9469 2605 9472
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 5736 9500 5764 9531
rect 6546 9528 6552 9540
rect 6604 9568 6610 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6604 9540 7113 9568
rect 6604 9528 6610 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7208 9568 7236 9608
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7524 9608 8217 9636
rect 7524 9596 7530 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 9692 9636 9720 9676
rect 10134 9636 10140 9648
rect 8205 9599 8263 9605
rect 8312 9608 9720 9636
rect 9784 9608 10140 9636
rect 8312 9568 8340 9608
rect 7208 9540 8340 9568
rect 7101 9531 7159 9537
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 9784 9577 9812 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 10244 9636 10272 9676
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 12345 9707 12403 9713
rect 12345 9704 12357 9707
rect 11664 9676 12357 9704
rect 11664 9664 11670 9676
rect 12345 9673 12357 9676
rect 12391 9673 12403 9707
rect 12710 9704 12716 9716
rect 12345 9667 12403 9673
rect 12544 9676 12716 9704
rect 12544 9636 12572 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 13722 9704 13728 9716
rect 13280 9676 13728 9704
rect 13280 9648 13308 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 14274 9664 14280 9716
rect 14332 9664 14338 9716
rect 10244 9608 10548 9636
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9456 9540 9781 9568
rect 9456 9528 9462 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10036 9571 10094 9577
rect 10036 9537 10048 9571
rect 10082 9568 10094 9571
rect 10410 9568 10416 9580
rect 10082 9540 10416 9568
rect 10082 9537 10094 9540
rect 10036 9531 10094 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10520 9568 10548 9608
rect 10704 9608 12572 9636
rect 10704 9568 10732 9608
rect 12618 9596 12624 9648
rect 12676 9596 12682 9648
rect 13262 9596 13268 9648
rect 13320 9596 13326 9648
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 10520 9540 10732 9568
rect 12084 9540 12265 9568
rect 6822 9500 6828 9512
rect 5736 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9500 6886 9512
rect 7466 9500 7472 9512
rect 6880 9472 7472 9500
rect 6880 9460 6886 9472
rect 7466 9460 7472 9472
rect 7524 9500 7530 9512
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 7524 9472 7573 9500
rect 7524 9460 7530 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 9364 9472 9505 9500
rect 9364 9460 9370 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 11790 9500 11796 9512
rect 10796 9472 11796 9500
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2004 9404 2789 9432
rect 2004 9392 2010 9404
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 2777 9395 2835 9401
rect 7282 9392 7288 9444
rect 7340 9392 7346 9444
rect 1578 9324 1584 9376
rect 1636 9324 1642 9376
rect 2222 9324 2228 9376
rect 2280 9324 2286 9376
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8386 9364 8392 9376
rect 8343 9336 8392 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9309 9367 9367 9373
rect 9309 9333 9321 9367
rect 9355 9364 9367 9367
rect 10042 9364 10048 9376
rect 9355 9336 10048 9364
rect 9355 9333 9367 9336
rect 9309 9327 9367 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10796 9364 10824 9472
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 12084 9509 12112 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12636 9568 12664 9596
rect 14292 9577 14320 9664
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 12636 9540 12817 9568
rect 12529 9531 12587 9537
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 12805 9531 12863 9537
rect 13004 9540 14197 9568
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 12544 9500 12572 9531
rect 12544 9472 12848 9500
rect 12069 9463 12127 9469
rect 11149 9435 11207 9441
rect 11149 9401 11161 9435
rect 11195 9432 11207 9435
rect 11882 9432 11888 9444
rect 11195 9404 11888 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 11882 9392 11888 9404
rect 11940 9432 11946 9444
rect 12084 9432 12112 9463
rect 11940 9404 12112 9432
rect 11940 9392 11946 9404
rect 10192 9336 10824 9364
rect 11517 9367 11575 9373
rect 10192 9324 10198 9336
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 11606 9364 11612 9376
rect 11563 9336 11612 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 12820 9364 12848 9472
rect 13004 9441 13032 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 13955 9472 14381 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 12989 9435 13047 9441
rect 12989 9401 13001 9435
rect 13035 9401 13047 9435
rect 13740 9432 13768 9463
rect 14001 9435 14059 9441
rect 14001 9432 14013 9435
rect 13740 9404 14013 9432
rect 12989 9395 13047 9401
rect 14001 9401 14013 9404
rect 14047 9401 14059 9435
rect 14001 9395 14059 9401
rect 13354 9364 13360 9376
rect 12820 9336 13360 9364
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 1578 9120 1584 9172
rect 1636 9120 1642 9172
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2280 9132 2329 9160
rect 2280 9120 2286 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2556 9132 2881 9160
rect 2556 9120 2562 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 4430 9160 4436 9172
rect 2869 9123 2927 9129
rect 2976 9132 4436 9160
rect 1596 9024 1624 9120
rect 2133 9027 2191 9033
rect 2133 9024 2145 9027
rect 1596 8996 2145 9024
rect 2133 8993 2145 8996
rect 2179 8993 2191 9027
rect 2133 8987 2191 8993
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2976 8965 3004 9132
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 6880 9132 8309 9160
rect 6880 9120 6886 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8570 9160 8576 9172
rect 8527 9132 8576 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9364 9132 9413 9160
rect 9364 9120 9370 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 12710 9120 12716 9172
rect 12768 9120 12774 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12860 9132 13093 9160
rect 12860 9120 12866 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 13262 9120 13268 9172
rect 13320 9120 13326 9172
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9160 13507 9163
rect 13630 9160 13636 9172
rect 13495 9132 13636 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 3973 9095 4031 9101
rect 3973 9061 3985 9095
rect 4019 9061 4031 9095
rect 3973 9055 4031 9061
rect 4249 9095 4307 9101
rect 4249 9061 4261 9095
rect 4295 9092 4307 9095
rect 4295 9064 4568 9092
rect 4295 9061 4307 9064
rect 4249 9055 4307 9061
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1728 8928 1961 8956
rect 1728 8916 1734 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8925 3019 8959
rect 2961 8919 3019 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3988 8956 4016 9055
rect 4540 9033 4568 9064
rect 4614 9052 4620 9104
rect 4672 9092 4678 9104
rect 5350 9092 5356 9104
rect 4672 9064 5356 9092
rect 4672 9052 4678 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 5537 9095 5595 9101
rect 5537 9061 5549 9095
rect 5583 9061 5595 9095
rect 5537 9055 5595 9061
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 5552 9024 5580 9055
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 4948 8996 5488 9024
rect 5552 8996 5825 9024
rect 4948 8984 4954 8996
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3988 8928 4077 8956
rect 3789 8919 3847 8925
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4908 8956 4936 8984
rect 4387 8928 4936 8956
rect 5261 8959 5319 8965
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1489 8891 1547 8897
rect 1489 8888 1501 8891
rect 992 8860 1501 8888
rect 992 8848 998 8860
rect 1489 8857 1501 8860
rect 1535 8857 1547 8891
rect 1489 8851 1547 8857
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 3804 8888 3832 8919
rect 5276 8888 5304 8919
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5460 8956 5488 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5460 8928 5641 8956
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 6454 8956 6460 8968
rect 5629 8919 5687 8925
rect 5727 8928 6460 8956
rect 5727 8888 5755 8928
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6840 8956 6868 9120
rect 6595 8928 6868 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7650 8956 7656 8968
rect 6972 8928 7656 8956
rect 6972 8916 6978 8928
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8956 8723 8959
rect 8846 8956 8852 8968
rect 8711 8928 8852 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 8846 8916 8852 8928
rect 8904 8956 8910 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8904 8928 9321 8956
rect 8904 8916 8910 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 9815 8928 10272 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 7006 8888 7012 8900
rect 2188 8860 5755 8888
rect 6288 8860 7012 8888
rect 2188 8848 2194 8860
rect 6288 8832 6316 8860
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 7184 8891 7242 8897
rect 7184 8857 7196 8891
rect 7230 8888 7242 8891
rect 7558 8888 7564 8900
rect 7230 8860 7564 8888
rect 7230 8857 7242 8860
rect 7184 8851 7242 8857
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 7668 8860 9689 8888
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 4614 8820 4620 8832
rect 1627 8792 4620 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 4982 8780 4988 8832
rect 5040 8780 5046 8832
rect 5166 8780 5172 8832
rect 5224 8780 5230 8832
rect 6270 8780 6276 8832
rect 6328 8780 6334 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7668 8820 7696 8860
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 9677 8851 9735 8857
rect 10244 8888 10272 8928
rect 11606 8916 11612 8968
rect 11664 8965 11670 8968
rect 11664 8956 11676 8965
rect 11664 8928 11709 8956
rect 11664 8919 11676 8928
rect 11664 8916 11670 8919
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11848 8928 11897 8956
rect 11848 8916 11854 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12216 8928 12357 8956
rect 12216 8916 12222 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12728 8956 12756 9120
rect 12989 9095 13047 9101
rect 12989 9061 13001 9095
rect 13035 9092 13047 9095
rect 13280 9092 13308 9120
rect 13035 9064 13308 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 12860 8996 13676 9024
rect 12860 8984 12866 8996
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 12728 8928 13277 8956
rect 12529 8919 12587 8925
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 12544 8888 12572 8919
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 13648 8965 13676 8996
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 15010 8956 15016 8968
rect 14323 8928 15016 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 13725 8891 13783 8897
rect 13725 8888 13737 8891
rect 10244 8860 12434 8888
rect 12544 8860 13737 8888
rect 10244 8832 10272 8860
rect 7432 8792 7696 8820
rect 7432 8780 7438 8792
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 10686 8820 10692 8832
rect 10551 8792 10692 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 12406 8820 12434 8860
rect 13725 8857 13737 8860
rect 13771 8857 13783 8891
rect 13725 8851 13783 8857
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 12406 8792 14105 8820
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 3326 8616 3332 8628
rect 1995 8588 3332 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3694 8576 3700 8628
rect 3752 8576 3758 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 3878 8616 3884 8628
rect 3835 8588 3884 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4982 8616 4988 8628
rect 4571 8588 4988 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 3712 8548 3740 8576
rect 1627 8520 3740 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 2004 8452 2053 8480
rect 2004 8440 2010 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2179 8452 2513 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4540 8480 4568 8579
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5408 8588 5457 8616
rect 5408 8576 5414 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 5445 8579 5503 8585
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6270 8616 6276 8628
rect 6227 8588 6276 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6454 8576 6460 8628
rect 6512 8576 6518 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 9122 8616 9128 8628
rect 8067 8588 9128 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 3743 8452 4568 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5184 8480 5212 8576
rect 5031 8452 5212 8480
rect 5261 8483 5319 8489
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5721 8483 5779 8489
rect 5307 8452 5672 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 2280 8384 2329 8412
rect 2280 8372 2286 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 3660 8384 4353 8412
rect 3660 8372 3666 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4816 8412 4844 8440
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4816 8384 5181 8412
rect 4341 8375 4399 8381
rect 5169 8381 5181 8384
rect 5215 8412 5227 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5215 8384 5549 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5644 8412 5672 8452
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6472 8480 6500 8576
rect 6656 8548 6684 8576
rect 6656 8520 6868 8548
rect 5767 8452 6500 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6546 8440 6552 8492
rect 6604 8478 6610 8492
rect 6840 8489 6868 8520
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 9769 8551 9827 8557
rect 7708 8520 9444 8548
rect 7708 8508 7714 8520
rect 6825 8483 6883 8489
rect 6604 8450 6647 8478
rect 6604 8440 6610 8450
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 8128 8489 8156 8520
rect 9416 8492 9444 8520
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 9858 8548 9864 8560
rect 9815 8520 9864 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 10100 8520 10517 8548
rect 10100 8508 10106 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 10505 8511 10563 8517
rect 10594 8508 10600 8560
rect 10652 8508 10658 8560
rect 8386 8489 8392 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 6972 8452 7757 8480
rect 6972 8440 6978 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8380 8480 8392 8489
rect 8347 8452 8392 8480
rect 8113 8443 8171 8449
rect 8380 8443 8392 8452
rect 6932 8412 6960 8440
rect 5644 8384 6960 8412
rect 7009 8415 7067 8421
rect 5537 8375 5595 8381
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 7055 8384 7665 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3234 8344 3240 8356
rect 3007 8316 3240 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 5074 8344 5080 8356
rect 3375 8316 5080 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6914 8344 6920 8356
rect 6687 8316 6920 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7190 8304 7196 8356
rect 7248 8304 7254 8356
rect 7852 8344 7880 8443
rect 8386 8440 8392 8443
rect 8444 8440 8450 8492
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 11698 8440 11704 8492
rect 11756 8480 11762 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 11756 8452 14105 8480
rect 11756 8440 11762 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9950 8412 9956 8424
rect 9723 8384 9956 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 9493 8347 9551 8353
rect 7852 8316 8156 8344
rect 8128 8276 8156 8316
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 9539 8316 9674 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 8478 8276 8484 8288
rect 8128 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 9646 8276 9674 8316
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 10192 8316 10241 8344
rect 10192 8304 10198 8316
rect 10229 8313 10241 8316
rect 10275 8344 10287 8347
rect 10796 8344 10824 8375
rect 12066 8372 12072 8424
rect 12124 8372 12130 8424
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 12216 8384 12265 8412
rect 12216 8372 12222 8384
rect 12253 8381 12265 8384
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 10275 8316 10824 8344
rect 10275 8313 10287 8316
rect 10229 8307 10287 8313
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14185 8347 14243 8353
rect 14185 8344 14197 8347
rect 13872 8316 14197 8344
rect 13872 8304 13878 8316
rect 14185 8313 14197 8316
rect 14231 8313 14243 8347
rect 14185 8307 14243 8313
rect 9950 8276 9956 8288
rect 9646 8248 9956 8276
rect 9950 8236 9956 8248
rect 10008 8276 10014 8288
rect 10410 8276 10416 8288
rect 10008 8248 10416 8276
rect 10008 8236 10014 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 11606 8236 11612 8288
rect 11664 8236 11670 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1452 8044 1593 8072
rect 1452 8032 1458 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3568 8044 3985 8072
rect 3568 8032 3574 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 9858 8032 9864 8084
rect 9916 8032 9922 8084
rect 10042 8032 10048 8084
rect 10100 8032 10106 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10594 8072 10600 8084
rect 10275 8044 10600 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 11609 8075 11667 8081
rect 11609 8041 11621 8075
rect 11655 8072 11667 8075
rect 12066 8072 12072 8084
rect 11655 8044 12072 8072
rect 11655 8041 11667 8044
rect 11609 8035 11667 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 2130 7964 2136 8016
rect 2188 7964 2194 8016
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 7973 4399 8007
rect 4341 7967 4399 7973
rect 9677 8007 9735 8013
rect 9677 7973 9689 8007
rect 9723 8004 9735 8007
rect 10060 8004 10088 8032
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9723 7976 10088 8004
rect 10244 7976 10333 8004
rect 9723 7973 9735 7976
rect 9677 7967 9735 7973
rect 2148 7936 2176 7964
rect 1780 7908 2176 7936
rect 4356 7936 4384 7967
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 4356 7908 5733 7936
rect 1780 7877 1808 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 6696 7908 6745 7936
rect 6696 7896 6702 7908
rect 6733 7905 6745 7908
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6914 7896 6920 7948
rect 6972 7896 6978 7948
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 9180 7908 9229 7936
rect 9180 7896 9186 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 3142 7868 3148 7880
rect 2179 7840 3148 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4246 7868 4252 7880
rect 4203 7840 4252 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 2400 7803 2458 7809
rect 2400 7769 2412 7803
rect 2446 7800 2458 7803
rect 2498 7800 2504 7812
rect 2446 7772 2504 7800
rect 2446 7769 2458 7772
rect 2400 7763 2458 7769
rect 2498 7760 2504 7772
rect 2556 7760 2562 7812
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 4080 7800 4108 7831
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6822 7868 6828 7880
rect 6595 7840 6828 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 2740 7772 4108 7800
rect 2740 7760 2746 7772
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 3050 7732 3056 7744
rect 2087 7704 3056 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 3510 7692 3516 7744
rect 3568 7692 3574 7744
rect 4080 7732 4108 7772
rect 4433 7803 4491 7809
rect 4433 7769 4445 7803
rect 4479 7800 4491 7803
rect 4890 7800 4896 7812
rect 4479 7772 4896 7800
rect 4479 7769 4491 7772
rect 4433 7763 4491 7769
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 4982 7760 4988 7812
rect 5040 7760 5046 7812
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 5132 7772 5273 7800
rect 5132 7760 5138 7772
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 5920 7800 5948 7831
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7156 7840 7665 7868
rect 7156 7828 7162 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8846 7868 8852 7880
rect 8711 7840 8852 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9876 7868 9904 7896
rect 9945 7873 10003 7879
rect 9945 7868 9957 7873
rect 9876 7840 9957 7868
rect 9945 7839 9957 7840
rect 9991 7839 10003 7873
rect 9945 7833 10003 7839
rect 10069 7871 10127 7877
rect 10069 7837 10081 7871
rect 10115 7868 10127 7871
rect 10244 7868 10272 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 11333 8007 11391 8013
rect 11333 7973 11345 8007
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 10115 7840 10272 7868
rect 10115 7837 10127 7840
rect 10069 7831 10127 7837
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10468 7840 10517 7868
rect 10468 7828 10474 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 5920 7772 7389 7800
rect 5261 7763 5319 7769
rect 7377 7769 7389 7772
rect 7423 7800 7435 7803
rect 10520 7800 10548 7831
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 10744 7840 11161 7868
rect 10744 7828 10750 7840
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 11348 7868 11376 7967
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11348 7840 11437 7868
rect 11149 7831 11207 7837
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 7423 7772 9674 7800
rect 10520 7772 14228 7800
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 4798 7732 4804 7744
rect 4080 7704 4804 7732
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5994 7692 6000 7744
rect 6052 7692 6058 7744
rect 7466 7692 7472 7744
rect 7524 7692 7530 7744
rect 9646 7732 9674 7772
rect 14200 7744 14228 7772
rect 11606 7732 11612 7744
rect 9646 7704 11612 7732
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 14182 7692 14188 7744
rect 14240 7692 14246 7744
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 4982 7528 4988 7540
rect 4755 7500 4988 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9398 7528 9404 7540
rect 9355 7500 9404 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10686 7488 10692 7540
rect 10744 7488 10750 7540
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 4387 7432 7849 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 7837 7429 7849 7432
rect 7883 7460 7895 7463
rect 8202 7460 8208 7472
rect 7883 7432 8208 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2038 7392 2044 7404
rect 1627 7364 2044 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 3568 7364 4629 7392
rect 3568 7352 3574 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2700 7324 2728 7352
rect 2004 7296 2728 7324
rect 2004 7284 2010 7296
rect 5184 7256 5212 7355
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 7064 7364 7113 7392
rect 7064 7352 7070 7364
rect 7101 7361 7113 7364
rect 7147 7361 7159 7395
rect 10704 7392 10732 7488
rect 7101 7355 7159 7361
rect 7199 7364 10732 7392
rect 14461 7395 14519 7401
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6604 7296 6929 7324
rect 6604 7284 6610 7296
rect 6917 7293 6929 7296
rect 6963 7324 6975 7327
rect 7199 7324 7227 7364
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14507 7364 14964 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 6963 7296 7227 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 7282 7284 7288 7336
rect 7340 7284 7346 7336
rect 14936 7268 14964 7364
rect 10226 7256 10232 7268
rect 2746 7228 4016 7256
rect 5184 7228 10232 7256
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 2746 7188 2774 7228
rect 3988 7200 4016 7228
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 14918 7216 14924 7268
rect 14976 7216 14982 7268
rect 1811 7160 2774 7188
rect 3053 7191 3111 7197
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3142 7188 3148 7200
rect 3099 7160 3148 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3970 7148 3976 7200
rect 4028 7148 4034 7200
rect 4982 7148 4988 7200
rect 5040 7148 5046 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5868 7160 6377 7188
rect 5868 7148 5874 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 7432 7160 7481 7188
rect 7432 7148 7438 7160
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 1854 6984 1860 6996
rect 1443 6956 1860 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 1854 6944 1860 6956
rect 1912 6944 1918 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4617 6987 4675 6993
rect 4617 6984 4629 6987
rect 4304 6956 4629 6984
rect 4304 6944 4310 6956
rect 4617 6953 4629 6956
rect 4663 6953 4675 6987
rect 4617 6947 4675 6953
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7282 6984 7288 6996
rect 7055 6956 7288 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 3142 6848 3148 6860
rect 2823 6820 3148 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 3142 6808 3148 6820
rect 3200 6848 3206 6860
rect 4172 6848 4200 6876
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 3200 6820 5457 6848
rect 3200 6808 3206 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9398 6848 9404 6860
rect 8812 6820 9404 6848
rect 8812 6808 8818 6820
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9723 6820 9996 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9968 6792 9996 6820
rect 2521 6783 2579 6789
rect 2521 6749 2533 6783
rect 2567 6780 2579 6783
rect 2869 6783 2927 6789
rect 2567 6752 2774 6780
rect 2567 6749 2579 6752
rect 2521 6743 2579 6749
rect 2746 6644 2774 6752
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 2958 6780 2964 6792
rect 2915 6752 2964 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3068 6712 3096 6743
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3292 6752 3525 6780
rect 3292 6740 3298 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3326 6712 3332 6724
rect 3068 6684 3332 6712
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 3528 6712 3556 6743
rect 4798 6740 4804 6792
rect 4856 6740 4862 6792
rect 5712 6783 5770 6789
rect 5712 6749 5724 6783
rect 5758 6780 5770 6783
rect 5994 6780 6000 6792
rect 5758 6752 6000 6780
rect 5758 6749 5770 6752
rect 5712 6743 5770 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6840 6752 6929 6780
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3528 6684 3893 6712
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 3881 6675 3939 6681
rect 3970 6672 3976 6724
rect 4028 6672 4034 6724
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4525 6715 4583 6721
rect 4525 6712 4537 6715
rect 4212 6684 4537 6712
rect 4212 6672 4218 6684
rect 4525 6681 4537 6684
rect 4571 6712 4583 6715
rect 4890 6712 4896 6724
rect 4571 6684 4896 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 4890 6672 4896 6684
rect 4948 6672 4954 6724
rect 5810 6672 5816 6724
rect 5868 6672 5874 6724
rect 5828 6644 5856 6672
rect 2746 6616 5856 6644
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6840 6653 6868 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7432 6752 8616 6780
rect 7432 6740 7438 6752
rect 8478 6672 8484 6724
rect 8536 6721 8542 6724
rect 8536 6675 8548 6721
rect 8588 6712 8616 6752
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 9033 6715 9091 6721
rect 9033 6712 9045 6715
rect 8588 6684 9045 6712
rect 9033 6681 9045 6684
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 9125 6715 9183 6721
rect 9125 6681 9137 6715
rect 9171 6712 9183 6715
rect 10410 6712 10416 6724
rect 9171 6684 10416 6712
rect 9171 6681 9183 6684
rect 9125 6675 9183 6681
rect 8536 6672 8542 6675
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6696 6616 6837 6644
rect 6696 6604 6702 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7558 6644 7564 6656
rect 7423 6616 7564 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10042 6644 10048 6656
rect 9999 6616 10048 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 1762 6400 1768 6452
rect 1820 6400 1826 6452
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 3068 6412 7880 6440
rect 2240 6344 2728 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1854 6304 1860 6316
rect 1627 6276 1860 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 2240 6313 2268 6344
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 1210 6196 1216 6248
rect 1268 6236 1274 6248
rect 2332 6236 2360 6267
rect 1268 6208 2360 6236
rect 2700 6236 2728 6344
rect 3068 6313 3096 6412
rect 7852 6372 7880 6412
rect 8478 6400 8484 6452
rect 8536 6400 8542 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9824 6412 10364 6440
rect 9824 6400 9830 6412
rect 9401 6375 9459 6381
rect 6932 6344 7788 6372
rect 7852 6344 8892 6372
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2823 6276 3065 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6638 6304 6644 6316
rect 6411 6276 6644 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 6932 6313 6960 6344
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7184 6307 7242 6313
rect 7184 6273 7196 6307
rect 7230 6304 7242 6307
rect 7650 6304 7656 6316
rect 7230 6276 7656 6304
rect 7230 6273 7242 6276
rect 7184 6267 7242 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7760 6304 7788 6344
rect 8864 6316 8892 6344
rect 9401 6341 9413 6375
rect 9447 6372 9459 6375
rect 9447 6344 9996 6372
rect 9447 6341 9459 6344
rect 9401 6335 9459 6341
rect 8754 6304 8760 6316
rect 7760 6276 8760 6304
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9968 6304 9996 6344
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 10100 6344 10272 6372
rect 10100 6332 10106 6344
rect 10244 6313 10272 6344
rect 10336 6313 10364 6412
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10560 6412 10977 6440
rect 10560 6400 10566 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12158 6440 12164 6452
rect 12023 6412 12164 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 14292 6372 14320 6400
rect 10428 6344 14320 6372
rect 10229 6307 10287 6313
rect 9968 6276 10088 6304
rect 3510 6236 3516 6248
rect 2700 6208 3516 6236
rect 1268 6196 1274 6208
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 7024 6236 7052 6264
rect 6564 6208 7052 6236
rect 9033 6239 9091 6245
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6168 2743 6171
rect 3418 6168 3424 6180
rect 2731 6140 3424 6168
rect 2731 6137 2743 6140
rect 2685 6131 2743 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 6564 6177 6592 6208
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 6549 6171 6607 6177
rect 6549 6137 6561 6171
rect 6595 6137 6607 6171
rect 6549 6131 6607 6137
rect 8297 6171 8355 6177
rect 8297 6137 8309 6171
rect 8343 6168 8355 6171
rect 9048 6168 9076 6199
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9766 6168 9772 6180
rect 8343 6140 9772 6168
rect 8343 6137 8355 6140
rect 8297 6131 8355 6137
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 9861 6171 9919 6177
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 9950 6168 9956 6180
rect 9907 6140 9956 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10060 6177 10088 6276
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10045 6171 10103 6177
rect 10045 6137 10057 6171
rect 10091 6137 10103 6171
rect 10045 6131 10103 6137
rect 2498 6060 2504 6112
rect 2556 6060 2562 6112
rect 2866 6060 2872 6112
rect 2924 6060 2930 6112
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 7558 6100 7564 6112
rect 6779 6072 7564 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 10428 6100 10456 6344
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10796 6276 10885 6304
rect 10594 6196 10600 6248
rect 10652 6196 10658 6248
rect 10796 6112 10824 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 14461 6307 14519 6313
rect 12115 6276 14320 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12360 6112 12388 6276
rect 14292 6177 14320 6276
rect 14461 6273 14473 6307
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14476 6236 14504 6267
rect 14918 6236 14924 6248
rect 14476 6208 14924 6236
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 14277 6171 14335 6177
rect 14277 6137 14289 6171
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 8904 6072 10456 6100
rect 8904 6060 8910 6072
rect 10778 6060 10784 6112
rect 10836 6060 10842 6112
rect 12342 6060 12348 6112
rect 12400 6060 12406 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1544 5868 1593 5896
rect 1544 5856 1550 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2556 5868 7604 5896
rect 2556 5856 2562 5868
rect 6825 5831 6883 5837
rect 6825 5797 6837 5831
rect 6871 5797 6883 5831
rect 7576 5828 7604 5868
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 8757 5899 8815 5905
rect 7852 5868 8708 5896
rect 7852 5828 7880 5868
rect 7576 5800 7880 5828
rect 7929 5831 7987 5837
rect 6825 5791 6883 5797
rect 7929 5797 7941 5831
rect 7975 5797 7987 5831
rect 8680 5828 8708 5868
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 8803 5868 9229 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9217 5865 9229 5868
rect 9263 5896 9275 5899
rect 9306 5896 9312 5908
rect 9263 5868 9312 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10594 5856 10600 5908
rect 10652 5856 10658 5908
rect 8680 5800 9536 5828
rect 7929 5791 7987 5797
rect 6840 5760 6868 5791
rect 7944 5760 7972 5791
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 6840 5732 7788 5760
rect 7944 5732 9413 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6380 5624 6408 5655
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6696 5664 7021 5692
rect 6696 5652 6702 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7760 5701 7788 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8202 5692 8208 5704
rect 8159 5664 8208 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 9508 5692 9536 5800
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 10612 5760 10640 5856
rect 9631 5732 10640 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9508 5664 10057 5692
rect 8297 5655 8355 5661
rect 10045 5661 10057 5664
rect 10091 5692 10103 5695
rect 10778 5692 10784 5704
rect 10091 5664 10784 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 6822 5624 6828 5636
rect 6380 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 7576 5624 7604 5652
rect 8312 5624 8340 5655
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 7576 5596 8340 5624
rect 6549 5559 6607 5565
rect 6549 5525 6561 5559
rect 6595 5556 6607 5559
rect 6914 5556 6920 5568
rect 6595 5528 6920 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 12158 5516 12164 5568
rect 12216 5516 12222 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7190 5352 7196 5364
rect 7147 5324 7196 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8202 5312 8208 5364
rect 8260 5312 8266 5364
rect 5736 5256 6868 5284
rect 5736 5225 5764 5256
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5721 5179 5779 5185
rect 5920 5188 6009 5216
rect 5920 5089 5948 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6840 5160 6868 5256
rect 7208 5225 7236 5312
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8312 5188 8953 5216
rect 6454 5108 6460 5160
rect 6512 5108 6518 5160
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6656 5080 6684 5111
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 8312 5148 8340 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 12434 5176 12440 5228
rect 12492 5176 12498 5228
rect 6880 5120 8340 5148
rect 8665 5151 8723 5157
rect 6880 5108 6886 5120
rect 8665 5117 8677 5151
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 6227 5052 6684 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 7374 5040 7380 5092
rect 7432 5080 7438 5092
rect 7561 5083 7619 5089
rect 7561 5080 7573 5083
rect 7432 5052 7573 5080
rect 7432 5040 7438 5052
rect 7561 5049 7573 5052
rect 7607 5049 7619 5083
rect 8680 5080 8708 5111
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 12452 5148 12480 5176
rect 8904 5120 12480 5148
rect 8904 5108 8910 5120
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8680 5052 9045 5080
rect 7561 5043 7619 5049
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6512 4780 7021 4808
rect 6512 4768 6518 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8202 4808 8208 4820
rect 8159 4780 8208 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 8846 4808 8852 4820
rect 8711 4780 8852 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14415 4780 14872 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 14844 4752 14872 4780
rect 6914 4700 6920 4752
rect 6972 4700 6978 4752
rect 7377 4743 7435 4749
rect 7377 4709 7389 4743
rect 7423 4740 7435 4743
rect 7423 4712 7696 4740
rect 7423 4709 7435 4712
rect 7377 4703 7435 4709
rect 6932 4672 6960 4700
rect 7668 4681 7696 4712
rect 14826 4700 14832 4752
rect 14884 4700 14890 4752
rect 7653 4675 7711 4681
rect 6932 4644 7236 4672
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7208 4613 7236 4644
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 9214 4672 9220 4684
rect 7653 4635 7711 4641
rect 8404 4644 9220 4672
rect 8404 4613 8432 4644
rect 9214 4632 9220 4644
rect 9272 4672 9278 4684
rect 9272 4644 12480 4672
rect 9272 4632 9278 4644
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 7515 4576 8309 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8570 4564 8576 4616
rect 8628 4606 8634 4616
rect 8628 4578 8671 4606
rect 8628 4564 8634 4578
rect 12452 4548 12480 4644
rect 14182 4564 14188 4616
rect 14240 4564 14246 4616
rect 12434 4496 12440 4548
rect 12492 4496 12498 4548
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 14274 4468 14280 4480
rect 7340 4440 14280 4468
rect 7340 4428 7346 4440
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 8570 4060 8576 4072
rect 1636 4032 8576 4060
rect 1636 4020 1642 4032
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 8956 4060 8984 4091
rect 8628 4032 8984 4060
rect 8628 4020 8634 4032
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9858 3924 9864 3936
rect 9171 3896 9864 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5442 3720 5448 3732
rect 5307 3692 5448 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 13998 3680 14004 3732
rect 14056 3720 14062 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14056 3692 14289 3720
rect 14056 3680 14062 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3621 1639 3655
rect 1581 3615 1639 3621
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1596 3516 1624 3615
rect 5258 3516 5264 3528
rect 1596 3488 5264 3516
rect 1397 3479 1455 3485
rect 5258 3476 5264 3488
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14507 3488 14596 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 14568 3392 14596 3488
rect 14550 3340 14556 3392
rect 14608 3340 14614 3392
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 5258 3136 5264 3188
rect 5316 3136 5322 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10008 3148 10548 3176
rect 10008 3136 10014 3148
rect 4154 3108 4160 3120
rect 2148 3080 4160 3108
rect 2148 3049 2176 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3040 1823 3043
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 1811 3012 2053 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 5276 3049 5304 3136
rect 10318 3108 10324 3120
rect 6748 3080 10324 3108
rect 6748 3049 6776 3080
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 10134 3040 10140 3052
rect 9631 3012 10140 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10520 3049 10548 3148
rect 13633 3111 13691 3117
rect 13633 3077 13645 3111
rect 13679 3108 13691 3111
rect 13814 3108 13820 3120
rect 13679 3080 13820 3108
rect 13679 3077 13691 3080
rect 13633 3071 13691 3077
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 13906 3068 13912 3120
rect 13964 3068 13970 3120
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 11882 3000 11888 3052
rect 11940 3000 11946 3052
rect 12434 3000 12440 3052
rect 12492 3000 12498 3052
rect 14458 2904 14464 2916
rect 13556 2876 14464 2904
rect 474 2796 480 2848
rect 532 2836 538 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 532 2808 1501 2836
rect 532 2796 538 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 4154 2796 4160 2848
rect 4212 2796 4218 2848
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5994 2836 6000 2848
rect 5491 2808 6000 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6546 2796 6552 2848
rect 6604 2796 6610 2848
rect 8205 2839 8263 2845
rect 8205 2805 8217 2839
rect 8251 2836 8263 2839
rect 8386 2836 8392 2848
rect 8251 2808 8392 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 8536 2808 9505 2836
rect 8536 2796 8542 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 11146 2836 11152 2848
rect 10643 2808 11152 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12066 2796 12072 2848
rect 12124 2796 12130 2848
rect 12618 2796 12624 2848
rect 12676 2796 12682 2848
rect 13556 2845 13584 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2805 13599 2839
rect 13541 2799 13599 2805
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14001 2839 14059 2845
rect 14001 2836 14013 2839
rect 13780 2808 14013 2836
rect 13780 2796 13786 2808
rect 14001 2805 14013 2808
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 3050 2592 3056 2644
rect 3108 2592 3114 2644
rect 14274 2592 14280 2644
rect 14332 2592 14338 2644
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 3068 2428 3096 2592
rect 12158 2564 12164 2576
rect 2639 2400 3096 2428
rect 3160 2536 12164 2564
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 1360 2332 1409 2360
rect 1360 2320 1366 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 1780 2292 1808 2323
rect 2222 2320 2228 2372
rect 2280 2320 2286 2372
rect 3050 2320 3056 2372
rect 3108 2320 3114 2372
rect 3160 2292 3188 2536
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 3436 2468 5028 2496
rect 3436 2437 3464 2468
rect 5000 2440 5028 2468
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6052 2468 9076 2496
rect 6052 2456 6058 2468
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 4212 2400 4261 2428
rect 4212 2388 4218 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4982 2388 4988 2440
rect 5040 2388 5046 2440
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6604 2400 6745 2428
rect 6604 2388 6610 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9048 2437 9076 2468
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9858 2428 9864 2440
rect 9815 2400 9864 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10284 2400 10609 2428
rect 10284 2388 10290 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11204 2400 11621 2428
rect 11204 2388 11210 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 12124 2400 12265 2428
rect 12124 2388 12130 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12676 2400 13093 2428
rect 12676 2388 12682 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14507 2400 14596 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 3878 2320 3884 2372
rect 3936 2320 3942 2372
rect 6362 2320 6368 2372
rect 6420 2320 6426 2372
rect 7190 2320 7196 2372
rect 7248 2320 7254 2372
rect 7561 2363 7619 2369
rect 7561 2329 7573 2363
rect 7607 2360 7619 2363
rect 8496 2360 8524 2388
rect 7607 2332 8524 2360
rect 7607 2329 7619 2332
rect 7561 2323 7619 2329
rect 14568 2304 14596 2400
rect 1780 2264 3188 2292
rect 4890 2252 4896 2304
rect 4948 2252 4954 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5721 2295 5779 2301
rect 5721 2292 5733 2295
rect 5592 2264 5733 2292
rect 5592 2252 5598 2264
rect 5721 2261 5733 2264
rect 5767 2261 5779 2295
rect 5721 2255 5779 2261
rect 8113 2295 8171 2301
rect 8113 2261 8125 2295
rect 8159 2292 8171 2295
rect 8202 2292 8208 2304
rect 8159 2264 8208 2292
rect 8159 2261 8171 2264
rect 8113 2255 8171 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8812 2264 9137 2292
rect 8812 2252 8818 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9732 2264 9873 2292
rect 9732 2252 9738 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 10689 2295 10747 2301
rect 10689 2292 10701 2295
rect 10468 2264 10701 2292
rect 10468 2252 10474 2264
rect 10689 2261 10701 2264
rect 10735 2261 10747 2295
rect 10689 2255 10747 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12308 2264 12541 2292
rect 12308 2252 12314 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 14550 2252 14556 2304
rect 14608 2252 14614 2304
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
<< via1 >>
rect 7656 17756 7708 17808
rect 8300 17756 8352 17808
rect 3056 17552 3108 17604
rect 4620 17552 4672 17604
rect 3240 17484 3292 17536
rect 6644 17484 6696 17536
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 940 17280 992 17332
rect 2412 17280 2464 17332
rect 3148 17280 3200 17332
rect 3056 17212 3108 17264
rect 5356 17280 5408 17332
rect 6092 17280 6144 17332
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 7656 17280 7708 17332
rect 9036 17280 9088 17332
rect 9772 17280 9824 17332
rect 10508 17280 10560 17332
rect 11152 17280 11204 17332
rect 11980 17280 12032 17332
rect 12716 17280 12768 17332
rect 13452 17280 13504 17332
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 2964 16940 3016 16992
rect 3240 16940 3292 16992
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 6828 17076 6880 17128
rect 7756 17187 7808 17196
rect 7756 17153 7765 17187
rect 7765 17153 7799 17187
rect 7799 17153 7808 17187
rect 7756 17144 7808 17153
rect 11704 17212 11756 17264
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 7564 17076 7616 17128
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12624 17144 12676 17196
rect 13268 17144 13320 17196
rect 13728 17144 13780 17196
rect 12072 17076 12124 17128
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 4712 16940 4764 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 8392 16940 8444 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 11060 16940 11112 16992
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 1676 16736 1728 16788
rect 3056 16736 3108 16788
rect 4068 16736 4120 16788
rect 4528 16779 4580 16788
rect 4528 16745 4537 16779
rect 4537 16745 4571 16779
rect 4571 16745 4580 16779
rect 4528 16736 4580 16745
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 1768 16532 1820 16584
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3884 16643 3936 16652
rect 3884 16609 3893 16643
rect 3893 16609 3927 16643
rect 3927 16609 3936 16643
rect 3884 16600 3936 16609
rect 4160 16600 4212 16652
rect 5724 16600 5776 16652
rect 3516 16532 3568 16584
rect 3792 16464 3844 16516
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 4896 16464 4948 16516
rect 6000 16464 6052 16516
rect 6552 16464 6604 16516
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 9220 16736 9272 16788
rect 11704 16779 11756 16788
rect 11704 16745 11713 16779
rect 11713 16745 11747 16779
rect 11747 16745 11756 16779
rect 11704 16736 11756 16745
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 13268 16736 13320 16788
rect 13728 16736 13780 16788
rect 14188 16736 14240 16788
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 10784 16532 10836 16541
rect 11152 16532 11204 16584
rect 11980 16532 12032 16584
rect 12532 16668 12584 16720
rect 8484 16464 8536 16516
rect 9128 16507 9180 16516
rect 9128 16473 9137 16507
rect 9137 16473 9171 16507
rect 9171 16473 9180 16507
rect 9128 16464 9180 16473
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 10692 16464 10744 16516
rect 12532 16532 12584 16584
rect 13176 16668 13228 16720
rect 13636 16532 13688 16584
rect 13268 16464 13320 16516
rect 13544 16507 13596 16516
rect 13544 16473 13553 16507
rect 13553 16473 13587 16507
rect 13587 16473 13596 16507
rect 13544 16464 13596 16473
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2044 16396 2096 16405
rect 2872 16396 2924 16448
rect 3424 16396 3476 16448
rect 5080 16396 5132 16448
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7564 16439 7616 16448
rect 7564 16405 7573 16439
rect 7573 16405 7607 16439
rect 7607 16405 7616 16439
rect 7564 16396 7616 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 9772 16396 9824 16448
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 13728 16396 13780 16448
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 1768 16192 1820 16244
rect 3424 16192 3476 16244
rect 4988 16192 5040 16244
rect 5724 16192 5776 16244
rect 8300 16192 8352 16244
rect 1952 16056 2004 16108
rect 4252 16124 4304 16176
rect 4712 16124 4764 16176
rect 5264 16124 5316 16176
rect 5816 16124 5868 16176
rect 5448 16056 5500 16108
rect 8852 16099 8904 16108
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 3516 15852 3568 15904
rect 6552 15988 6604 16040
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9956 16192 10008 16244
rect 10692 16192 10744 16244
rect 10784 16192 10836 16244
rect 12164 16192 12216 16244
rect 12256 16192 12308 16244
rect 9772 16124 9824 16176
rect 13544 16192 13596 16244
rect 15016 16192 15068 16244
rect 9036 15988 9088 16040
rect 10416 16099 10468 16108
rect 10416 16065 10425 16099
rect 10425 16065 10459 16099
rect 10459 16065 10468 16099
rect 10416 16056 10468 16065
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 11060 15988 11112 16040
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 12348 16056 12400 16108
rect 13360 16056 13412 16108
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 6460 15852 6512 15904
rect 11060 15852 11112 15904
rect 11704 15852 11756 15904
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 13452 15852 13504 15861
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 2320 15648 2372 15700
rect 3148 15648 3200 15700
rect 4160 15691 4212 15700
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 4804 15648 4856 15700
rect 5448 15648 5500 15700
rect 3424 15512 3476 15564
rect 3516 15555 3568 15564
rect 3516 15521 3525 15555
rect 3525 15521 3559 15555
rect 3559 15521 3568 15555
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 9128 15648 9180 15700
rect 10692 15648 10744 15700
rect 11152 15648 11204 15700
rect 12808 15648 12860 15700
rect 13360 15648 13412 15700
rect 13452 15648 13504 15700
rect 3516 15512 3568 15521
rect 2964 15444 3016 15496
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 4712 15444 4764 15496
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 7564 15512 7616 15564
rect 8852 15512 8904 15564
rect 5448 15444 5500 15496
rect 7012 15444 7064 15496
rect 7472 15444 7524 15496
rect 8392 15444 8444 15496
rect 10600 15512 10652 15564
rect 4068 15376 4120 15428
rect 3332 15308 3384 15360
rect 5448 15351 5500 15360
rect 5448 15317 5457 15351
rect 5457 15317 5491 15351
rect 5491 15317 5500 15351
rect 5448 15308 5500 15317
rect 6460 15376 6512 15428
rect 7104 15376 7156 15428
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 11612 15444 11664 15496
rect 6920 15308 6972 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 9312 15308 9364 15360
rect 11704 15376 11756 15428
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 13728 15419 13780 15428
rect 13728 15385 13737 15419
rect 13737 15385 13771 15419
rect 13771 15385 13780 15419
rect 13728 15376 13780 15385
rect 13820 15419 13872 15428
rect 13820 15385 13829 15419
rect 13829 15385 13863 15419
rect 13863 15385 13872 15419
rect 13820 15376 13872 15385
rect 11244 15308 11296 15360
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 3056 15104 3108 15156
rect 3240 15104 3292 15156
rect 2228 15036 2280 15088
rect 3332 14968 3384 15020
rect 4344 15104 4396 15156
rect 10692 15104 10744 15156
rect 11612 15104 11664 15156
rect 12164 15104 12216 15156
rect 13360 15104 13412 15156
rect 13820 15104 13872 15156
rect 4804 15036 4856 15088
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 3608 14832 3660 14884
rect 4804 14832 4856 14884
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 6000 14832 6052 14884
rect 10416 14968 10468 15020
rect 11060 14968 11112 15020
rect 13360 14968 13412 15020
rect 14188 14968 14240 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 11888 14900 11940 14952
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5172 14764 5224 14816
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 7196 14764 7248 14816
rect 7840 14764 7892 14816
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9404 14764 9456 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 11704 14832 11756 14884
rect 13544 14900 13596 14952
rect 12440 14764 12492 14816
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 12808 14764 12860 14816
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 940 14356 992 14408
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 5264 14492 5316 14544
rect 5816 14560 5868 14612
rect 6828 14560 6880 14612
rect 7196 14560 7248 14612
rect 7748 14560 7800 14612
rect 8760 14560 8812 14612
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 5908 14492 5960 14544
rect 7104 14424 7156 14476
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 7840 14424 7892 14476
rect 9036 14467 9088 14476
rect 9036 14433 9045 14467
rect 9045 14433 9079 14467
rect 9079 14433 9088 14467
rect 9036 14424 9088 14433
rect 10048 14424 10100 14476
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 4160 14220 4212 14272
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 11244 14356 11296 14408
rect 11796 14356 11848 14408
rect 12716 14356 12768 14408
rect 14556 14356 14608 14408
rect 8852 14288 8904 14340
rect 9404 14288 9456 14340
rect 9864 14220 9916 14272
rect 11888 14220 11940 14272
rect 12440 14220 12492 14272
rect 13636 14220 13688 14272
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 1952 14016 2004 14068
rect 3424 14016 3476 14068
rect 3608 14016 3660 14068
rect 4804 14016 4856 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 6000 14016 6052 14068
rect 6184 14016 6236 14068
rect 6552 14016 6604 14068
rect 8760 14016 8812 14068
rect 2044 13880 2096 13932
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 9312 13991 9364 14000
rect 9312 13957 9330 13991
rect 9330 13957 9364 13991
rect 9312 13948 9364 13957
rect 5908 13880 5960 13932
rect 6460 13880 6512 13932
rect 7748 13880 7800 13932
rect 9036 13880 9088 13932
rect 11060 14016 11112 14068
rect 11704 14016 11756 14068
rect 11888 14016 11940 14068
rect 12808 14016 12860 14068
rect 5632 13744 5684 13796
rect 6000 13744 6052 13796
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 3608 13719 3660 13728
rect 3608 13685 3617 13719
rect 3617 13685 3651 13719
rect 3651 13685 3660 13719
rect 3608 13676 3660 13685
rect 4528 13676 4580 13728
rect 7564 13676 7616 13728
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 12532 13676 12584 13728
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 940 13268 992 13320
rect 1584 13268 1636 13320
rect 3056 13268 3108 13320
rect 3424 13268 3476 13320
rect 4068 13336 4120 13388
rect 4804 13336 4856 13388
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 1952 13132 2004 13184
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 2780 13132 2832 13141
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4528 13268 4580 13320
rect 5264 13404 5316 13456
rect 7196 13404 7248 13456
rect 7748 13472 7800 13524
rect 10508 13472 10560 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 13636 13472 13688 13524
rect 7564 13379 7616 13388
rect 5448 13268 5500 13320
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 7656 13336 7708 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 6184 13268 6236 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 8852 13268 8904 13320
rect 9312 13268 9364 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 11060 13336 11112 13388
rect 11796 13336 11848 13388
rect 7104 13200 7156 13252
rect 10508 13200 10560 13252
rect 14188 13268 14240 13320
rect 14004 13200 14056 13252
rect 4712 13132 4764 13184
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 6092 13132 6144 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 11888 13132 11940 13184
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 2780 12928 2832 12980
rect 4712 12860 4764 12912
rect 4160 12792 4212 12844
rect 6184 12860 6236 12912
rect 6276 12860 6328 12912
rect 6092 12792 6144 12844
rect 6460 12792 6512 12844
rect 7104 12860 7156 12912
rect 7196 12860 7248 12912
rect 9036 12928 9088 12980
rect 9680 12928 9732 12980
rect 1952 12724 2004 12776
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5448 12724 5500 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 5632 12656 5684 12708
rect 8208 12860 8260 12912
rect 10600 12928 10652 12980
rect 11980 12928 12032 12980
rect 4712 12588 4764 12640
rect 4896 12588 4948 12640
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 10048 12792 10100 12844
rect 11888 12792 11940 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 10508 12656 10560 12708
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13084 12724 13136 12776
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 11704 12588 11756 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 14096 12656 14148 12708
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 4712 12384 4764 12436
rect 6000 12427 6052 12436
rect 6000 12393 6009 12427
rect 6009 12393 6043 12427
rect 6043 12393 6052 12427
rect 6000 12384 6052 12393
rect 4528 12316 4580 12368
rect 2504 12248 2556 12300
rect 3608 12248 3660 12300
rect 3976 12291 4028 12300
rect 3976 12257 3985 12291
rect 3985 12257 4019 12291
rect 4019 12257 4028 12291
rect 3976 12248 4028 12257
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 2780 12223 2832 12232
rect 2780 12189 2789 12223
rect 2789 12189 2823 12223
rect 2823 12189 2832 12223
rect 2780 12180 2832 12189
rect 3332 12180 3384 12232
rect 4068 12180 4120 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 7564 12316 7616 12368
rect 8760 12316 8812 12368
rect 5632 12248 5684 12300
rect 7472 12248 7524 12300
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 7012 12180 7064 12232
rect 9312 12384 9364 12436
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10416 12248 10468 12300
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 11152 12180 11204 12232
rect 12716 12316 12768 12368
rect 13176 12316 13228 12368
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 13452 12248 13504 12300
rect 13636 12248 13688 12300
rect 12624 12180 12676 12232
rect 5816 12044 5868 12096
rect 7564 12044 7616 12096
rect 10784 12112 10836 12164
rect 13728 12155 13780 12164
rect 13728 12121 13737 12155
rect 13737 12121 13771 12155
rect 13771 12121 13780 12155
rect 13728 12112 13780 12121
rect 10508 12044 10560 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11060 12044 11112 12096
rect 11704 12044 11756 12096
rect 12348 12044 12400 12096
rect 13544 12044 13596 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 2780 11840 2832 11892
rect 940 11704 992 11756
rect 1492 11704 1544 11756
rect 3332 11704 3384 11756
rect 9036 11840 9088 11892
rect 10048 11840 10100 11892
rect 10692 11840 10744 11892
rect 10784 11840 10836 11892
rect 13268 11840 13320 11892
rect 6920 11815 6972 11824
rect 6920 11781 6929 11815
rect 6929 11781 6963 11815
rect 6963 11781 6972 11815
rect 6920 11772 6972 11781
rect 5080 11704 5132 11756
rect 5356 11704 5408 11756
rect 8484 11704 8536 11756
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 7472 11636 7524 11688
rect 3976 11568 4028 11620
rect 7380 11568 7432 11620
rect 7656 11568 7708 11620
rect 3056 11500 3108 11552
rect 4252 11500 4304 11552
rect 4988 11500 5040 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 10508 11704 10560 11756
rect 11520 11704 11572 11756
rect 12256 11772 12308 11824
rect 12348 11772 12400 11824
rect 12624 11704 12676 11756
rect 13176 11704 13228 11756
rect 10324 11568 10376 11620
rect 10968 11568 11020 11620
rect 12440 11500 12492 11552
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 1492 11296 1544 11348
rect 1584 11296 1636 11348
rect 4988 11296 5040 11348
rect 5080 11296 5132 11348
rect 4160 11228 4212 11280
rect 3056 11160 3108 11212
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 8392 11296 8444 11348
rect 8484 11296 8536 11348
rect 5172 11160 5224 11212
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 5540 11092 5592 11101
rect 7656 11160 7708 11212
rect 2504 11067 2556 11076
rect 2504 11033 2522 11067
rect 2522 11033 2556 11067
rect 2504 11024 2556 11033
rect 3240 10956 3292 11008
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 5632 10956 5684 11008
rect 6460 11092 6512 11144
rect 6920 11092 6972 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 10232 11228 10284 11280
rect 11980 11296 12032 11348
rect 12072 11296 12124 11348
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 13268 11296 13320 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 13728 11296 13780 11348
rect 11060 11228 11112 11280
rect 11152 11228 11204 11280
rect 8668 11092 8720 11144
rect 10508 11092 10560 11144
rect 9680 11067 9732 11076
rect 9680 11033 9689 11067
rect 9689 11033 9723 11067
rect 9723 11033 9732 11067
rect 9680 11024 9732 11033
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11060 11024 11112 11076
rect 7656 10956 7708 11008
rect 11704 11024 11756 11076
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 12716 10956 12768 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 10232 10752 10284 10804
rect 11060 10752 11112 10804
rect 13360 10752 13412 10804
rect 1860 10684 1912 10736
rect 2412 10616 2464 10668
rect 4252 10684 4304 10736
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 6368 10616 6420 10668
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2504 10548 2556 10600
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 8668 10684 8720 10736
rect 7656 10616 7708 10668
rect 8392 10616 8444 10668
rect 9680 10616 9732 10668
rect 11888 10684 11940 10736
rect 12716 10684 12768 10736
rect 6828 10548 6880 10557
rect 7564 10548 7616 10600
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 8484 10548 8536 10557
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 5540 10523 5592 10532
rect 5540 10489 5549 10523
rect 5549 10489 5583 10523
rect 5583 10489 5592 10523
rect 5540 10480 5592 10489
rect 6552 10480 6604 10532
rect 6736 10480 6788 10532
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 12440 10616 12492 10668
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6000 10412 6052 10464
rect 6368 10412 6420 10464
rect 6828 10412 6880 10464
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 9956 10412 10008 10464
rect 10232 10412 10284 10464
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 12808 10412 12860 10464
rect 13912 10412 13964 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 3424 10208 3476 10260
rect 5632 10208 5684 10260
rect 5724 10208 5776 10260
rect 6000 10208 6052 10260
rect 8484 10208 8536 10260
rect 9220 10208 9272 10260
rect 10048 10208 10100 10260
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 10968 10208 11020 10260
rect 11704 10208 11756 10260
rect 13636 10208 13688 10260
rect 3332 10072 3384 10124
rect 5172 10072 5224 10124
rect 3148 10004 3200 10056
rect 5264 10004 5316 10056
rect 6736 10183 6788 10192
rect 6736 10149 6745 10183
rect 6745 10149 6779 10183
rect 6779 10149 6788 10183
rect 6736 10140 6788 10149
rect 6460 10004 6512 10056
rect 940 9936 992 9988
rect 4804 9868 4856 9920
rect 6920 10004 6972 10056
rect 7104 9979 7156 9988
rect 7104 9945 7138 9979
rect 7138 9945 7156 9979
rect 7104 9936 7156 9945
rect 10232 10140 10284 10192
rect 9220 10072 9272 10124
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 10324 10047 10376 10056
rect 8852 9936 8904 9988
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 11612 10140 11664 10192
rect 11612 9936 11664 9988
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 12808 10004 12860 10056
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 13728 10004 13780 10056
rect 14924 10004 14976 10056
rect 11888 9868 11940 9920
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 7104 9664 7156 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2136 9528 2188 9580
rect 3884 9571 3936 9580
rect 3884 9537 3902 9571
rect 3902 9537 3936 9571
rect 3884 9528 3936 9537
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 2504 9460 2556 9512
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 6552 9528 6604 9580
rect 7472 9596 7524 9648
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 9404 9528 9456 9580
rect 10140 9596 10192 9648
rect 11612 9664 11664 9716
rect 12716 9664 12768 9716
rect 13728 9664 13780 9716
rect 14280 9664 14332 9716
rect 10416 9528 10468 9580
rect 12624 9596 12676 9648
rect 13268 9639 13320 9648
rect 13268 9605 13277 9639
rect 13277 9605 13311 9639
rect 13311 9605 13320 9639
rect 13268 9596 13320 9605
rect 6828 9460 6880 9512
rect 7472 9460 7524 9512
rect 9312 9460 9364 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 1952 9392 2004 9444
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 8392 9324 8444 9376
rect 10048 9324 10100 9376
rect 10140 9324 10192 9376
rect 11796 9460 11848 9512
rect 11888 9392 11940 9444
rect 11612 9324 11664 9376
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 13360 9324 13412 9376
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 1584 9120 1636 9172
rect 2228 9120 2280 9172
rect 2504 9120 2556 9172
rect 1676 8916 1728 8968
rect 4436 9120 4488 9172
rect 6828 9120 6880 9172
rect 8576 9120 8628 9172
rect 9312 9120 9364 9172
rect 12716 9120 12768 9172
rect 12808 9120 12860 9172
rect 13268 9120 13320 9172
rect 13636 9120 13688 9172
rect 4620 9052 4672 9104
rect 5356 9052 5408 9104
rect 4896 8984 4948 9036
rect 940 8848 992 8900
rect 2136 8848 2188 8900
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 6460 8916 6512 8968
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7656 8916 7708 8968
rect 8852 8916 8904 8968
rect 7012 8848 7064 8900
rect 7564 8848 7616 8900
rect 4620 8780 4672 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5172 8823 5224 8832
rect 5172 8789 5181 8823
rect 5181 8789 5215 8823
rect 5215 8789 5224 8823
rect 5172 8780 5224 8789
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 7380 8780 7432 8832
rect 11612 8959 11664 8968
rect 11612 8925 11630 8959
rect 11630 8925 11664 8959
rect 11612 8916 11664 8925
rect 11796 8916 11848 8968
rect 12164 8916 12216 8968
rect 12808 8984 12860 9036
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 15016 8916 15068 8968
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 10232 8780 10284 8832
rect 10692 8780 10744 8832
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 3332 8576 3384 8628
rect 3700 8576 3752 8628
rect 3884 8576 3936 8628
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 1952 8440 2004 8492
rect 4988 8576 5040 8628
rect 5172 8576 5224 8628
rect 5356 8576 5408 8628
rect 6276 8576 6328 8628
rect 6460 8576 6512 8628
rect 6644 8576 6696 8628
rect 9128 8576 9180 8628
rect 4804 8440 4856 8492
rect 2228 8372 2280 8424
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 3608 8372 3660 8424
rect 6552 8481 6604 8492
rect 6552 8447 6561 8481
rect 6561 8447 6595 8481
rect 6595 8447 6604 8481
rect 7656 8508 7708 8560
rect 6552 8440 6604 8447
rect 6920 8440 6972 8492
rect 9864 8508 9916 8560
rect 10048 8508 10100 8560
rect 10600 8551 10652 8560
rect 10600 8517 10609 8551
rect 10609 8517 10643 8551
rect 10643 8517 10652 8551
rect 10600 8508 10652 8517
rect 8392 8483 8444 8492
rect 8392 8449 8426 8483
rect 8426 8449 8444 8483
rect 3240 8304 3292 8356
rect 5080 8304 5132 8356
rect 6920 8304 6972 8356
rect 7196 8347 7248 8356
rect 7196 8313 7205 8347
rect 7205 8313 7239 8347
rect 7239 8313 7248 8347
rect 7196 8304 7248 8313
rect 8392 8440 8444 8449
rect 9404 8440 9456 8492
rect 11704 8440 11756 8492
rect 9956 8372 10008 8424
rect 8484 8236 8536 8288
rect 10140 8304 10192 8356
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 12164 8372 12216 8424
rect 13820 8304 13872 8356
rect 9956 8236 10008 8288
rect 10416 8236 10468 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 1400 8032 1452 8084
rect 3516 8032 3568 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 10048 8032 10100 8084
rect 10600 8032 10652 8084
rect 12072 8032 12124 8084
rect 2136 7964 2188 8016
rect 6644 7896 6696 7948
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 9128 7896 9180 7948
rect 9864 7896 9916 7948
rect 3148 7828 3200 7880
rect 2504 7760 2556 7812
rect 2688 7760 2740 7812
rect 4252 7828 4304 7880
rect 3056 7692 3108 7744
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4896 7760 4948 7812
rect 4988 7803 5040 7812
rect 4988 7769 4997 7803
rect 4997 7769 5031 7803
rect 5031 7769 5040 7803
rect 4988 7760 5040 7769
rect 5080 7803 5132 7812
rect 5080 7769 5089 7803
rect 5089 7769 5123 7803
rect 5123 7769 5132 7803
rect 5080 7760 5132 7769
rect 6828 7828 6880 7880
rect 7104 7828 7156 7880
rect 8852 7828 8904 7880
rect 10416 7828 10468 7880
rect 10692 7828 10744 7880
rect 4804 7692 4856 7744
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 11612 7692 11664 7744
rect 14188 7692 14240 7744
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 4988 7488 5040 7540
rect 9404 7488 9456 7540
rect 10692 7488 10744 7540
rect 8208 7420 8260 7472
rect 2044 7352 2096 7404
rect 2688 7352 2740 7404
rect 3516 7352 3568 7404
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 7012 7352 7064 7404
rect 6552 7284 6604 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 10232 7216 10284 7268
rect 14924 7216 14976 7268
rect 3148 7148 3200 7200
rect 3976 7148 4028 7200
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5816 7148 5868 7200
rect 7380 7148 7432 7200
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 1860 6944 1912 6996
rect 4252 6944 4304 6996
rect 7288 6944 7340 6996
rect 4160 6876 4212 6928
rect 3148 6808 3200 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 9404 6808 9456 6860
rect 2964 6740 3016 6792
rect 3240 6740 3292 6792
rect 3332 6672 3384 6724
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 6000 6740 6052 6792
rect 3976 6715 4028 6724
rect 3976 6681 3985 6715
rect 3985 6681 4019 6715
rect 4019 6681 4028 6715
rect 3976 6672 4028 6681
rect 4160 6672 4212 6724
rect 4896 6672 4948 6724
rect 5816 6672 5868 6724
rect 6644 6604 6696 6656
rect 7380 6740 7432 6792
rect 8484 6715 8536 6724
rect 8484 6681 8502 6715
rect 8502 6681 8536 6715
rect 8484 6672 8536 6681
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 9956 6740 10008 6792
rect 10416 6672 10468 6724
rect 7564 6604 7616 6656
rect 10048 6604 10100 6656
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 1860 6264 1912 6316
rect 1216 6196 1268 6248
rect 8484 6443 8536 6452
rect 8484 6409 8493 6443
rect 8493 6409 8527 6443
rect 8527 6409 8536 6443
rect 8484 6400 8536 6409
rect 9772 6400 9824 6452
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 7012 6264 7064 6316
rect 7656 6264 7708 6316
rect 8760 6264 8812 6316
rect 8852 6264 8904 6316
rect 10048 6332 10100 6384
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 10508 6400 10560 6452
rect 12164 6400 12216 6452
rect 14280 6400 14332 6452
rect 3516 6196 3568 6248
rect 3424 6128 3476 6180
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 9772 6128 9824 6180
rect 9956 6128 10008 6180
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 7564 6060 7616 6112
rect 8852 6060 8904 6112
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 14924 6196 14976 6248
rect 10784 6060 10836 6112
rect 12348 6060 12400 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 1492 5856 1544 5908
rect 2504 5856 2556 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 9312 5856 9364 5908
rect 10600 5856 10652 5908
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 7564 5652 7616 5704
rect 8208 5652 8260 5704
rect 6828 5584 6880 5636
rect 10784 5652 10836 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 6920 5516 6972 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 12164 5559 12216 5568
rect 12164 5525 12173 5559
rect 12173 5525 12207 5559
rect 12207 5525 12216 5559
rect 12164 5516 12216 5525
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 7196 5312 7248 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 7472 5176 7524 5228
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 6828 5108 6880 5160
rect 12440 5176 12492 5228
rect 7380 5040 7432 5092
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 6460 4768 6512 4820
rect 8208 4768 8260 4820
rect 8852 4768 8904 4820
rect 6920 4700 6972 4752
rect 14832 4700 14884 4752
rect 940 4564 992 4616
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 9220 4632 9272 4684
rect 8576 4609 8628 4616
rect 8576 4575 8585 4609
rect 8585 4575 8619 4609
rect 8619 4575 8628 4609
rect 8576 4564 8628 4575
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 12440 4496 12492 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 7288 4428 7340 4480
rect 14280 4428 14332 4480
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 1584 4020 1636 4072
rect 8576 4020 8628 4072
rect 9864 3884 9916 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 5448 3680 5500 3732
rect 14004 3680 14056 3732
rect 940 3476 992 3528
rect 5264 3476 5316 3528
rect 14556 3340 14608 3392
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 5264 3136 5316 3188
rect 9956 3136 10008 3188
rect 4160 3068 4212 3120
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 10324 3068 10376 3120
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 10140 3000 10192 3052
rect 13820 3068 13872 3120
rect 13912 3111 13964 3120
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 480 2796 532 2848
rect 4160 2839 4212 2848
rect 4160 2805 4169 2839
rect 4169 2805 4203 2839
rect 4203 2805 4212 2839
rect 4160 2796 4212 2805
rect 6000 2796 6052 2848
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 8392 2796 8444 2848
rect 8484 2796 8536 2848
rect 11152 2796 11204 2848
rect 12072 2839 12124 2848
rect 12072 2805 12081 2839
rect 12081 2805 12115 2839
rect 12115 2805 12124 2839
rect 12072 2796 12124 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 14464 2864 14516 2916
rect 13728 2796 13780 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 3056 2592 3108 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 1308 2320 1360 2372
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 3056 2363 3108 2372
rect 3056 2329 3065 2363
rect 3065 2329 3099 2363
rect 3099 2329 3108 2363
rect 3056 2320 3108 2329
rect 12164 2524 12216 2576
rect 6000 2456 6052 2508
rect 4160 2388 4212 2440
rect 4712 2388 4764 2440
rect 4988 2388 5040 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 6552 2388 6604 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 8484 2388 8536 2440
rect 9864 2388 9916 2440
rect 10232 2388 10284 2440
rect 11152 2388 11204 2440
rect 12072 2388 12124 2440
rect 12624 2388 12676 2440
rect 3884 2363 3936 2372
rect 3884 2329 3893 2363
rect 3893 2329 3927 2363
rect 3927 2329 3936 2363
rect 3884 2320 3936 2329
rect 6368 2363 6420 2372
rect 6368 2329 6377 2363
rect 6377 2329 6411 2363
rect 6411 2329 6420 2363
rect 6368 2320 6420 2329
rect 7196 2363 7248 2372
rect 7196 2329 7205 2363
rect 7205 2329 7239 2363
rect 7239 2329 7248 2363
rect 7196 2320 7248 2329
rect 4896 2295 4948 2304
rect 4896 2261 4905 2295
rect 4905 2261 4939 2295
rect 4939 2261 4948 2295
rect 4896 2252 4948 2261
rect 5540 2252 5592 2304
rect 8208 2252 8260 2304
rect 8760 2252 8812 2304
rect 9680 2252 9732 2304
rect 10416 2252 10468 2304
rect 11152 2252 11204 2304
rect 12256 2252 12308 2304
rect 12900 2252 12952 2304
rect 14556 2252 14608 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
<< metal2 >>
rect 938 19200 994 20000
rect 1674 19200 1730 20000
rect 2410 19200 2466 20000
rect 3146 19200 3202 20000
rect 3882 19200 3938 20000
rect 4618 19200 4674 20000
rect 5354 19200 5410 20000
rect 6090 19200 6146 20000
rect 6826 19200 6882 20000
rect 7562 19200 7618 20000
rect 8298 19200 8354 20000
rect 9034 19200 9090 20000
rect 9770 19200 9826 20000
rect 10506 19200 10562 20000
rect 11242 19200 11298 20000
rect 11978 19200 12034 20000
rect 12714 19200 12770 20000
rect 13450 19200 13506 20000
rect 14186 19200 14242 20000
rect 14922 19200 14978 20000
rect 952 17338 980 19200
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 940 17332 992 17338
rect 940 17274 992 17280
rect 1412 16590 1440 17983
rect 1688 17898 1716 19200
rect 1688 17870 1808 17898
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16794 1716 16934
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1780 16590 1808 17870
rect 2424 17338 2452 19200
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 3068 17270 3096 17546
rect 3160 17338 3188 19200
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 3252 17134 3280 17478
rect 3896 17184 3924 19200
rect 4632 17610 4660 19200
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 5368 17338 5396 19200
rect 6104 17338 6132 19200
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 3804 17156 3924 17184
rect 5724 17196 5776 17202
rect 3240 17128 3292 17134
rect 2976 17054 3096 17082
rect 3240 17070 3292 17076
rect 2976 16998 3004 17054
rect 1952 16992 2004 16998
rect 1872 16952 1952 16980
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16250 1808 16390
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 940 14408 992 14414
rect 940 14350 992 14356
rect 952 13977 980 14350
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 938 13968 994 13977
rect 938 13903 994 13912
rect 1596 13326 1624 14214
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 952 12617 980 13262
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 938 12608 994 12617
rect 938 12543 994 12552
rect 1596 12238 1624 13126
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 952 11257 980 11698
rect 1504 11354 1532 11698
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11354 1624 11494
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 938 11248 994 11257
rect 938 11183 994 11192
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 952 9897 980 9930
rect 938 9888 994 9897
rect 938 9823 994 9832
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8537 980 8842
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 1412 8090 1440 9522
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9178 1624 9318
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 8974 1716 15846
rect 1872 10742 1900 16952
rect 1952 16934 2004 16940
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 1950 16688 2006 16697
rect 1950 16623 2006 16632
rect 1964 16114 1992 16623
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1964 13190 1992 14010
rect 2056 13938 2084 16390
rect 2240 15094 2268 16934
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 3068 16794 3096 17054
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2872 16448 2924 16454
rect 2924 16396 3096 16402
rect 2872 16390 3096 16396
rect 2884 16374 3096 16390
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15706 2360 15982
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 3068 15586 3096 16374
rect 3160 15706 3188 16526
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3068 15558 3188 15586
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2976 14804 3004 15438
rect 3068 15162 3096 15438
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2976 14776 3096 14804
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12782 1992 13126
rect 2516 12986 2544 13670
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 3068 13326 3096 14776
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12986 2820 13126
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1964 10606 1992 12718
rect 2516 12306 2544 12922
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 10674 2452 12038
rect 2792 11898 2820 12174
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 3068 11218 3096 11494
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2516 10810 2544 11018
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 1964 9450 1992 10542
rect 2516 10266 2544 10542
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 3160 10062 3188 15558
rect 3252 15162 3280 16934
rect 3516 16584 3568 16590
rect 3436 16544 3516 16572
rect 3436 16454 3464 16544
rect 3516 16526 3568 16532
rect 3804 16522 3832 17156
rect 5724 17138 5776 17144
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16794 4108 17070
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 4540 16794 4568 16934
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3436 15570 3464 16186
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15570 3556 15846
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3344 15026 3372 15302
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 14074 3464 14350
rect 3620 14074 3648 14826
rect 3896 14260 3924 16594
rect 4172 15706 4200 16594
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4724 16182 4752 16934
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 15337 4108 15370
rect 4066 15328 4122 15337
rect 4066 15263 4122 15272
rect 4264 15144 4292 16118
rect 4724 15502 4752 16118
rect 4816 15706 4844 16526
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4344 15156 4396 15162
rect 4264 15116 4344 15144
rect 4344 15098 4396 15104
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4816 14890 4844 15030
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14278 4200 14758
rect 3712 14232 3924 14260
rect 4160 14272 4212 14278
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3620 13530 3648 13670
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3436 12434 3464 13262
rect 3436 12406 3556 12434
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11014 3280 12038
rect 3344 11762 3372 12174
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10810 3280 10950
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3344 10130 3372 11698
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10266 3464 10406
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 2148 8906 2176 9522
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9178 2268 9318
rect 2516 9178 2544 9454
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1398 7032 1454 7041
rect 1398 6967 1454 6976
rect 1216 6248 1268 6254
rect 1216 6190 1268 6196
rect 1228 5817 1256 6190
rect 1214 5808 1270 5817
rect 1214 5743 1270 5752
rect 1412 5710 1440 6967
rect 1504 5914 1532 8434
rect 1780 6458 1808 8434
rect 1964 7342 1992 8434
rect 2148 8022 2176 8842
rect 2240 8430 2268 9114
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2516 7546 2544 7754
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2700 7410 2728 7754
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1860 6996 1912 7002
rect 1964 6984 1992 7278
rect 1912 6956 1992 6984
rect 1860 6938 1912 6944
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1872 6322 1900 6938
rect 2056 6458 2084 7346
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 3068 6882 3096 7686
rect 3160 7206 3188 7822
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2976 6854 3096 6882
rect 3160 6866 3188 7142
rect 3148 6860 3200 6866
rect 2976 6798 3004 6854
rect 3148 6802 3200 6808
rect 3252 6798 3280 8298
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3344 6730 3372 8570
rect 3528 8514 3556 12406
rect 3620 12306 3648 13466
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3712 8634 3740 14232
rect 4160 14214 4212 14220
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12434 3832 13126
rect 3804 12406 4016 12434
rect 3988 12306 4016 12406
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 4080 12238 4108 13330
rect 4172 12850 4200 14214
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4816 14074 4844 14826
rect 4908 14396 4936 16458
rect 5000 16250 5028 16526
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4908 14368 5028 14396
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13326 4568 13670
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4816 13274 4844 13330
rect 4816 13246 4936 13274
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 4724 12918 4752 13126
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4632 12434 4660 12718
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12442 4752 12582
rect 4540 12406 4660 12434
rect 4712 12436 4764 12442
rect 4540 12374 4568 12406
rect 4712 12378 4764 12384
rect 4528 12368 4580 12374
rect 4724 12322 4752 12378
rect 4528 12310 4580 12316
rect 4632 12294 4752 12322
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4632 12084 4660 12294
rect 4712 12232 4764 12238
rect 4816 12220 4844 13126
rect 4908 12646 4936 13246
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4764 12192 4844 12220
rect 4908 12220 4936 12582
rect 5000 12322 5028 14368
rect 5092 12434 5120 16390
rect 5276 16182 5304 16934
rect 5736 16658 5764 17138
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5460 16114 5488 16390
rect 5736 16250 5764 16594
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5828 16182 5856 16934
rect 6012 16522 6040 16934
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15706 5488 16050
rect 6564 16046 6592 16458
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 15366 5488 15438
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5184 13938 5212 14758
rect 5276 14550 5304 14758
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5276 13462 5304 14350
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12782 5488 13262
rect 5552 12782 5580 15506
rect 6472 15434 6500 15846
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5828 14074 5856 14554
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5920 13938 5948 14486
rect 6012 14074 6040 14826
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 14074 6224 14214
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6472 13938 6500 15370
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6564 14074 6592 14962
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5092 12406 5212 12434
rect 5000 12294 5120 12322
rect 4988 12232 5040 12238
rect 4908 12192 4988 12220
rect 4712 12174 4764 12180
rect 4988 12174 5040 12180
rect 4632 12056 4752 12084
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3988 11150 4016 11562
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3896 8634 3924 9522
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3436 8486 3556 8514
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 3436 6186 3464 8486
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3528 8090 3556 8366
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3620 7970 3648 8366
rect 3528 7942 3648 7970
rect 3528 7750 3556 7942
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7410 3556 7686
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3528 6254 3556 7346
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6730 4016 7142
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2872 6112 2924 6118
rect 2924 6072 3096 6100
rect 2872 6054 2924 6060
rect 2516 5914 2544 6054
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4457 980 4558
rect 1584 4480 1636 4486
rect 938 4448 994 4457
rect 1584 4422 1636 4428
rect 938 4383 994 4392
rect 1596 4078 1624 4422
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 952 3097 980 3470
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 480 2848 532 2854
rect 480 2790 532 2796
rect 492 800 520 2790
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 3068 2650 3096 6072
rect 4080 3058 4108 11018
rect 4172 10606 4200 11222
rect 4264 10742 4292 11494
rect 4724 11082 4752 12056
rect 5092 11914 5120 12294
rect 4908 11886 5120 11914
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 9518 4200 10542
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 6934 4200 9454
rect 4448 9178 4476 9522
rect 4620 9376 4672 9382
rect 4672 9336 4752 9364
rect 4620 9318 4672 9324
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4632 8838 4660 9046
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4264 7002 4292 7822
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 3126 4200 6666
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 4172 2446 4200 2790
rect 4724 2446 4752 9336
rect 4816 8498 4844 9862
rect 4908 9042 4936 11886
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 11354 5028 11494
rect 5092 11354 5120 11698
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5184 11218 5212 12406
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5276 11744 5304 12174
rect 5356 11756 5408 11762
rect 5276 11716 5356 11744
rect 5356 11698 5408 11704
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10130 5212 11154
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5276 10062 5304 10950
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5368 9110 5396 11698
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5000 8634 5028 8774
rect 5184 8634 5212 8774
rect 5368 8634 5396 8910
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5092 7818 5120 8298
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 6798 4844 7686
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4908 6730 4936 7754
rect 5000 7546 5028 7754
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 5000 2446 5028 7142
rect 5460 3738 5488 12718
rect 5644 12714 5672 13738
rect 6012 13308 6040 13738
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6184 13320 6236 13326
rect 6012 13280 6184 13308
rect 6184 13262 6236 13268
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12850 6132 13126
rect 6196 12918 6224 13262
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12918 6316 13126
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6472 12850 6500 13262
rect 6092 12844 6144 12850
rect 6012 12804 6092 12832
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5644 12306 5672 12650
rect 6012 12442 6040 12804
rect 6092 12786 6144 12792
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10538 5580 11086
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5644 10266 5672 10950
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10266 5764 10406
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5828 7426 5856 12038
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5920 9722 5948 10610
rect 6380 10470 6408 10610
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6012 10266 6040 10406
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6472 10062 6500 11086
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6564 9586 6592 10474
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6460 8968 6512 8974
rect 6512 8928 6592 8956
rect 6460 8910 6512 8916
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6288 8634 6316 8774
rect 6472 8634 6500 8774
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6564 8498 6592 8928
rect 6656 8634 6684 17478
rect 6840 17134 6868 19200
rect 7576 17134 7604 19200
rect 8312 17814 8340 19200
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 7668 17338 7696 17750
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 9048 17338 9076 19200
rect 9784 17338 9812 19200
rect 10520 17338 10548 19200
rect 11256 17626 11284 19200
rect 11164 17598 11284 17626
rect 11164 17338 11192 17598
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 11992 17338 12020 19200
rect 12346 18048 12402 18057
rect 12346 17983 12402 17992
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 7756 17196 7808 17202
rect 7668 17156 7756 17184
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 12900 6776 16934
rect 7668 16590 7696 17156
rect 7756 17138 7808 17144
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7024 15502 7052 16390
rect 7576 15570 7604 16390
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14618 6868 14894
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6748 12872 6868 12900
rect 6840 10606 6868 12872
rect 6932 11830 6960 15302
rect 7116 14482 7144 15370
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14618 7236 14758
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12238 7052 13126
rect 7116 12918 7144 13194
rect 7208 12918 7236 13398
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7484 12730 7512 15438
rect 7668 15366 7696 16526
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 8312 16250 8340 16390
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8404 15502 8432 16934
rect 8496 16522 8524 16934
rect 9232 16794 9260 17138
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 8496 15706 8524 16458
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8864 15570 8892 16050
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7760 14618 7788 14962
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7852 14482 7880 14758
rect 8772 14618 8800 14758
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 9048 14482 9076 15982
rect 9140 15706 9168 16458
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16182 9812 16390
rect 9968 16250 9996 16458
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 7852 14260 7880 14418
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 7668 14232 7880 14260
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 13394 7604 13670
rect 7668 13394 7696 14232
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 8772 14074 8800 14350
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7760 13530 7788 13874
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 7484 12702 7696 12730
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 12306 7512 12582
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7576 12102 7604 12310
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 10198 6776 10474
rect 6828 10464 6880 10470
rect 6932 10452 6960 11086
rect 6880 10424 6960 10452
rect 6828 10406 6880 10412
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6840 9518 6868 10406
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5644 7398 5856 7426
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 3194 5304 3470
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5644 2446 5672 7398
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6730 5856 7142
rect 6012 6798 6040 7686
rect 6564 7342 6592 8434
rect 6656 7954 6684 8570
rect 6840 8514 6868 9114
rect 6932 8974 6960 9998
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9722 7144 9930
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7300 9450 7328 11086
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6840 8498 6960 8514
rect 6840 8492 6972 8498
rect 6840 8486 6920 8492
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6840 7886 6868 8486
rect 6920 8434 6972 8440
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 7954 6960 8298
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 6322 6684 6598
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6656 5710 6684 6258
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6840 5642 6868 7822
rect 7024 7410 7052 8842
rect 7392 8838 7420 11562
rect 7484 9654 7512 11630
rect 7576 10606 7604 12038
rect 7668 11626 7696 12702
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11218 7696 11562
rect 8220 11558 8248 12854
rect 8312 12306 8340 13330
rect 8864 13326 8892 14282
rect 9048 13938 9076 14418
rect 9324 14006 9352 15302
rect 10428 15026 10456 16050
rect 10612 15570 10640 16526
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 16250 10732 16458
rect 10796 16250 10824 16526
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10704 15706 10732 16050
rect 11072 16046 11100 16934
rect 11716 16794 11744 17206
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 11900 16794 11928 17138
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11164 16130 11192 16526
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 11164 16102 11284 16130
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14346 9444 14758
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 10060 14482 10088 14894
rect 10428 14618 10456 14962
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8772 12374 8800 13262
rect 9048 12986 9076 13874
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9876 13394 9904 14214
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10674 7696 10950
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7484 8786 7512 9454
rect 7576 8906 7604 10406
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7484 8758 7604 8786
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7116 6338 7144 7822
rect 7024 6322 7144 6338
rect 7012 6316 7144 6322
rect 7064 6310 7144 6316
rect 7012 6258 7064 6264
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 5166 6868 5578
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6472 4826 6500 5102
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6932 4758 6960 5510
rect 7208 5370 7236 8298
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 7002 7328 7278
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7392 6798 7420 7142
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7392 5098 7420 6734
rect 7484 5234 7512 7686
rect 7576 6662 7604 8758
rect 7668 8566 7696 8910
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 8220 7478 8248 11494
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5710 7604 6054
rect 7668 5914 7696 6258
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 8220 5370 8248 5646
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 8220 4826 8248 5306
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 7104 4616 7156 4622
rect 7156 4576 7328 4604
rect 7104 4558 7156 4564
rect 7300 4486 7328 4576
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 8312 3058 8340 12242
rect 9048 11898 9076 12922
rect 9324 12442 9352 13262
rect 9692 12986 9720 13262
rect 9680 12980 9732 12986
rect 9732 12940 9904 12968
rect 9680 12922 9732 12928
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11354 8524 11698
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8404 10674 8432 11290
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8680 10742 8708 11086
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 9692 10674 9720 11018
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 8496 10266 8524 10542
rect 9232 10266 9260 10542
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8498 8432 9318
rect 8588 9178 8616 9998
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8864 9586 8892 9930
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8864 8974 8892 9522
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 8090 8524 8230
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8864 7886 8892 8910
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 7954 9076 8774
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9140 7954 9168 8570
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8496 6458 8524 6666
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8772 6322 8800 6802
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8864 6118 8892 6258
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4826 8892 5102
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 9232 4690 9260 10066
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9324 9178 9352 9454
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 8498 9444 9522
rect 9680 9512 9732 9518
rect 9876 9500 9904 12940
rect 10060 12850 10088 14418
rect 10520 13530 10548 15438
rect 10704 15162 10732 15438
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 11072 15026 11100 15846
rect 11164 15706 11192 15982
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11256 15366 11284 16102
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 11624 15162 11652 15438
rect 11716 15434 11744 15846
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14414 11284 14758
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 11716 14074 11744 14826
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10428 12306 10456 13262
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12714 10548 13194
rect 10612 12986 10640 13262
rect 10704 13138 10732 13806
rect 11072 13394 11100 14010
rect 11716 13530 11744 14010
rect 11808 13870 11836 14350
rect 11900 14278 11928 14894
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14074 11928 14214
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 13394 11836 13806
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11888 13184 11940 13190
rect 10704 13110 10916 13138
rect 11888 13126 11940 13132
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10060 11898 10088 12242
rect 10520 12186 10548 12650
rect 10152 12158 10548 12186
rect 10784 12164 10836 12170
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9732 9472 9904 9500
rect 9680 9454 9732 9460
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 7546 9444 8434
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9876 8090 9904 8502
rect 9968 8430 9996 10406
rect 10060 10266 10088 10542
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10152 9874 10180 12158
rect 10784 12106 10836 12112
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10520 11762 10548 12038
rect 10704 11898 10732 12038
rect 10796 11898 10824 12106
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 10810 10272 11222
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10198 10272 10406
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10336 10062 10364 11562
rect 10888 11234 10916 13110
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11900 12850 11928 13126
rect 11992 12986 12020 16526
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11532 12434 11560 12718
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11532 12406 11652 12434
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10520 11206 10916 11234
rect 10520 11150 10548 11206
rect 10980 11150 11008 11562
rect 11072 11286 11100 12038
rect 11164 11286 11192 12174
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11520 11756 11572 11762
rect 11624 11744 11652 12406
rect 11716 12102 11744 12582
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11572 11716 11652 11744
rect 11520 11698 11572 11704
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10152 9846 10364 9874
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 9382 10180 9590
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10060 8566 10088 9318
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 7948 9916 7954
rect 9968 7936 9996 8230
rect 10060 8090 10088 8502
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9916 7908 9996 7936
rect 9864 7890 9916 7896
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9416 6866 9444 7482
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9784 6458 9812 6734
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9784 6186 9812 6394
rect 9968 6186 9996 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6390 10088 6598
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8588 4078 8616 4558
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 6012 2514 6040 2790
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6564 2446 6592 2790
rect 8404 2446 8432 2790
rect 8496 2446 8524 2790
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 9876 2446 9904 3878
rect 9968 3194 9996 6122
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10152 3058 10180 8298
rect 10244 7274 10272 8774
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10244 2446 10272 5510
rect 10336 3126 10364 9846
rect 10428 9586 10456 11018
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7886 10456 8230
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10520 6458 10548 11086
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10810 11100 11018
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 10266 10824 10542
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10266 11008 10406
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11624 10198 11652 11154
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 10266 11744 11018
rect 11900 10742 11928 12582
rect 11978 12336 12034 12345
rect 11978 12271 12034 12280
rect 11992 11354 12020 12271
rect 12084 11354 12112 17070
rect 12176 16250 12204 17138
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16250 12296 16390
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12360 16114 12388 17983
rect 12728 17338 12756 19200
rect 13464 17338 13492 19200
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 12636 16794 12664 17138
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 13280 16794 13308 17138
rect 13740 16794 13768 17138
rect 14200 16794 14228 19200
rect 14936 17898 14964 19200
rect 14936 17870 15056 17898
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 12532 16720 12584 16726
rect 13176 16720 13228 16726
rect 13174 16688 13176 16697
rect 13228 16688 13230 16697
rect 12584 16668 12664 16674
rect 12532 16662 12664 16668
rect 12544 16646 12664 16662
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 15162 12204 15438
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14278 12480 14758
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12544 13818 12572 16526
rect 12452 13790 12572 13818
rect 12452 12345 12480 13790
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 12850 12572 13670
rect 12532 12844 12584 12850
rect 12636 12832 12664 16646
rect 13174 16623 13230 16632
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 15706 12848 15982
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12728 14414 12756 14758
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12820 14074 12848 14758
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 13280 12866 13308 16458
rect 13556 16250 13584 16458
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13372 15706 13400 16050
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 15706 13492 15846
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13372 15162 13400 15642
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13372 14618 13400 14962
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13556 14618 13584 14894
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13648 14278 13676 16526
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 15434 13768 16390
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 15028 16250 15056 17870
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14646 15464 14702 15473
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 14568 15422 14646 15450
rect 13832 15162 13860 15370
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14200 15026 14228 15302
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14292 14618 14320 14962
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14568 14414 14596 15422
rect 14646 15399 14702 15408
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 13530 13676 14214
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14462 13968 14518 13977
rect 14462 13903 14464 13912
rect 14516 13903 14518 13912
rect 14464 13874 14516 13880
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 14200 13326 14228 13806
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 12820 12838 13308 12866
rect 13360 12844 13412 12850
rect 12636 12804 12756 12832
rect 12532 12786 12584 12792
rect 12438 12336 12494 12345
rect 12256 12300 12308 12306
rect 12438 12271 12494 12280
rect 12256 12242 12308 12248
rect 12268 11830 12296 12242
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11830 12388 12038
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11612 10192 11664 10198
rect 11664 10140 11744 10146
rect 11612 10134 11744 10140
rect 11624 10118 11744 10134
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 11624 9722 11652 9930
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 8974 11652 9318
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10612 8090 10640 8502
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10704 7886 10732 8774
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11716 8498 11744 10118
rect 11808 9518 11836 10542
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11808 8974 11836 9454
rect 11900 9450 11928 9862
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7546 10732 7822
rect 11624 7750 11652 8230
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10612 5914 10640 6190
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10796 5710 10824 6054
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 11888 3052 11940 3058
rect 11992 3040 12020 11290
rect 12452 10674 12480 11494
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8430 12204 8910
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12084 8090 12112 8366
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 6458 12204 8366
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5710 12388 6054
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 11940 3012 12020 3040
rect 11888 2994 11940 3000
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 11164 2446 11192 2790
rect 12084 2446 12112 2790
rect 12176 2582 12204 5510
rect 12452 5234 12480 9998
rect 12544 9738 12572 12786
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12238 12664 12582
rect 12728 12374 12756 12804
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12636 11354 12664 11698
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10742 12756 10950
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12544 9710 12664 9738
rect 12728 9722 12756 10678
rect 12820 10470 12848 12838
rect 13360 12786 13412 12792
rect 13084 12776 13136 12782
rect 13136 12724 13308 12730
rect 13084 12718 13308 12724
rect 13096 12702 13308 12718
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11762 13216 12310
rect 13280 11898 13308 12702
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 13280 11354 13308 11834
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13372 11150 13400 12786
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12306 13492 12582
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11354 13584 12038
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10810 13400 11086
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12636 9654 12664 9710
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12636 9058 12664 9590
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12820 9178 12848 9998
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 13280 9178 13308 9590
rect 13372 9382 13400 10746
rect 13648 10266 13676 12242
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11354 13768 12106
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 12636 9042 12848 9058
rect 12636 9036 12860 9042
rect 12636 9030 12808 9036
rect 12808 8978 12860 8984
rect 13372 8974 13400 9318
rect 13648 9178 13676 9998
rect 13740 9722 13768 9998
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12452 3058 12480 4490
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 13832 3126 13860 8298
rect 13924 3126 13952 10406
rect 14016 3738 14044 13194
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14108 12442 14136 12650
rect 14476 12617 14504 12718
rect 14462 12608 14518 12617
rect 14462 12543 14518 12552
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14462 11248 14518 11257
rect 14462 11183 14518 11192
rect 14476 10674 14504 11183
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14924 10056 14976 10062
rect 14922 10024 14924 10033
rect 14976 10024 14978 10033
rect 14922 9959 14978 9968
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9722 14320 9862
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 15028 8537 15056 8910
rect 15014 8528 15070 8537
rect 15014 8463 15070 8472
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 4622 14228 7686
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14280 7200 14332 7206
rect 14936 7177 14964 7210
rect 14280 7142 14332 7148
rect 14922 7168 14978 7177
rect 14292 6458 14320 7142
rect 14922 7103 14978 7112
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14936 5817 14964 6190
rect 14922 5808 14978 5817
rect 14922 5743 14978 5752
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14188 4616 14240 4622
rect 14844 4593 14872 4694
rect 14188 4558 14240 4564
rect 14830 4584 14886 4593
rect 14830 4519 14886 4528
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12636 2446 12664 2790
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4988 2440 5040 2446
rect 5632 2440 5684 2446
rect 4988 2382 5040 2388
rect 1308 2372 1360 2378
rect 2228 2372 2280 2378
rect 1308 2314 1360 2320
rect 2148 2332 2228 2360
rect 1320 800 1348 2314
rect 2148 800 2176 2332
rect 3056 2372 3108 2378
rect 2228 2314 2280 2320
rect 2976 2332 3056 2360
rect 2976 800 3004 2332
rect 3884 2372 3936 2378
rect 3056 2314 3108 2320
rect 3804 2332 3884 2360
rect 3804 800 3832 2332
rect 3884 2314 3936 2320
rect 5460 2366 5580 2394
rect 5632 2382 5684 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 9864 2440 9916 2446
rect 8484 2382 8536 2388
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 4632 870 4752 898
rect 4632 800 4660 870
rect 478 0 534 800
rect 1306 0 1362 800
rect 2134 0 2190 800
rect 2962 0 3018 800
rect 3790 0 3846 800
rect 4618 0 4674 800
rect 4724 762 4752 870
rect 4908 762 4936 2246
rect 5460 800 5488 2366
rect 5552 2310 5580 2366
rect 6368 2372 6420 2378
rect 6288 2332 6368 2360
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 6288 800 6316 2332
rect 6368 2314 6420 2320
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 9600 2366 9720 2394
rect 9864 2382 9916 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 7208 1170 7236 2314
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 7116 1142 7236 1170
rect 7116 800 7144 1142
rect 7944 870 8064 898
rect 7944 800 7972 870
rect 4724 734 4936 762
rect 5446 0 5502 800
rect 6274 0 6330 800
rect 7102 0 7158 800
rect 7930 0 7986 800
rect 8036 762 8064 870
rect 8220 762 8248 2246
rect 8772 800 8800 2246
rect 9600 800 9628 2366
rect 9692 2310 9720 2366
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 10428 800 10456 2246
rect 11164 1170 11192 2246
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 12268 1170 12296 2246
rect 11164 1142 11284 1170
rect 11256 800 11284 1142
rect 12084 1142 12296 1170
rect 12084 800 12112 1142
rect 12912 800 12940 2246
rect 13740 800 13768 2790
rect 14292 2650 14320 4422
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 3074 14596 3334
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14646 3088 14702 3097
rect 14568 3046 14646 3074
rect 14646 3023 14702 3032
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14476 1442 14504 2858
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14568 1714 14596 2246
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 14646 1728 14702 1737
rect 14568 1686 14646 1714
rect 14646 1663 14702 1672
rect 14476 1414 14596 1442
rect 14568 800 14596 1414
rect 8036 734 8248 762
rect 8758 0 8814 800
rect 9586 0 9642 800
rect 10414 0 10470 800
rect 11242 0 11298 800
rect 12070 0 12126 800
rect 12898 0 12954 800
rect 13726 0 13782 800
rect 14554 0 14610 800
<< via2 >>
rect 1398 17992 1454 18048
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 938 13912 994 13968
rect 938 12552 994 12608
rect 938 11192 994 11248
rect 938 9832 994 9888
rect 938 8472 994 8528
rect 1950 16632 2006 16688
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4066 15272 4122 15328
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 1398 6976 1454 7032
rect 1214 5752 1270 5808
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 938 4392 994 4448
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 938 3032 994 3088
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 12346 17992 12402 18048
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11978 12280 12034 12336
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 13174 16668 13176 16688
rect 13176 16668 13228 16688
rect 13228 16668 13230 16688
rect 13174 16632 13230 16668
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14646 15408 14702 15464
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14462 13932 14518 13968
rect 14462 13912 14464 13932
rect 14464 13912 14516 13932
rect 14516 13912 14518 13932
rect 12438 12280 12494 12336
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14462 12552 14518 12608
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14462 11192 14518 11248
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14922 10004 14924 10024
rect 14924 10004 14976 10024
rect 14976 10004 14978 10024
rect 14922 9968 14978 10004
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 15014 8472 15070 8528
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14922 7112 14978 7168
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14922 5752 14978 5808
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14830 4528 14886 4584
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 14646 3032 14702 3088
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 14646 1672 14702 1728
<< metal3 >>
rect 0 18050 800 18080
rect 1393 18050 1459 18053
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 0 17960 800 17990
rect 1393 17987 1459 17990
rect 12341 18050 12407 18053
rect 15200 18050 16000 18080
rect 12341 18048 16000 18050
rect 12341 17992 12346 18048
rect 12402 17992 16000 18048
rect 12341 17990 16000 17992
rect 12341 17987 12407 17990
rect 15200 17960 16000 17990
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 12940 16831 13256 16832
rect 0 16690 800 16720
rect 1945 16690 2011 16693
rect 0 16688 2011 16690
rect 0 16632 1950 16688
rect 2006 16632 2011 16688
rect 0 16630 2011 16632
rect 0 16600 800 16630
rect 1945 16627 2011 16630
rect 13169 16690 13235 16693
rect 15200 16690 16000 16720
rect 13169 16688 16000 16690
rect 13169 16632 13174 16688
rect 13230 16632 16000 16688
rect 13169 16630 16000 16632
rect 13169 16627 13235 16630
rect 15200 16600 16000 16630
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 14641 15466 14707 15469
rect 14641 15464 15210 15466
rect 14641 15408 14646 15464
rect 14702 15408 15210 15464
rect 14641 15406 15210 15408
rect 14641 15403 14707 15406
rect 15150 15360 15210 15406
rect 0 15330 800 15360
rect 4061 15330 4127 15333
rect 0 15328 4127 15330
rect 0 15272 4066 15328
rect 4122 15272 4127 15328
rect 0 15270 4127 15272
rect 15150 15270 16000 15360
rect 0 15240 800 15270
rect 4061 15267 4127 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 15200 15240 16000 15270
rect 14653 15199 14969 15200
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 0 13970 800 14000
rect 933 13970 999 13973
rect 0 13968 999 13970
rect 0 13912 938 13968
rect 994 13912 999 13968
rect 0 13910 999 13912
rect 0 13880 800 13910
rect 933 13907 999 13910
rect 14457 13970 14523 13973
rect 15200 13970 16000 14000
rect 14457 13968 16000 13970
rect 14457 13912 14462 13968
rect 14518 13912 16000 13968
rect 14457 13910 16000 13912
rect 14457 13907 14523 13910
rect 15200 13880 16000 13910
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 0 12610 800 12640
rect 933 12610 999 12613
rect 0 12608 999 12610
rect 0 12552 938 12608
rect 994 12552 999 12608
rect 0 12550 999 12552
rect 0 12520 800 12550
rect 933 12547 999 12550
rect 14457 12610 14523 12613
rect 15200 12610 16000 12640
rect 14457 12608 16000 12610
rect 14457 12552 14462 12608
rect 14518 12552 16000 12608
rect 14457 12550 16000 12552
rect 14457 12547 14523 12550
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 15200 12520 16000 12550
rect 12940 12479 13256 12480
rect 11973 12338 12039 12341
rect 12433 12338 12499 12341
rect 11973 12336 12499 12338
rect 11973 12280 11978 12336
rect 12034 12280 12438 12336
rect 12494 12280 12499 12336
rect 11973 12278 12499 12280
rect 11973 12275 12039 12278
rect 12433 12275 12499 12278
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 14653 11935 14969 11936
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 0 11250 800 11280
rect 933 11250 999 11253
rect 0 11248 999 11250
rect 0 11192 938 11248
rect 994 11192 999 11248
rect 0 11190 999 11192
rect 0 11160 800 11190
rect 933 11187 999 11190
rect 14457 11250 14523 11253
rect 15200 11250 16000 11280
rect 14457 11248 16000 11250
rect 14457 11192 14462 11248
rect 14518 11192 16000 11248
rect 14457 11190 16000 11192
rect 14457 11187 14523 11190
rect 15200 11160 16000 11190
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 14917 10026 14983 10029
rect 14917 10024 15210 10026
rect 14917 9968 14922 10024
rect 14978 9968 15210 10024
rect 14917 9966 15210 9968
rect 14917 9963 14983 9966
rect 15150 9920 15210 9966
rect 0 9890 800 9920
rect 933 9890 999 9893
rect 0 9888 999 9890
rect 0 9832 938 9888
rect 994 9832 999 9888
rect 0 9830 999 9832
rect 15150 9830 16000 9920
rect 0 9800 800 9830
rect 933 9827 999 9830
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 15200 9800 16000 9830
rect 14653 9759 14969 9760
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 15009 8530 15075 8533
rect 15200 8530 16000 8560
rect 15009 8528 16000 8530
rect 15009 8472 15014 8528
rect 15070 8472 16000 8528
rect 15009 8470 16000 8472
rect 15009 8467 15075 8470
rect 15200 8440 16000 8470
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 0 7170 800 7200
rect 14917 7170 14983 7173
rect 15200 7170 16000 7200
rect 0 7080 858 7170
rect 14917 7168 16000 7170
rect 14917 7112 14922 7168
rect 14978 7112 16000 7168
rect 14917 7110 16000 7112
rect 14917 7107 14983 7110
rect 798 7034 858 7080
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 15200 7080 16000 7110
rect 12940 7039 13256 7040
rect 1393 7034 1459 7037
rect 798 7032 1459 7034
rect 798 6976 1398 7032
rect 1454 6976 1459 7032
rect 798 6974 1459 6976
rect 1393 6971 1459 6974
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 0 5810 800 5840
rect 1209 5810 1275 5813
rect 0 5808 1275 5810
rect 0 5752 1214 5808
rect 1270 5752 1275 5808
rect 0 5750 1275 5752
rect 0 5720 800 5750
rect 1209 5747 1275 5750
rect 14917 5810 14983 5813
rect 15200 5810 16000 5840
rect 14917 5808 16000 5810
rect 14917 5752 14922 5808
rect 14978 5752 16000 5808
rect 14917 5750 16000 5752
rect 14917 5747 14983 5750
rect 15200 5720 16000 5750
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 14825 4586 14891 4589
rect 14825 4584 15210 4586
rect 14825 4528 14830 4584
rect 14886 4528 15210 4584
rect 14825 4526 15210 4528
rect 14825 4523 14891 4526
rect 15150 4480 15210 4526
rect 0 4450 800 4480
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 0 4390 999 4392
rect 15150 4390 16000 4480
rect 0 4360 800 4390
rect 933 4387 999 4390
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 15200 4360 16000 4390
rect 14653 4319 14969 4320
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 14641 3090 14707 3093
rect 15200 3090 16000 3120
rect 14641 3088 16000 3090
rect 14641 3032 14646 3088
rect 14702 3032 16000 3088
rect 14641 3030 16000 3032
rect 14641 3027 14707 3030
rect 15200 3000 16000 3030
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 14641 1730 14707 1733
rect 15200 1730 16000 1760
rect 14641 1728 16000 1730
rect 14641 1672 14646 1728
rect 14702 1672 16000 1728
rect 14641 1670 16000 1672
rect 14641 1667 14707 1670
rect 15200 1640 16000 1670
<< via3 >>
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 16896 2977 17456
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 17440 4690 17456
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 16896 6404 17456
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 17440 8117 17456
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 16896 9831 17456
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 17440 11544 17456
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 16896 13258 17456
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 17440 14971 17456
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__inv_2  _161_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform -1 0 3680 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1688980957
transform 1 0 4324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1688980957
transform -1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform -1 0 2668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1688980957
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1688980957
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1688980957
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1688980957
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1688980957
transform -1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1688980957
transform -1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1688980957
transform -1 0 5336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1688980957
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1688980957
transform -1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1688980957
transform -1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1688980957
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1688980957
transform -1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1688980957
transform -1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1688980957
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1688980957
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1688980957
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1688980957
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1688980957
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1688980957
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1688980957
transform -1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1688980957
transform -1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1688980957
transform -1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1688980957
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1688980957
transform 1 0 7452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1688980957
transform -1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform -1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1688980957
transform -1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1688980957
transform -1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1688980957
transform -1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1688980957
transform -1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1688980957
transform -1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1688980957
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1688980957
transform -1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform 1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1688980957
transform -1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1688980957
transform 1 0 7820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1688980957
transform -1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1688980957
transform 1 0 6440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1688980957
transform 1 0 8280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform -1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1688980957
transform -1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1688980957
transform -1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1688980957
transform -1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1688980957
transform -1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1688980957
transform 1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1688980957
transform -1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1688980957
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1688980957
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1688980957
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1688980957
transform -1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1688980957
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform -1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform -1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1688980957
transform -1 0 12052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform -1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1688980957
transform -1 0 10580 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1688980957
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1688980957
transform -1 0 10212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1688980957
transform -1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1688980957
transform -1 0 10672 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1688980957
transform -1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1688980957
transform -1 0 7636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1688980957
transform -1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1688980957
transform -1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1688980957
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1688980957
transform -1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1688980957
transform -1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1688980957
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1688980957
transform 1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1688980957
transform 1 0 5244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1688980957
transform -1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1688980957
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1688980957
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _273_
timestamp 1688980957
transform -1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1688980957
transform -1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1688980957
transform -1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1688980957
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1688980957
transform -1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1688980957
transform -1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1688980957
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1688980957
transform -1 0 10580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1688980957
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1688980957
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1688980957
transform -1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1688980957
transform 1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1688980957
transform -1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1688980957
transform -1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1688980957
transform 1 0 3036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1688980957
transform -1 0 3036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1688980957
transform -1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1688980957
transform -1 0 5520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1688980957
transform -1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1688980957
transform -1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1688980957
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1688980957
transform -1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1688980957
transform 1 0 14260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1688980957
transform 1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1688980957
transform 1 0 1472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1688980957
transform -1 0 10488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1688980957
transform -1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1688980957
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1688980957
transform 1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1688980957
transform 1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1688980957
transform -1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1688980957
transform 1 0 11592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1688980957
transform -1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1688980957
transform 1 0 11592 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1688980957
transform 1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1688980957
transform -1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1688980957
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1688980957
transform 1 0 1564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1688980957
transform -1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform -1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1688980957
transform 1 0 5244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1688980957
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform -1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1688980957
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1688980957
transform -1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1688980957
transform -1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1688980957
transform -1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1688980957
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1688980957
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform -1 0 2944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1688980957
transform 1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1688980957
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1688980957
transform -1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1688980957
transform -1 0 4324 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _357_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 1688980957
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _359_
timestamp 1688980957
transform 1 0 8740 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _360_
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _361_
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _362_
timestamp 1688980957
transform 1 0 6808 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _364_
timestamp 1688980957
transform -1 0 8740 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1688980957
transform 1 0 6256 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1688980957
transform 1 0 9016 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1688980957
transform -1 0 9660 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1688980957
transform -1 0 11960 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1688980957
transform 1 0 11776 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1688980957
transform 1 0 11776 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _375_
timestamp 1688980957
transform -1 0 12328 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1688980957
transform 1 0 6900 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _378_
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1688980957
transform 1 0 2116 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1688980957
transform -1 0 2852 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _381_
timestamp 1688980957
transform -1 0 11960 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1688980957
transform 1 0 2760 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1688980957
transform -1 0 2852 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _384_
timestamp 1688980957
transform -1 0 4232 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1688980957
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1688980957
transform -1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1688980957
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _401_
timestamp 1688980957
transform -1 0 12420 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1688980957
transform -1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1688980957
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1688980957
transform -1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1688980957
transform -1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1688980957
transform -1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1688980957
transform -1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1688980957
transform -1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1688980957
transform -1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _412_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _412__63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _413_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _414_
timestamp 1688980957
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _415_
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _416_
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _417_
timestamp 1688980957
transform 1 0 3864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _418_
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _419_
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _420_
timestamp 1688980957
transform -1 0 13984 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _421_
timestamp 1688980957
transform 1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _422_
timestamp 1688980957
transform 1 0 11224 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _423__64
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _423_
timestamp 1688980957
transform -1 0 11316 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _424_
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _425_
timestamp 1688980957
transform -1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _426_
timestamp 1688980957
transform 1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _427_
timestamp 1688980957
transform 1 0 11040 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _428_
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _429_
timestamp 1688980957
transform 1 0 9844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _430_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _431_
timestamp 1688980957
transform 1 0 6072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _432_
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _433__65
timestamp 1688980957
transform 1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _433_
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _434_
timestamp 1688980957
transform 1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _435_
timestamp 1688980957
transform 1 0 7544 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _436_
timestamp 1688980957
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _437_
timestamp 1688980957
transform 1 0 9568 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _438_
timestamp 1688980957
transform -1 0 9752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _439_
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _440_
timestamp 1688980957
transform 1 0 6808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _441_
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _442_
timestamp 1688980957
transform 1 0 9752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _443_
timestamp 1688980957
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _443__66
timestamp 1688980957
transform -1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _444_
timestamp 1688980957
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _445_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _446_
timestamp 1688980957
transform -1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _447_
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _448__67
timestamp 1688980957
transform -1 0 11224 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _448_
timestamp 1688980957
transform 1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _449_
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _450_
timestamp 1688980957
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _451_
timestamp 1688980957
transform 1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _452__68
timestamp 1688980957
transform 1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _452_
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _453_
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _454_
timestamp 1688980957
transform 1 0 12788 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _455_
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _456_
timestamp 1688980957
transform -1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _457__69
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _457_
timestamp 1688980957
transform -1 0 11408 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _458_
timestamp 1688980957
transform 1 0 12420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _459_
timestamp 1688980957
transform -1 0 13984 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _460_
timestamp 1688980957
transform -1 0 13984 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _461_
timestamp 1688980957
transform 1 0 12328 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _462_
timestamp 1688980957
transform -1 0 13892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _463_
timestamp 1688980957
transform 1 0 12328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _464_
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _465_
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _465__70
timestamp 1688980957
transform -1 0 6992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _466_
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _467_
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _468_
timestamp 1688980957
transform -1 0 9476 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _469_
timestamp 1688980957
transform 1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _470_
timestamp 1688980957
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _471_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _472_
timestamp 1688980957
transform 1 0 6808 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _473_
timestamp 1688980957
transform 1 0 5336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _474_
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _475_
timestamp 1688980957
transform 1 0 5152 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _476_
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _477__71
timestamp 1688980957
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _477_
timestamp 1688980957
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _478_
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _479_
timestamp 1688980957
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _480_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _481_
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _482_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _483_
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _484_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _485_
timestamp 1688980957
transform -1 0 8924 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _486_
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _487_
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _488_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _489__72
timestamp 1688980957
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _489_
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _490_
timestamp 1688980957
transform -1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _491_
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _492_
timestamp 1688980957
transform -1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _493_
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _494_
timestamp 1688980957
transform -1 0 5244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _495_
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _496_
timestamp 1688980957
transform -1 0 3772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _497_
timestamp 1688980957
transform -1 0 2668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _498_
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _499_
timestamp 1688980957
transform -1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _500_
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _501__73
timestamp 1688980957
transform -1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _501_
timestamp 1688980957
transform 1 0 2576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _502_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _503_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _504_
timestamp 1688980957
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _505_
timestamp 1688980957
transform -1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _506_
timestamp 1688980957
transform -1 0 4876 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _507_
timestamp 1688980957
transform 1 0 2576 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _508_
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _509_
timestamp 1688980957
transform 1 0 1840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _510_
timestamp 1688980957
transform -1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _511_
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_18
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_36
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_91
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_43
timestamp 1688980957
transform 1 0 5060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_79
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_87
timestamp 1688980957
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_120
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_126
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 1688980957
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 1688980957
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1688980957
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_47
timestamp 1688980957
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_59
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_71
timestamp 1688980957
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_88
timestamp 1688980957
transform 1 0 9200 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_100
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_61
timestamp 1688980957
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_80
timestamp 1688980957
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_47
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_74
timestamp 1688980957
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_88
timestamp 1688980957
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_100
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1688980957
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1688980957
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_63
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_75
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_100
timestamp 1688980957
transform 1 0 10304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_112
timestamp 1688980957
transform 1 0 11408 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_145
timestamp 1688980957
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_8
timestamp 1688980957
transform 1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_22
timestamp 1688980957
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_34
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_46
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_79
timestamp 1688980957
transform 1 0 8372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_120
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_132
timestamp 1688980957
transform 1 0 13248 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_140
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1688980957
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_41
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_72
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_103
timestamp 1688980957
transform 1 0 10580 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_115
timestamp 1688980957
transform 1 0 11684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_127
timestamp 1688980957
transform 1 0 12788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_122
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_134
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_144
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_17
timestamp 1688980957
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_60
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_95
timestamp 1688980957
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_118
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_144
timestamp 1688980957
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_34
timestamp 1688980957
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_47
timestamp 1688980957
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_68
timestamp 1688980957
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_130
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_7
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_22
timestamp 1688980957
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_78
timestamp 1688980957
transform 1 0 8280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_88
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_96
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_106
timestamp 1688980957
transform 1 0 10856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1688980957
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_94
timestamp 1688980957
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_135
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_44
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_144
timestamp 1688980957
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_6
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_34
timestamp 1688980957
transform 1 0 4232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_46
timestamp 1688980957
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_132
timestamp 1688980957
transform 1 0 13248 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_8
timestamp 1688980957
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_24
timestamp 1688980957
transform 1 0 3312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_56
timestamp 1688980957
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_91
timestamp 1688980957
transform 1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_130
timestamp 1688980957
transform 1 0 13064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_144
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_102
timestamp 1688980957
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_116
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_44
timestamp 1688980957
transform 1 0 5152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_54
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_117
timestamp 1688980957
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1688980957
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_17
timestamp 1688980957
transform 1 0 2668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_38
timestamp 1688980957
transform 1 0 4600 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_52
timestamp 1688980957
transform 1 0 5888 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_76
timestamp 1688980957
transform 1 0 8096 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_97
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_132
timestamp 1688980957
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_6
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_18
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_24
timestamp 1688980957
transform 1 0 3312 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_38
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_36
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_47
timestamp 1688980957
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_70
timestamp 1688980957
transform 1 0 7544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_99
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_35
timestamp 1688980957
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_44
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_72
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_118
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_144
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_66
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_83
timestamp 1688980957
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_87
timestamp 1688980957
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_91
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_117
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_130
timestamp 1688980957
transform 1 0 13064 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_138
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_38
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_129
timestamp 1688980957
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_144
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_29
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_46
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_101
timestamp 1688980957
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_144
timestamp 1688980957
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 9200 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 14260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 10212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 4508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 7636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 13340 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 1840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 7728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 2024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 9016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform -1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1688980957
transform -1 0 14536 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1688980957
transform -1 0 14536 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 13432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform -1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform -1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform -1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform -1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output36 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform -1 0 2760 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 3588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 4416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform -1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform -1 0 8556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output49
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output53
timestamp 1688980957
transform -1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform -1 0 10396 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1688980957
transform -1 0 11132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output57
timestamp 1688980957
transform -1 0 12052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 12788 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 13984 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal3 s 15200 3000 16000 3120 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 15200 4360 16000 4480 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 3 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 4 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 5 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 6 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 7 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 8 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 9 nsew signal input
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 10 nsew signal input
flabel metal2 s 478 0 534 800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 11 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 12 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 13 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 14 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 15 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 16 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 17 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 18 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 19 nsew signal tristate
flabel metal3 s 15200 5720 16000 5840 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 20 nsew signal input
flabel metal3 s 15200 7080 16000 7200 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 21 nsew signal input
flabel metal3 s 15200 8440 16000 8560 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 22 nsew signal input
flabel metal3 s 15200 9800 16000 9920 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 23 nsew signal input
flabel metal3 s 15200 11160 16000 11280 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 24 nsew signal input
flabel metal3 s 15200 12520 16000 12640 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 25 nsew signal input
flabel metal3 s 15200 13880 16000 14000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 26 nsew signal input
flabel metal3 s 15200 15240 16000 15360 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 27 nsew signal input
flabel metal3 s 15200 16600 16000 16720 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 28 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 29 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 30 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 31 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 32 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 33 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 34 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 35 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 36 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 37 nsew signal tristate
flabel metal2 s 1674 19200 1730 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 38 nsew signal input
flabel metal2 s 2410 19200 2466 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 39 nsew signal input
flabel metal2 s 3146 19200 3202 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 40 nsew signal input
flabel metal2 s 3882 19200 3938 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 41 nsew signal input
flabel metal2 s 4618 19200 4674 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 42 nsew signal input
flabel metal2 s 5354 19200 5410 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 43 nsew signal input
flabel metal2 s 6090 19200 6146 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 44 nsew signal input
flabel metal2 s 6826 19200 6882 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 45 nsew signal input
flabel metal2 s 7562 19200 7618 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 46 nsew signal input
flabel metal2 s 9034 19200 9090 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 47 nsew signal tristate
flabel metal2 s 9770 19200 9826 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 48 nsew signal tristate
flabel metal2 s 10506 19200 10562 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 49 nsew signal tristate
flabel metal2 s 11242 19200 11298 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 50 nsew signal tristate
flabel metal2 s 11978 19200 12034 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 51 nsew signal tristate
flabel metal2 s 12714 19200 12770 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 52 nsew signal tristate
flabel metal2 s 13450 19200 13506 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 53 nsew signal tristate
flabel metal2 s 14186 19200 14242 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 54 nsew signal tristate
flabel metal2 s 14922 19200 14978 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 55 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 56 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 57 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 prog_clk
port 58 nsew signal input
flabel metal3 s 15200 1640 16000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 59 nsew signal input
flabel metal3 s 15200 17960 16000 18080 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 60 nsew signal input
flabel metal2 s 938 19200 994 20000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 61 nsew signal input
flabel metal2 s 8298 19200 8354 20000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 62 nsew signal input
flabel metal4 s 2657 2128 2977 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 6084 2128 6404 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 9511 2128 9831 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 12938 2128 13258 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 4370 2128 4690 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
rlabel metal1 7958 16864 7958 16864 0 vdd
rlabel via1 8037 17408 8037 17408 0 vss
rlabel metal1 3358 14042 3358 14042 0 _000_
rlabel metal1 4002 13226 4002 13226 0 _001_
rlabel metal1 2392 13294 2392 13294 0 _002_
rlabel metal2 4002 11356 4002 11356 0 _003_
rlabel metal1 1564 13906 1564 13906 0 _004_
rlabel metal1 2484 10030 2484 10030 0 _005_
rlabel metal1 4048 8942 4048 8942 0 _006_
rlabel metal1 4462 6970 4462 6970 0 _007_
rlabel metal1 11408 7854 11408 7854 0 _008_
rlabel metal1 1840 7378 1840 7378 0 _009_
rlabel metal1 1518 8058 1518 8058 0 _010_
rlabel metal2 1794 7446 1794 7446 0 _011_
rlabel metal1 5428 8602 5428 8602 0 _012_
rlabel metal1 6578 6188 6578 6188 0 _013_
rlabel metal1 5980 5202 5980 5202 0 _014_
rlabel metal1 10258 6324 10258 6324 0 _015_
rlabel metal1 7222 4624 7222 4624 0 _016_
rlabel metal1 7774 5712 7774 5712 0 _017_
rlabel metal1 4968 14382 4968 14382 0 _018_
rlabel metal1 7222 14042 7222 14042 0 _019_
rlabel metal1 8050 14586 8050 14586 0 _020_
rlabel metal1 9292 12206 9292 12206 0 _021_
rlabel metal2 4784 12206 4784 12206 0 _022_
rlabel metal1 6348 12682 6348 12682 0 _023_
rlabel metal1 13616 9554 13616 9554 0 _024_
rlabel metal1 13018 8942 13018 8942 0 _025_
rlabel metal1 14352 11322 14352 11322 0 _026_
rlabel metal2 13570 11696 13570 11696 0 _027_
rlabel metal1 10396 13906 10396 13906 0 _028_
rlabel metal1 12098 15130 12098 15130 0 _029_
rlabel metal1 10212 12818 10212 12818 0 _030_
rlabel metal1 11408 14994 11408 14994 0 _031_
rlabel metal1 7456 16558 7456 16558 0 _032_
rlabel metal1 9154 16082 9154 16082 0 _033_
rlabel metal1 10442 15674 10442 15674 0 _034_
rlabel metal1 5198 10030 5198 10030 0 _035_
rlabel metal1 8556 9146 8556 9146 0 _036_
rlabel metal2 7314 10268 7314 10268 0 _037_
rlabel metal1 10178 7854 10178 7854 0 _038_
rlabel metal2 8510 8160 8510 8160 0 _039_
rlabel metal2 5934 10166 5934 10166 0 _040_
rlabel metal1 10580 10030 10580 10030 0 _041_
rlabel metal1 10994 10642 10994 10642 0 _042_
rlabel metal1 12236 10030 12236 10030 0 _043_
rlabel metal1 11178 11866 11178 11866 0 _044_
rlabel metal1 2944 14994 2944 14994 0 _045_
rlabel metal1 5198 15470 5198 15470 0 _046_
rlabel metal1 4462 13294 4462 13294 0 _047_
rlabel metal1 6210 17136 6210 17136 0 _048_
rlabel metal1 3910 15606 3910 15606 0 _049_
rlabel metal1 3726 16762 3726 16762 0 _050_
rlabel metal1 5888 16490 5888 16490 0 _051_
rlabel metal1 5612 15470 5612 15470 0 _052_
rlabel metal1 3036 15130 3036 15130 0 _053_
rlabel metal1 5060 12886 5060 12886 0 _054_
rlabel metal2 4186 16150 4186 16150 0 _055_
rlabel metal1 6210 16150 6210 16150 0 _056_
rlabel metal1 2530 15674 2530 15674 0 _057_
rlabel metal2 13754 15912 13754 15912 0 _058_
rlabel metal1 4738 16218 4738 16218 0 _059_
rlabel metal1 11960 10234 11960 10234 0 _060_
rlabel metal1 10810 11730 10810 11730 0 _061_
rlabel metal2 10810 10404 10810 10404 0 _062_
rlabel metal1 11316 10778 11316 10778 0 _063_
rlabel metal1 5658 10098 5658 10098 0 _064_
rlabel metal1 12006 9690 12006 9690 0 _065_
rlabel metal1 11684 11254 11684 11254 0 _066_
rlabel metal1 10120 10234 10120 10234 0 _067_
rlabel metal1 8786 11186 8786 11186 0 _068_
rlabel metal1 6164 10098 6164 10098 0 _069_
rlabel metal1 10442 8058 10442 8058 0 _070_
rlabel metal1 9200 7922 9200 7922 0 _071_
rlabel metal1 8464 10234 8464 10234 0 _072_
rlabel metal1 7636 11118 7636 11118 0 _073_
rlabel metal1 5474 10234 5474 10234 0 _074_
rlabel metal2 9890 8296 9890 8296 0 _075_
rlabel metal1 9384 9146 9384 9146 0 _076_
rlabel metal1 9154 10234 9154 10234 0 _077_
rlabel metal1 6854 10642 6854 10642 0 _078_
rlabel metal1 6486 11186 6486 11186 0 _079_
rlabel metal1 9706 16218 9706 16218 0 _080_
rlabel metal1 10856 16218 10856 16218 0 _081_
rlabel metal1 7820 15538 7820 15538 0 _082_
rlabel metal1 9476 15674 9476 15674 0 _083_
rlabel metal1 10166 16116 10166 16116 0 _084_
rlabel metal1 8234 17204 8234 17204 0 _085_
rlabel metal1 11592 15130 11592 15130 0 _086_
rlabel metal1 10534 12954 10534 12954 0 _087_
rlabel metal1 10580 15130 10580 15130 0 _088_
rlabel metal2 9890 13804 9890 13804 0 _089_
rlabel metal1 12374 15572 12374 15572 0 _090_
rlabel metal1 11224 13362 11224 13362 0 _091_
rlabel metal2 13570 14756 13570 14756 0 _092_
rlabel metal1 11270 13838 11270 13838 0 _093_
rlabel metal1 14030 11832 14030 11832 0 _094_
rlabel metal2 14122 12546 14122 12546 0 _095_
rlabel metal1 12972 9146 12972 9146 0 _096_
rlabel metal1 13754 9452 13754 9452 0 _097_
rlabel metal1 13984 11254 13984 11254 0 _098_
rlabel metal1 13018 12274 13018 12274 0 _099_
rlabel metal1 13570 9146 13570 9146 0 _100_
rlabel metal1 12558 8908 12558 8908 0 _101_
rlabel metal1 8050 12104 8050 12104 0 _102_
rlabel metal1 7314 12852 7314 12852 0 _103_
rlabel metal1 7452 14450 7452 14450 0 _104_
rlabel metal1 5750 12172 5750 12172 0 _105_
rlabel metal1 9246 14892 9246 14892 0 _106_
rlabel metal1 5566 14518 5566 14518 0 _107_
rlabel metal1 8326 13226 8326 13226 0 _108_
rlabel metal1 6578 12852 6578 12852 0 _109_
rlabel metal1 6072 14042 6072 14042 0 _110_
rlabel metal1 5290 13362 5290 13362 0 _111_
rlabel metal1 6762 14450 6762 14450 0 _112_
rlabel metal1 5382 13940 5382 13940 0 _113_
rlabel metal1 9706 6358 9706 6358 0 _114_
rlabel metal1 8694 5746 8694 5746 0 _115_
rlabel metal1 7452 5202 7452 5202 0 _116_
rlabel metal1 7682 4692 7682 4692 0 _117_
rlabel metal1 6670 5100 6670 5100 0 _118_
rlabel metal1 5704 9010 5704 9010 0 _119_
rlabel metal2 10442 6562 10442 6562 0 _120_
rlabel metal1 8326 5644 8326 5644 0 _121_
rlabel metal1 7176 6970 7176 6970 0 _122_
rlabel metal1 8694 5100 8694 5100 0 _123_
rlabel metal1 7360 8398 7360 8398 0 _124_
rlabel metal1 6118 8466 6118 8466 0 _125_
rlabel metal1 2277 7174 2277 7174 0 _126_
rlabel metal2 3358 7650 3358 7650 0 _127_
rlabel metal1 5060 7922 5060 7922 0 _128_
rlabel metal1 1886 9010 1886 9010 0 _129_
rlabel metal1 11868 8058 11868 8058 0 _130_
rlabel metal1 4554 9044 4554 9044 0 _131_
rlabel metal1 4876 7514 4876 7514 0 _132_
rlabel metal1 2346 8466 2346 8466 0 _133_
rlabel metal1 3772 8058 3772 8058 0 _134_
rlabel metal1 2116 9486 2116 9486 0 _135_
rlabel metal2 6946 8126 6946 8126 0 _136_
rlabel metal1 5106 8466 5106 8466 0 _137_
rlabel metal1 3312 11050 3312 11050 0 _138_
rlabel metal2 2530 10404 2530 10404 0 _139_
rlabel metal2 3818 12789 3818 12789 0 _140_
rlabel metal1 1886 13838 1886 13838 0 _141_
rlabel metal1 2691 13430 2691 13430 0 _142_
rlabel metal1 4370 14484 4370 14484 0 _143_
rlabel metal1 4646 11016 4646 11016 0 _144_
rlabel metal2 2806 12036 2806 12036 0 _145_
rlabel metal2 4646 12585 4646 12585 0 _146_
rlabel metal1 2070 12716 2070 12716 0 _147_
rlabel metal1 4094 13940 4094 13940 0 _148_
rlabel metal1 3542 13906 3542 13906 0 _149_
rlabel metal1 14536 3502 14536 3502 0 ccff_head
rlabel metal1 14628 4794 14628 4794 0 ccff_tail
rlabel metal3 820 3060 820 3060 0 chanx_left_in[0]
rlabel metal3 820 4420 820 4420 0 chanx_left_in[1]
rlabel metal3 958 5780 958 5780 0 chanx_left_in[2]
rlabel metal3 751 7140 751 7140 0 chanx_left_in[3]
rlabel metal3 820 8500 820 8500 0 chanx_left_in[4]
rlabel metal3 820 9860 820 9860 0 chanx_left_in[5]
rlabel metal3 820 11220 820 11220 0 chanx_left_in[6]
rlabel metal3 820 12580 820 12580 0 chanx_left_in[7]
rlabel metal3 820 13940 820 13940 0 chanx_left_in[8]
rlabel metal2 506 1792 506 1792 0 chanx_left_out[0]
rlabel metal2 1334 1554 1334 1554 0 chanx_left_out[1]
rlabel metal2 2162 1554 2162 1554 0 chanx_left_out[2]
rlabel metal2 2990 1554 2990 1554 0 chanx_left_out[3]
rlabel metal2 3818 1554 3818 1554 0 chanx_left_out[4]
rlabel metal2 4646 823 4646 823 0 chanx_left_out[5]
rlabel metal2 5474 1571 5474 1571 0 chanx_left_out[6]
rlabel metal2 6302 1554 6302 1554 0 chanx_left_out[7]
rlabel metal2 7130 959 7130 959 0 chanx_left_out[8]
rlabel metal1 14490 6256 14490 6256 0 chanx_right_in[0]
rlabel metal1 14720 7378 14720 7378 0 chanx_right_in[1]
rlabel metal1 14674 8942 14674 8942 0 chanx_right_in[2]
rlabel metal1 14720 10030 14720 10030 0 chanx_right_in[3]
rlabel metal2 14490 10931 14490 10931 0 chanx_right_in[4]
rlabel metal2 14490 12665 14490 12665 0 chanx_right_in[5]
rlabel via2 14490 13923 14490 13923 0 chanx_right_in[6]
rlabel metal1 14536 14382 14536 14382 0 chanx_right_in[7]
rlabel metal1 13156 16694 13156 16694 0 chanx_right_in[8]
rlabel metal2 7958 823 7958 823 0 chanx_right_out[0]
rlabel metal2 8786 1520 8786 1520 0 chanx_right_out[1]
rlabel metal2 9614 1571 9614 1571 0 chanx_right_out[2]
rlabel metal2 10442 1520 10442 1520 0 chanx_right_out[3]
rlabel metal2 11270 959 11270 959 0 chanx_right_out[4]
rlabel metal2 12098 959 12098 959 0 chanx_right_out[5]
rlabel metal2 12926 1520 12926 1520 0 chanx_right_out[6]
rlabel metal2 13754 1792 13754 1792 0 chanx_right_out[7]
rlabel metal2 14582 1095 14582 1095 0 chanx_right_out[8]
rlabel metal1 1978 16626 1978 16626 0 chany_top_in[0]
rlabel metal1 1794 17204 1794 17204 0 chany_top_in[1]
rlabel metal1 2300 17170 2300 17170 0 chany_top_in[2]
rlabel metal1 2622 16524 2622 16524 0 chany_top_in[3]
rlabel metal1 2622 17204 2622 17204 0 chany_top_in[4]
rlabel metal1 3082 17170 3082 17170 0 chany_top_in[5]
rlabel metal1 4232 17170 4232 17170 0 chany_top_in[6]
rlabel metal1 6394 17136 6394 17136 0 chany_top_in[7]
rlabel metal1 6946 17136 6946 17136 0 chany_top_in[8]
rlabel metal1 9200 17306 9200 17306 0 chany_top_out[0]
rlabel metal1 9890 17306 9890 17306 0 chany_top_out[1]
rlabel metal1 10626 17306 10626 17306 0 chany_top_out[2]
rlabel metal1 11408 17306 11408 17306 0 chany_top_out[3]
rlabel metal1 12144 17306 12144 17306 0 chany_top_out[4]
rlabel metal1 12880 17306 12880 17306 0 chany_top_out[5]
rlabel metal1 13662 17306 13662 17306 0 chany_top_out[6]
rlabel metal1 14030 16762 14030 16762 0 chany_top_out[7]
rlabel metal2 14996 17884 14996 17884 0 chany_top_out[8]
rlabel metal1 7866 12920 7866 12920 0 clknet_0_prog_clk
rlabel metal1 4140 6834 4140 6834 0 clknet_2_0__leaf_prog_clk
rlabel metal1 6026 12274 6026 12274 0 clknet_2_1__leaf_prog_clk
rlabel metal1 11868 8942 11868 8942 0 clknet_2_2__leaf_prog_clk
rlabel metal2 9062 15232 9062 15232 0 clknet_2_3__leaf_prog_clk
rlabel metal3 1050 18020 1050 18020 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1326 16660 1326 16660 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 12098 9452 12098 9452 0 mem_left_track_1.DFF_0_.D
rlabel metal1 10626 8806 10626 8806 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 1748 6290 1748 6290 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 2714 6290 2714 6290 0 mem_left_track_1.DFF_2_.Q
rlabel metal1 4922 11798 4922 11798 0 mem_left_track_17.DFF_0_.D
rlabel metal1 6808 9554 6808 9554 0 mem_left_track_17.DFF_0_.Q
rlabel metal1 8970 9996 8970 9996 0 mem_left_track_17.DFF_1_.Q
rlabel metal2 1978 9996 1978 9996 0 mem_left_track_9.DFF_0_.Q
rlabel metal1 1978 11730 1978 11730 0 mem_left_track_9.DFF_1_.Q
rlabel metal1 13248 11866 13248 11866 0 mem_right_track_0.DFF_0_.D
rlabel metal1 9430 13294 9430 13294 0 mem_right_track_0.DFF_0_.Q
rlabel metal2 6210 13090 6210 13090 0 mem_right_track_0.DFF_1_.Q
rlabel metal1 7682 12070 7682 12070 0 mem_right_track_0.DFF_2_.Q
rlabel metal1 9062 6188 9062 6188 0 mem_right_track_16.DFF_0_.D
rlabel metal1 7544 9486 7544 9486 0 mem_right_track_16.DFF_0_.Q
rlabel metal2 10994 11356 10994 11356 0 mem_right_track_16.DFF_1_.Q
rlabel metal1 6394 5644 6394 5644 0 mem_right_track_8.DFF_0_.Q
rlabel metal1 6854 5678 6854 5678 0 mem_right_track_8.DFF_1_.Q
rlabel metal1 13570 13498 13570 13498 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 3864 15470 3864 15470 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 5612 17170 5612 17170 0 mem_top_track_0.DFF_2_.Q
rlabel metal1 10488 14994 10488 14994 0 mem_top_track_14.DFF_0_.D
rlabel metal1 11822 13906 11822 13906 0 mem_top_track_14.DFF_0_.Q
rlabel metal2 13386 14790 13386 14790 0 mem_top_track_14.DFF_1_.Q
rlabel metal2 12558 13260 12558 13260 0 mem_top_track_16.DFF_0_.Q
rlabel metal2 13386 11968 13386 11968 0 mem_top_track_16.DFF_1_.Q
rlabel metal1 9982 15402 9982 15402 0 mem_top_track_2.DFF_0_.Q
rlabel metal1 8096 16082 8096 16082 0 mem_top_track_2.DFF_1_.Q
rlabel metal1 9430 14382 9430 14382 0 mem_top_track_8.DFF_0_.Q
rlabel metal1 5014 8398 5014 8398 0 mux_left_track_1.INVTX1_0_.out
rlabel metal2 4968 14382 4968 14382 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 4968 17510 4968 17510 0 mux_left_track_1.INVTX1_2_.out
rlabel metal1 12236 8398 12236 8398 0 mux_left_track_1.INVTX1_3_.out
rlabel metal2 2530 9316 2530 9316 0 mux_left_track_1.INVTX1_4_.out
rlabel metal1 1840 8942 1840 8942 0 mux_left_track_1.INVTX1_5_.out
rlabel metal1 4784 8602 4784 8602 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5934 7820 5934 7820 0 mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 2300 9146 2300 9146 0 mux_left_track_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 5106 8058 5106 8058 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 3404 6766 3404 6766 0 mux_left_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 2162 3060 2162 3060 0 mux_left_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 5796 10030 5796 10030 0 mux_left_track_17.INVTX1_0_.out
rlabel metal1 4324 16422 4324 16422 0 mux_left_track_17.INVTX1_1_.out
rlabel metal2 6854 11730 6854 11730 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 7544 8806 7544 8806 0 mux_left_track_17.INVTX1_3_.out
rlabel metal1 9752 12954 9752 12954 0 mux_left_track_17.INVTX1_4_.out
rlabel metal1 6716 11254 6716 11254 0 mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7912 10642 7912 10642 0 mux_left_track_17.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9844 10438 9844 10438 0 mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9890 7990 9890 7990 0 mux_left_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 10212 8330 10212 8330 0 mux_left_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3956 14994 3956 14994 0 mux_left_track_9.INVTX1_0_.out
rlabel metal1 5382 14484 5382 14484 0 mux_left_track_9.INVTX1_1_.out
rlabel metal1 6946 14382 6946 14382 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 3036 13294 3036 13294 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 2323 12818 2323 12818 0 mux_left_track_9.INVTX1_4_.out
rlabel metal1 2024 13906 2024 13906 0 mux_left_track_9.INVTX1_5_.out
rlabel metal1 4048 14246 4048 14246 0 mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 3634 13600 3634 13600 0 mux_left_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 2530 13328 2530 13328 0 mux_left_track_9.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 4784 12614 4784 12614 0 mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2990 11016 2990 11016 0 mux_left_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 4094 7038 4094 7038 0 mux_left_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 14214 15028 14214 15028 0 mux_right_track_0.INVTX1_3_.out
rlabel metal1 5382 12750 5382 12750 0 mux_right_track_0.INVTX1_4_.out
rlabel metal1 5474 12206 5474 12206 0 mux_right_track_0.INVTX1_5_.out
rlabel metal1 6440 14586 6440 14586 0 mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 8096 14518 8096 14518 0 mux_right_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 6256 12818 6256 12818 0 mux_right_track_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 8004 14450 8004 14450 0 mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7268 12614 7268 12614 0 mux_right_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 8326 8194 8326 8194 0 mux_right_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 10810 13124 10810 13124 0 mux_right_track_16.INVTX1_3_.out
rlabel metal1 10258 12274 10258 12274 0 mux_right_track_16.INVTX1_4_.out
rlabel metal2 6762 10336 6762 10336 0 mux_right_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9660 11050 9660 11050 0 mux_right_track_16.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 10764 10438 10764 10438 0 mux_right_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10672 11866 10672 11866 0 mux_right_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 11592 10098 11592 10098 0 mux_right_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 6762 4794 6762 4794 0 mux_right_track_8.INVTX1_3_.out
rlabel metal1 12466 5168 12466 5168 0 mux_right_track_8.INVTX1_4_.out
rlabel metal1 7912 4590 7912 4590 0 mux_right_track_8.INVTX1_5_.out
rlabel metal1 6256 8602 6256 8602 0 mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7176 5338 7176 5338 0 mux_right_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 8234 5508 8234 5508 0 mux_right_track_8.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 7452 7174 7452 7174 0 mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9292 5882 9292 5882 0 mux_right_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 9936 6154 9936 6154 0 mux_right_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 2162 16116 2162 16116 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 14122 15130 14122 15130 0 mux_top_track_0.INVTX1_2_.out
rlabel metal2 3818 14246 3818 14246 0 mux_top_track_0.INVTX1_4_.out
rlabel metal1 4186 15538 4186 15538 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5566 15572 5566 15572 0 mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 5704 15674 5704 15674 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 4554 16864 4554 16864 0 mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 6670 16014 6670 16014 0 mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3542 13464 3542 13464 0 mux_top_track_14.INVTX1_1_.out
rlabel metal1 12834 14892 12834 14892 0 mux_top_track_14.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13248 15674 13248 15674 0 mux_top_track_14.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 14168 9486 14168 9486 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 1702 12104 1702 12104 0 mux_top_track_16.INVTX1_3_.out
rlabel metal1 13294 9656 13294 9656 0 mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13570 10234 13570 10234 0 mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13478 11662 13478 11662 0 mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel via1 12558 16677 12558 16677 0 mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 8050 17068 8050 17068 0 mux_top_track_2.INVTX1_0_.out
rlabel metal2 11086 16490 11086 16490 0 mux_top_track_2.INVTX1_2_.out
rlabel metal2 8510 16320 8510 16320 0 mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9844 16490 9844 16490 0 mux_top_track_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9936 16626 9936 16626 0 mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10442 13498 10442 13498 0 mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 11546 15402 11546 15402 0 mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 14168 3706 14168 3706 0 net1
rlabel metal1 1656 13294 1656 13294 0 net10
rlabel metal1 8372 13498 8372 13498 0 net100
rlabel metal2 2530 7650 2530 7650 0 net101
rlabel metal1 6210 15130 6210 15130 0 net102
rlabel metal1 14306 6222 14306 6222 0 net11
rlabel metal1 14306 6392 14306 6392 0 net12
rlabel metal1 13271 8806 13271 8806 0 net13
rlabel metal1 14306 9622 14306 9622 0 net14
rlabel metal1 12650 11118 12650 11118 0 net15
rlabel metal1 13754 12750 13754 12750 0 net16
rlabel metal2 14214 13566 14214 13566 0 net17
rlabel metal2 14306 14790 14306 14790 0 net18
rlabel metal1 13570 16762 13570 16762 0 net19
rlabel metal1 1610 3570 1610 3570 0 net2
rlabel via1 2898 16405 2898 16405 0 net20
rlabel metal2 1932 16966 1932 16966 0 net21
rlabel metal2 2254 16014 2254 16014 0 net22
rlabel metal1 2852 16558 2852 16558 0 net23
rlabel metal1 3450 16592 3450 16592 0 net24
rlabel metal1 4738 14994 4738 14994 0 net25
rlabel metal1 3404 17170 3404 17170 0 net26
rlabel metal1 6624 17170 6624 17170 0 net27
rlabel metal1 8510 15470 8510 15470 0 net28
rlabel metal1 1610 16456 1610 16456 0 net29
rlabel metal1 8970 4080 8970 4080 0 net3
rlabel metal1 1840 16082 1840 16082 0 net30
rlabel metal2 14306 3536 14306 3536 0 net31
rlabel metal1 14122 15504 14122 15504 0 net32
rlabel metal2 1702 16864 1702 16864 0 net33
rlabel metal1 7452 17170 7452 17170 0 net34
rlabel metal1 9591 8330 9591 8330 0 net35
rlabel metal1 1932 3026 1932 3026 0 net36
rlabel metal1 1794 2312 1794 2312 0 net37
rlabel metal1 2852 2414 2852 2414 0 net38
rlabel metal1 3450 2448 3450 2448 0 net39
rlabel metal2 2530 5984 2530 5984 0 net4
rlabel metal1 4232 2414 4232 2414 0 net40
rlabel metal1 4784 2414 4784 2414 0 net41
rlabel metal2 5750 7412 5750 7412 0 net42
rlabel metal1 6670 2414 6670 2414 0 net43
rlabel metal1 8050 2346 8050 2346 0 net44
rlabel metal1 8326 2822 8326 2822 0 net45
rlabel metal1 9062 2448 9062 2448 0 net46
rlabel metal1 9844 2414 9844 2414 0 net47
rlabel metal1 10442 2414 10442 2414 0 net48
rlabel metal1 11408 2414 11408 2414 0 net49
rlabel metal1 1564 5882 1564 5882 0 net5
rlabel metal1 12190 2414 12190 2414 0 net50
rlabel metal1 12880 2414 12880 2414 0 net51
rlabel metal1 13708 10438 13708 10438 0 net52
rlabel metal1 13754 3094 13754 3094 0 net53
rlabel metal1 8970 16762 8970 16762 0 net54
rlabel metal2 11730 17000 11730 17000 0 net55
rlabel metal1 11546 17102 11546 17102 0 net56
rlabel metal2 11914 16966 11914 16966 0 net57
rlabel metal1 11960 16218 11960 16218 0 net58
rlabel metal2 12650 16966 12650 16966 0 net59
rlabel metal2 12466 13056 12466 13056 0 net6
rlabel metal1 13110 16762 13110 16762 0 net60
rlabel metal1 13616 16218 13616 16218 0 net61
rlabel metal1 13271 16150 13271 16150 0 net62
rlabel metal1 2530 17068 2530 17068 0 net63
rlabel metal2 11546 12585 11546 12585 0 net64
rlabel metal2 9062 8364 9062 8364 0 net65
rlabel metal1 10534 15538 10534 15538 0 net66
rlabel metal1 11224 15538 11224 15538 0 net67
rlabel metal1 12650 15470 12650 15470 0 net68
rlabel metal2 11914 12988 11914 12988 0 net69
rlabel metal1 12466 4590 12466 4590 0 net7
rlabel metal1 7130 12818 7130 12818 0 net70
rlabel metal1 10120 5746 10120 5746 0 net71
rlabel metal2 3082 7293 3082 7293 0 net72
rlabel metal1 2530 10642 2530 10642 0 net73
rlabel metal1 7401 8874 7401 8874 0 net74
rlabel metal1 4354 10710 4354 10710 0 net75
rlabel metal1 11458 14382 11458 14382 0 net76
rlabel metal1 6803 15470 6803 15470 0 net77
rlabel metal2 8510 6562 8510 6562 0 net78
rlabel via1 11642 8942 11642 8942 0 net79
rlabel metal2 1610 11424 1610 11424 0 net8
rlabel metal2 12742 14586 12742 14586 0 net80
rlabel metal1 12650 12172 12650 12172 0 net81
rlabel metal1 12834 14008 12834 14008 0 net82
rlabel via1 9342 13974 9342 13974 0 net83
rlabel metal1 9379 14314 9379 14314 0 net84
rlabel metal1 11990 10710 11990 10710 0 net85
rlabel metal1 3864 8602 3864 8602 0 net86
rlabel metal1 8376 16150 8376 16150 0 net87
rlabel metal2 7682 6086 7682 6086 0 net88
rlabel metal1 7084 9690 7084 9690 0 net89
rlabel metal2 1610 12682 1610 12682 0 net9
rlabel metal2 12650 11526 12650 11526 0 net90
rlabel metal1 10253 9554 10253 9554 0 net91
rlabel metal1 5883 6766 5883 6766 0 net92
rlabel metal1 7866 9622 7866 9622 0 net93
rlabel metal1 5101 16150 5101 16150 0 net94
rlabel metal1 2655 6766 2655 6766 0 net95
rlabel metal2 2530 10914 2530 10914 0 net96
rlabel metal1 6849 12206 6849 12206 0 net97
rlabel metal1 2882 11798 2882 11798 0 net98
rlabel via1 8413 8466 8413 8466 0 net99
rlabel metal2 4094 15351 4094 15351 0 prog_clk
rlabel metal1 14536 2414 14536 2414 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 12374 17051 12374 17051 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 1242 17170 1242 17170 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 7682 17238 7682 17238 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
<< properties >>
string FIXED_BBOX 0 0 16000 20000
<< end >>
