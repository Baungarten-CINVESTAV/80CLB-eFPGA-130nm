VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN bottom_width_0_height_0_subtile_0__pin_I_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_I_2_
  PIN bottom_width_0_height_0_subtile_0__pin_I_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_I_6_
  PIN bottom_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_O_0_
  PIN bottom_width_0_height_0_subtile_0__pin_clk_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_clk_0_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 110.200 150.000 110.800 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 134.680 150.000 135.280 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END clk
  PIN left_width_0_height_0_subtile_0__pin_I_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END left_width_0_height_0_subtile_0__pin_I_3_
  PIN left_width_0_height_0_subtile_0__pin_I_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END left_width_0_height_0_subtile_0__pin_I_7_
  PIN left_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END left_width_0_height_0_subtile_0__pin_O_1_
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END prog_clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END reset
  PIN right_width_0_height_0_subtile_0__pin_I_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 12.280 150.000 12.880 ;
    END
  END right_width_0_height_0_subtile_0__pin_I_1_
  PIN right_width_0_height_0_subtile_0__pin_I_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 146.000 36.760 150.000 37.360 ;
    END
  END right_width_0_height_0_subtile_0__pin_I_5_
  PIN right_width_0_height_0_subtile_0__pin_I_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 150.000 61.840 ;
    END
  END right_width_0_height_0_subtile_0__pin_I_9_
  PIN right_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.720 150.000 86.320 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_3_
  PIN set
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END set
  PIN top_width_0_height_0_subtile_0__pin_I_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 146.000 19.230 150.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I_0_
  PIN top_width_0_height_0_subtile_0__pin_I_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 146.000 56.490 150.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I_4_
  PIN top_width_0_height_0_subtile_0__pin_I_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_I_8_
  PIN top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.730 146.000 131.010 150.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_2_
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 138.960 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 4.670 8.200 145.240 139.360 ;
      LAYER met2 ;
        RECT 4.690 145.720 18.670 146.000 ;
        RECT 19.510 145.720 55.930 146.000 ;
        RECT 56.770 145.720 93.190 146.000 ;
        RECT 94.030 145.720 130.450 146.000 ;
        RECT 131.290 145.720 145.210 146.000 ;
        RECT 4.690 4.280 145.210 145.720 ;
        RECT 4.690 3.670 18.670 4.280 ;
        RECT 19.510 3.670 55.930 4.280 ;
        RECT 56.770 3.670 93.190 4.280 ;
        RECT 94.030 3.670 130.450 4.280 ;
        RECT 131.290 3.670 145.210 4.280 ;
      LAYER met3 ;
        RECT 4.000 137.040 146.000 138.885 ;
        RECT 4.400 135.680 146.000 137.040 ;
        RECT 4.400 135.640 145.600 135.680 ;
        RECT 4.000 134.280 145.600 135.640 ;
        RECT 4.000 119.360 146.000 134.280 ;
        RECT 4.400 117.960 146.000 119.360 ;
        RECT 4.000 111.200 146.000 117.960 ;
        RECT 4.000 109.800 145.600 111.200 ;
        RECT 4.000 101.680 146.000 109.800 ;
        RECT 4.400 100.280 146.000 101.680 ;
        RECT 4.000 86.720 146.000 100.280 ;
        RECT 4.000 85.320 145.600 86.720 ;
        RECT 4.000 84.000 146.000 85.320 ;
        RECT 4.400 82.600 146.000 84.000 ;
        RECT 4.000 66.320 146.000 82.600 ;
        RECT 4.400 64.920 146.000 66.320 ;
        RECT 4.000 62.240 146.000 64.920 ;
        RECT 4.000 60.840 145.600 62.240 ;
        RECT 4.000 48.640 146.000 60.840 ;
        RECT 4.400 47.240 146.000 48.640 ;
        RECT 4.000 37.760 146.000 47.240 ;
        RECT 4.000 36.360 145.600 37.760 ;
        RECT 4.000 30.960 146.000 36.360 ;
        RECT 4.400 29.560 146.000 30.960 ;
        RECT 4.000 13.280 146.000 29.560 ;
        RECT 4.000 11.880 145.600 13.280 ;
        RECT 4.000 9.700 146.000 11.880 ;
      LAYER met4 ;
        RECT 24.215 10.240 39.050 90.265 ;
        RECT 41.450 10.240 56.415 90.265 ;
        RECT 58.815 10.240 73.780 90.265 ;
        RECT 76.180 10.240 91.145 90.265 ;
        RECT 93.545 10.240 108.510 90.265 ;
        RECT 110.910 10.240 125.875 90.265 ;
        RECT 128.275 10.240 130.345 90.265 ;
        RECT 24.215 9.695 130.345 10.240 ;
  END
END grid_clb
END LIBRARY

