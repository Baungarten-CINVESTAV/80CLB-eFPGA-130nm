magic
tech sky130A
magscale 1 2
timestamp 1707850049
<< viali >>
rect 1409 9605 1443 9639
rect 1961 9605 1995 9639
rect 2973 9605 3007 9639
rect 3985 9605 4019 9639
rect 4997 9605 5031 9639
rect 6377 9605 6411 9639
rect 7021 9605 7055 9639
rect 8033 9605 8067 9639
rect 9505 9605 9539 9639
rect 1777 9537 1811 9571
rect 2329 9537 2363 9571
rect 3341 9537 3375 9571
rect 4353 9537 4387 9571
rect 5365 9537 5399 9571
rect 6745 9537 6779 9571
rect 7389 9537 7423 9571
rect 8401 9537 8435 9571
rect 8585 9537 8619 9571
rect 9137 9537 9171 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10333 9401 10367 9435
rect 8769 9333 8803 9367
rect 9781 9333 9815 9367
rect 3341 9129 3375 9163
rect 4353 9129 4387 9163
rect 7481 9129 7515 9163
rect 9137 9129 9171 9163
rect 10241 9129 10275 9163
rect 4721 8993 4755 9027
rect 5549 8993 5583 9027
rect 9321 8993 9355 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 3525 8925 3559 8959
rect 4077 8925 4111 8959
rect 4537 8925 4571 8959
rect 4905 8925 4939 8959
rect 5457 8925 5491 8959
rect 7389 8925 7423 8959
rect 7665 8925 7699 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 9505 8925 9539 8959
rect 9873 8857 9907 8891
rect 10149 8857 10183 8891
rect 1593 8789 1627 8823
rect 1869 8789 1903 8823
rect 2145 8789 2179 8823
rect 4261 8789 4295 8823
rect 5365 8789 5399 8823
rect 6469 8789 6503 8823
rect 7297 8789 7331 8823
rect 4905 8585 4939 8619
rect 9873 8585 9907 8619
rect 10149 8585 10183 8619
rect 1409 8449 1443 8483
rect 4997 8449 5031 8483
rect 5549 8449 5583 8483
rect 6469 8449 6503 8483
rect 8125 8449 8159 8483
rect 9597 8449 9631 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 5733 8381 5767 8415
rect 6653 8381 6687 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 8309 8381 8343 8415
rect 1593 8313 1627 8347
rect 6193 8313 6227 8347
rect 6837 8313 6871 8347
rect 8033 8313 8067 8347
rect 8493 8313 8527 8347
rect 9781 8313 9815 8347
rect 5089 8041 5123 8075
rect 6561 8041 6595 8075
rect 7573 8041 7607 8075
rect 7757 8041 7791 8075
rect 5457 7973 5491 8007
rect 5733 7973 5767 8007
rect 7205 7973 7239 8007
rect 5825 7905 5859 7939
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 4997 7837 5031 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 6745 7837 6779 7871
rect 7021 7837 7055 7871
rect 7389 7837 7423 7871
rect 7665 7837 7699 7871
rect 8953 7837 8987 7871
rect 9209 7837 9243 7871
rect 10333 7701 10367 7735
rect 4721 7497 4755 7531
rect 7941 7497 7975 7531
rect 10425 7497 10459 7531
rect 1409 7361 1443 7395
rect 4537 7361 4571 7395
rect 5080 7361 5114 7395
rect 8125 7361 8159 7395
rect 10333 7361 10367 7395
rect 4813 7293 4847 7327
rect 7021 7293 7055 7327
rect 7849 7293 7883 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 6193 7225 6227 7259
rect 1593 7157 1627 7191
rect 6469 7157 6503 7191
rect 7205 7157 7239 7191
rect 9965 7157 9999 7191
rect 5273 6953 5307 6987
rect 9413 6953 9447 6987
rect 5181 6885 5215 6919
rect 10333 6885 10367 6919
rect 3801 6749 3835 6783
rect 5917 6749 5951 6783
rect 6193 6749 6227 6783
rect 6377 6749 6411 6783
rect 6633 6749 6667 6783
rect 7849 6749 7883 6783
rect 8585 6749 8619 6783
rect 8953 6749 8987 6783
rect 9781 6749 9815 6783
rect 9965 6749 9999 6783
rect 10057 6749 10091 6783
rect 10517 6749 10551 6783
rect 4068 6681 4102 6715
rect 6009 6613 6043 6647
rect 7757 6613 7791 6647
rect 8493 6613 8527 6647
rect 8677 6613 8711 6647
rect 9137 6613 9171 6647
rect 2329 6409 2363 6443
rect 6009 6409 6043 6443
rect 7113 6409 7147 6443
rect 10333 6409 10367 6443
rect 8502 6341 8536 6375
rect 1409 6273 1443 6307
rect 2513 6273 2547 6307
rect 3985 6273 4019 6307
rect 4445 6273 4479 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 8769 6273 8803 6307
rect 10517 6273 10551 6307
rect 5089 6205 5123 6239
rect 8861 6205 8895 6239
rect 9045 6205 9079 6239
rect 9597 6205 9631 6239
rect 6745 6137 6779 6171
rect 1593 6069 1627 6103
rect 4077 6069 4111 6103
rect 4261 6069 4295 6103
rect 4629 6069 4663 6103
rect 4905 6069 4939 6103
rect 5733 6069 5767 6103
rect 6929 6069 6963 6103
rect 7389 6069 7423 6103
rect 9413 6069 9447 6103
rect 10241 6069 10275 6103
rect 5641 5865 5675 5899
rect 5549 5797 5583 5831
rect 4169 5729 4203 5763
rect 5089 5729 5123 5763
rect 3433 5661 3467 5695
rect 3893 5661 3927 5695
rect 4353 5661 4387 5695
rect 4905 5661 4939 5695
rect 5825 5661 5859 5695
rect 6193 5661 6227 5695
rect 8677 5661 8711 5695
rect 10158 5661 10192 5695
rect 10425 5661 10459 5695
rect 4813 5593 4847 5627
rect 6469 5593 6503 5627
rect 3617 5525 3651 5559
rect 3985 5525 4019 5559
rect 6285 5525 6319 5559
rect 7757 5525 7791 5559
rect 8493 5525 8527 5559
rect 9045 5525 9079 5559
rect 3065 5321 3099 5355
rect 5089 5321 5123 5355
rect 9137 5321 9171 5355
rect 10425 5321 10459 5355
rect 4353 5253 4387 5287
rect 7849 5253 7883 5287
rect 1409 5185 1443 5219
rect 1777 5185 1811 5219
rect 4629 5185 4663 5219
rect 5365 5185 5399 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6469 5185 6503 5219
rect 6745 5185 6779 5219
rect 7297 5185 7331 5219
rect 9781 5185 9815 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 4445 5117 4479 5151
rect 7113 5117 7147 5151
rect 7757 5117 7791 5151
rect 5917 5049 5951 5083
rect 6561 5049 6595 5083
rect 10057 5049 10091 5083
rect 1593 4981 1627 5015
rect 1961 4981 1995 5015
rect 5181 4981 5215 5015
rect 6193 4981 6227 5015
rect 6837 4981 6871 5015
rect 9965 4981 9999 5015
rect 4445 4777 4479 4811
rect 4997 4777 5031 4811
rect 7665 4777 7699 4811
rect 3341 4709 3375 4743
rect 10057 4709 10091 4743
rect 3525 4641 3559 4675
rect 3985 4641 4019 4675
rect 4813 4641 4847 4675
rect 6469 4641 6503 4675
rect 7205 4641 7239 4675
rect 7757 4641 7791 4675
rect 7941 4641 7975 4675
rect 8401 4641 8435 4675
rect 9689 4641 9723 4675
rect 3157 4573 3191 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 4629 4573 4663 4607
rect 6285 4573 6319 4607
rect 7021 4573 7055 4607
rect 8677 4573 8711 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 8585 4505 8619 4539
rect 6929 4437 6963 4471
rect 8953 4437 8987 4471
rect 4169 4233 4203 4267
rect 4537 4233 4571 4267
rect 7205 4233 7239 4267
rect 9781 4165 9815 4199
rect 9873 4165 9907 4199
rect 1409 4097 1443 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 4905 4097 4939 4131
rect 5917 4097 5951 4131
rect 6009 4097 6043 4131
rect 6561 4097 6595 4131
rect 7573 4097 7607 4131
rect 7665 4097 7699 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 9597 4097 9631 4131
rect 6745 4029 6779 4063
rect 7849 4029 7883 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 1593 3961 1627 3995
rect 4721 3961 4755 3995
rect 7481 3961 7515 3995
rect 8861 3961 8895 3995
rect 10333 3961 10367 3995
rect 8309 3893 8343 3927
rect 8585 3893 8619 3927
rect 3065 3689 3099 3723
rect 5549 3689 5583 3723
rect 5917 3689 5951 3723
rect 8309 3689 8343 3723
rect 10333 3689 10367 3723
rect 6377 3553 6411 3587
rect 7849 3553 7883 3587
rect 8769 3553 8803 3587
rect 8953 3553 8987 3587
rect 2697 3485 2731 3519
rect 2973 3485 3007 3519
rect 4905 3485 4939 3519
rect 5089 3485 5123 3519
rect 6101 3485 6135 3519
rect 6285 3485 6319 3519
rect 6644 3485 6678 3519
rect 8033 3485 8067 3519
rect 9220 3417 9254 3451
rect 2881 3349 2915 3383
rect 7757 3349 7791 3383
rect 5273 3145 5307 3179
rect 5917 3145 5951 3179
rect 6745 3145 6779 3179
rect 7389 3145 7423 3179
rect 8125 3145 8159 3179
rect 9137 3145 9171 3179
rect 9873 3077 9907 3111
rect 10425 3077 10459 3111
rect 1409 3009 1443 3043
rect 1777 3009 1811 3043
rect 2053 3009 2087 3043
rect 2513 3009 2547 3043
rect 5089 3009 5123 3043
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 6193 3009 6227 3043
rect 6561 3009 6595 3043
rect 6653 3009 6687 3043
rect 6929 3009 6963 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8217 3009 8251 3043
rect 9413 3009 9447 3043
rect 8493 2941 8527 2975
rect 9781 2941 9815 2975
rect 1593 2873 1627 2907
rect 2329 2873 2363 2907
rect 6101 2873 6135 2907
rect 6377 2873 6411 2907
rect 7849 2873 7883 2907
rect 8309 2873 8343 2907
rect 9597 2873 9631 2907
rect 1961 2805 1995 2839
rect 2237 2805 2271 2839
rect 4905 2805 4939 2839
rect 5641 2805 5675 2839
rect 7113 2805 7147 2839
rect 9597 2601 9631 2635
rect 5733 2533 5767 2567
rect 8585 2533 8619 2567
rect 7849 2465 7883 2499
rect 1777 2397 1811 2431
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4077 2397 4111 2431
rect 5365 2397 5399 2431
rect 5917 2397 5951 2431
rect 6193 2397 6227 2431
rect 6469 2397 6503 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8769 2397 8803 2431
rect 9781 2397 9815 2431
rect 1409 2329 1443 2363
rect 4997 2329 5031 2363
rect 8125 2329 8159 2363
rect 9137 2329 9171 2363
rect 10149 2329 10183 2363
rect 2145 2261 2179 2295
rect 3157 2261 3191 2295
rect 4169 2261 4203 2295
rect 6101 2261 6135 2295
rect 6561 2261 6595 2295
rect 7205 2261 7239 2295
rect 8217 2261 8251 2295
rect 9229 2261 9263 2295
rect 10241 2261 10275 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 9582 9704 9588 9716
rect 8588 9676 9588 9704
rect 842 9596 848 9648
rect 900 9636 906 9648
rect 1397 9639 1455 9645
rect 1397 9636 1409 9639
rect 900 9608 1409 9636
rect 900 9596 906 9608
rect 1397 9605 1409 9608
rect 1443 9605 1455 9639
rect 1397 9599 1455 9605
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 1949 9639 2007 9645
rect 1949 9636 1961 9639
rect 1912 9608 1961 9636
rect 1912 9596 1918 9608
rect 1949 9605 1961 9608
rect 1995 9605 2007 9639
rect 1949 9599 2007 9605
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2924 9608 2973 9636
rect 2924 9596 2930 9608
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 2961 9599 3019 9605
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3936 9608 3985 9636
rect 3936 9596 3942 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 3973 9599 4031 9605
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4948 9608 4997 9636
rect 4948 9596 4954 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 6236 9608 6377 9636
rect 6236 9596 6242 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6972 9608 7021 9636
rect 6972 9596 6978 9608
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 7009 9599 7067 9605
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 7984 9608 8033 9636
rect 7984 9596 7990 9608
rect 8021 9605 8033 9608
rect 8067 9605 8079 9639
rect 8021 9599 8079 9605
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 4338 9528 4344 9580
rect 4396 9528 4402 9580
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 8588 9577 8616 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8996 9608 9505 9636
rect 8996 9596 9002 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9968 9608 10640 9636
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 8404 9500 8432 9531
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9968 9577 9996 9608
rect 10612 9580 10640 9608
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 8938 9500 8944 9512
rect 8404 9472 8944 9500
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 10008 9404 10333 9432
rect 10008 9392 10014 9404
rect 10321 9401 10333 9404
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 8757 9367 8815 9373
rect 8757 9333 8769 9367
rect 8803 9364 8815 9367
rect 9030 9364 9036 9376
rect 8803 9336 9036 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 9272 9336 9781 9364
rect 9272 9324 9278 9336
rect 9769 9333 9781 9336
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 3326 9120 3332 9172
rect 3384 9120 3390 9172
rect 4338 9120 4344 9172
rect 4396 9120 4402 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7432 9132 7481 9160
rect 7432 9120 7438 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 9122 9120 9128 9172
rect 9180 9120 9186 9172
rect 9214 9120 9220 9172
rect 9272 9120 9278 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9364 9132 10241 9160
rect 9364 9120 9370 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 5626 9092 5632 9104
rect 3528 9064 5632 9092
rect 2774 9024 2780 9036
rect 1872 8996 2780 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1872 8956 1900 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 1719 8928 1900 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1946 8916 1952 8968
rect 2004 8916 2010 8968
rect 3528 8965 3556 9064
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 4755 8996 5549 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 9232 9024 9260 9120
rect 10134 9092 10140 9104
rect 9324 9064 10140 9092
rect 9324 9033 9352 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 5537 8987 5595 8993
rect 7392 8996 9260 9024
rect 9309 9027 9367 9033
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4080 8888 4108 8919
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 7392 8965 7420 8996
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 5460 8888 5488 8919
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 8956 8965 8984 8996
rect 9309 8993 9321 9027
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 11054 8956 11060 8968
rect 9539 8928 11060 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 9232 8888 9260 8919
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 1872 8860 5488 8888
rect 8680 8860 9260 8888
rect 1578 8780 1584 8832
rect 1636 8780 1642 8832
rect 1872 8829 1900 8860
rect 8680 8832 8708 8860
rect 9858 8848 9864 8900
rect 9916 8848 9922 8900
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 10100 8860 10149 8888
rect 10100 8848 10106 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 2130 8780 2136 8832
rect 2188 8780 2194 8832
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 5258 8820 5264 8832
rect 4295 8792 5264 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5353 8823 5411 8829
rect 5353 8789 5365 8823
rect 5399 8820 5411 8823
rect 5534 8820 5540 8832
rect 5399 8792 5540 8820
rect 5399 8789 5411 8792
rect 5353 8783 5411 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6972 8792 7297 8820
rect 6972 8780 6978 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 6454 8576 6460 8628
rect 6512 8576 6518 8628
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 8996 8588 9873 8616
rect 8996 8576 9002 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8585 10195 8619
rect 10137 8579 10195 8585
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 6270 8548 6276 8560
rect 1636 8520 6276 8548
rect 1636 8508 1642 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5166 8480 5172 8492
rect 5031 8452 5172 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 6472 8489 6500 8576
rect 6748 8548 6776 8576
rect 10152 8548 10180 8579
rect 6748 8520 10180 8548
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 6604 8452 8125 8480
rect 6604 8440 6610 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9364 8452 9597 8480
rect 9364 8440 9370 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9585 8443 9643 8449
rect 9784 8452 10057 8480
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5684 8384 5733 8412
rect 5684 8372 5690 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 5721 8375 5779 8381
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6840 8384 7389 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 3786 8344 3792 8356
rect 1627 8316 3792 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 6840 8353 6868 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 7558 8372 7564 8424
rect 7616 8372 7622 8424
rect 8294 8372 8300 8424
rect 8352 8372 8358 8424
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6227 8316 6837 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8067 8316 8493 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8481 8313 8493 8316
rect 8527 8344 8539 8347
rect 8662 8344 8668 8356
rect 8527 8316 8668 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 9784 8353 9812 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 10192 8452 10333 8480
rect 10192 8440 10198 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8313 9827 8347
rect 9769 8307 9827 8313
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5626 8072 5632 8084
rect 5123 8044 5632 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6638 8072 6644 8084
rect 6595 8044 6644 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 8294 8072 8300 8084
rect 7791 8044 8300 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 5445 8007 5503 8013
rect 5445 7973 5457 8007
rect 5491 7973 5503 8007
rect 5445 7967 5503 7973
rect 4430 7896 4436 7948
rect 4488 7936 4494 7948
rect 5166 7936 5172 7948
rect 4488 7908 5172 7936
rect 4488 7896 4494 7908
rect 5166 7896 5172 7908
rect 5224 7936 5230 7948
rect 5224 7908 5304 7936
rect 5224 7896 5230 7908
rect 5276 7877 5304 7908
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5261 7871 5319 7877
rect 5031 7840 5212 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5184 7744 5212 7840
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5460 7868 5488 7967
rect 5534 7964 5540 8016
rect 5592 7964 5598 8016
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 8004 5779 8007
rect 7193 8007 7251 8013
rect 5767 7976 6316 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 5552 7936 5580 7964
rect 6288 7945 6316 7976
rect 7193 7973 7205 8007
rect 7239 7973 7251 8007
rect 7193 7967 7251 7973
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 5552 7908 5825 7936
rect 5813 7905 5825 7908
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6914 7936 6920 7948
rect 6503 7908 6920 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5460 7840 5549 7868
rect 5261 7831 5319 7837
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 5276 7732 5304 7831
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7208 7868 7236 7967
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7064 7840 7144 7868
rect 7208 7840 7389 7868
rect 7064 7828 7070 7840
rect 7116 7800 7144 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7668 7800 7696 7831
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9197 7871 9255 7877
rect 9197 7868 9209 7871
rect 9088 7840 9209 7868
rect 9088 7828 9094 7840
rect 9197 7837 9209 7840
rect 9243 7837 9255 7871
rect 9197 7831 9255 7837
rect 7116 7772 7696 7800
rect 7834 7732 7840 7744
rect 5276 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7732 7898 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 7892 7704 10333 7732
rect 7892 7692 7898 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 6638 7528 6644 7540
rect 4755 7500 6644 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 6788 7500 7941 7528
rect 6788 7488 6794 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 9916 7500 10425 7528
rect 9916 7488 9922 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 5074 7401 5080 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 3844 7364 4537 7392
rect 3844 7352 3850 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 5068 7355 5080 7401
rect 5074 7352 5080 7355
rect 5132 7352 5138 7404
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 5960 7364 8125 7392
rect 5960 7352 5966 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 8113 7355 8171 7361
rect 9968 7364 10333 7392
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 4062 7188 4068 7200
rect 1627 7160 4068 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4816 7188 4844 7287
rect 7006 7284 7012 7336
rect 7064 7284 7070 7336
rect 7834 7284 7840 7336
rect 7892 7284 7898 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 8076 7296 9597 7324
rect 8076 7284 8082 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 9858 7324 9864 7336
rect 9815 7296 9864 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 7024 7256 7052 7284
rect 6227 7228 7052 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 5442 7188 5448 7200
rect 4816 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6454 7148 6460 7200
rect 6512 7148 6518 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 6972 7160 7205 7188
rect 6972 7148 6978 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 9968 7197 9996 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9456 7160 9965 7188
rect 9456 7148 9462 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5261 6987 5319 6993
rect 5261 6984 5273 6987
rect 5132 6956 5273 6984
rect 5132 6944 5138 6956
rect 5261 6953 5273 6956
rect 5307 6953 5319 6987
rect 5261 6947 5319 6953
rect 9398 6944 9404 6996
rect 9456 6944 9462 6996
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 5902 6916 5908 6928
rect 5224 6888 5908 6916
rect 5224 6876 5230 6888
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 10321 6919 10379 6925
rect 10321 6885 10333 6919
rect 10367 6885 10379 6919
rect 10321 6879 10379 6885
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5592 6820 6408 6848
rect 5592 6808 5598 6820
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 5552 6780 5580 6808
rect 6380 6792 6408 6820
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 10336 6848 10364 6879
rect 10870 6848 10876 6860
rect 7708 6820 10364 6848
rect 10520 6820 10876 6848
rect 7708 6808 7714 6820
rect 3844 6752 5580 6780
rect 3844 6740 3850 6752
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 6621 6783 6679 6789
rect 6621 6780 6633 6783
rect 6512 6752 6633 6780
rect 6512 6740 6518 6752
rect 6621 6749 6633 6752
rect 6667 6749 6679 6783
rect 6621 6743 6679 6749
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 8588 6789 8616 6820
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 8987 6752 9720 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 4056 6715 4114 6721
rect 4056 6681 4068 6715
rect 4102 6712 4114 6715
rect 6932 6712 6960 6740
rect 4102 6684 6960 6712
rect 4102 6681 4114 6684
rect 4056 6675 4114 6681
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5684 6616 6009 6644
rect 5684 6604 5690 6616
rect 5997 6613 6009 6616
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7852 6644 7880 6743
rect 9692 6656 9720 6752
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 10520 6789 10548 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9999 6752 10057 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 7800 6616 7880 6644
rect 7800 6604 7806 6616
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8168 6616 8493 6644
rect 8168 6604 8174 6616
rect 8481 6613 8493 6616
rect 8527 6613 8539 6647
rect 8481 6607 8539 6613
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 9122 6604 9128 6656
rect 9180 6604 9186 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2498 6440 2504 6452
rect 2363 6412 2504 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 5626 6400 5632 6452
rect 5684 6400 5690 6452
rect 5718 6400 5724 6452
rect 5776 6400 5782 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6178 6440 6184 6452
rect 6043 6412 6184 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 5442 6372 5448 6384
rect 2746 6344 5448 6372
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2746 6304 2774 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 2547 6276 2774 6304
rect 3973 6307 4031 6313
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4019 6276 4108 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4080 6248 4108 6276
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5261 6307 5319 6313
rect 5031 6276 5212 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4724 6168 4752 6267
rect 5074 6196 5080 6248
rect 5132 6196 5138 6248
rect 5184 6236 5212 6276
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5644 6304 5672 6400
rect 5307 6276 5672 6304
rect 5736 6304 5764 6400
rect 7116 6372 7144 6403
rect 7742 6400 7748 6452
rect 7800 6400 7806 6452
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 9824 6412 10333 6440
rect 9824 6400 9830 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 6564 6344 7144 6372
rect 6564 6313 6592 6344
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5736 6276 5825 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5736 6236 5764 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7055 6276 7297 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7285 6273 7297 6276
rect 7331 6304 7343 6307
rect 7760 6304 7788 6400
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8490 6375 8548 6381
rect 8490 6372 8502 6375
rect 8168 6344 8502 6372
rect 8168 6332 8174 6344
rect 8490 6341 8502 6344
rect 8536 6341 8548 6375
rect 8490 6335 8548 6341
rect 7331 6276 7788 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 5184 6208 5764 6236
rect 8680 6236 8708 6400
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 8938 6304 8944 6316
rect 8803 6276 8944 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9140 6304 9168 6400
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 9140 6276 10517 6304
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8680 6208 8861 6236
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 9030 6196 9036 6248
rect 9088 6196 9094 6248
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 9674 6236 9680 6248
rect 9631 6208 9680 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 6733 6171 6791 6177
rect 4724 6140 5856 6168
rect 5828 6112 5856 6140
rect 6733 6137 6745 6171
rect 6779 6168 6791 6171
rect 7466 6168 7472 6180
rect 6779 6140 7472 6168
rect 6779 6137 6791 6140
rect 6733 6131 6791 6137
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 9600 6168 9628 6199
rect 9674 6196 9680 6208
rect 9732 6236 9738 6248
rect 10318 6236 10324 6248
rect 9732 6208 10324 6236
rect 9732 6196 9738 6208
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 9048 6140 9628 6168
rect 1578 6060 1584 6112
rect 1636 6060 1642 6112
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4154 6100 4160 6112
rect 4111 6072 4160 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 4246 6060 4252 6112
rect 4304 6060 4310 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4396 6072 4629 6100
rect 4396 6060 4402 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4617 6063 4675 6069
rect 4893 6103 4951 6109
rect 4893 6069 4905 6103
rect 4939 6100 4951 6103
rect 4982 6100 4988 6112
rect 4939 6072 4988 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 6914 6060 6920 6112
rect 6972 6060 6978 6112
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 9048 6100 9076 6140
rect 7423 6072 9076 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 9398 6060 9404 6112
rect 9456 6060 9462 6112
rect 10226 6060 10232 6112
rect 10284 6060 10290 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 4982 5856 4988 5908
rect 5040 5856 5046 5908
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5408 5868 5641 5896
rect 5408 5856 5414 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 5629 5859 5687 5865
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 8956 5868 10456 5896
rect 4264 5828 4292 5856
rect 3436 5800 4292 5828
rect 3436 5701 3464 5800
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 4356 5760 4384 5856
rect 4203 5732 4384 5760
rect 5000 5760 5028 5856
rect 5537 5831 5595 5837
rect 5537 5797 5549 5831
rect 5583 5828 5595 5831
rect 5718 5828 5724 5840
rect 5583 5800 5724 5828
rect 5583 5797 5595 5800
rect 5537 5791 5595 5797
rect 5718 5788 5724 5800
rect 5776 5828 5782 5840
rect 6564 5828 6592 5856
rect 8956 5840 8984 5868
rect 5776 5800 6592 5828
rect 5776 5788 5782 5800
rect 8938 5788 8944 5840
rect 8996 5788 9002 5840
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 5000 5732 5089 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 7558 5760 7564 5772
rect 5077 5723 5135 5729
rect 6104 5732 7564 5760
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 4246 5692 4252 5704
rect 3936 5664 4252 5692
rect 3936 5652 3942 5664
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 4982 5692 4988 5704
rect 4939 5664 4988 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 4356 5624 4384 5655
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 6104 5692 6132 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7668 5732 8892 5760
rect 5868 5664 6132 5692
rect 6181 5695 6239 5701
rect 5868 5652 5874 5664
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 7668 5692 7696 5732
rect 6227 5664 7696 5692
rect 8665 5695 8723 5701
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 8711 5664 8800 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 3620 5596 4384 5624
rect 4801 5627 4859 5633
rect 3620 5565 3648 5596
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 5074 5624 5080 5636
rect 4847 5596 5080 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6196 5624 6224 5655
rect 5500 5596 6224 5624
rect 5500 5584 5506 5596
rect 6454 5584 6460 5636
rect 6512 5584 6518 5636
rect 8772 5568 8800 5664
rect 8864 5636 8892 5732
rect 10428 5701 10456 5868
rect 10146 5695 10204 5701
rect 10146 5661 10158 5695
rect 10192 5661 10204 5695
rect 10146 5655 10204 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 8846 5584 8852 5636
rect 8904 5584 8910 5636
rect 10152 5624 10180 5655
rect 10226 5624 10232 5636
rect 10152 5596 10232 5624
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 3605 5559 3663 5565
rect 3605 5525 3617 5559
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 4246 5556 4252 5568
rect 4019 5528 4252 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 6270 5516 6276 5568
rect 6328 5516 6334 5568
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 8662 5556 8668 5568
rect 8527 5528 8668 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8812 5528 9045 5556
rect 8812 5516 8818 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 9033 5519 9091 5525
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1578 5312 1584 5364
rect 1636 5312 1642 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3786 5352 3792 5364
rect 3099 5324 3792 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 5074 5312 5080 5364
rect 5132 5312 5138 5364
rect 8938 5312 8944 5364
rect 8996 5352 9002 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8996 5324 9137 5352
rect 8996 5312 9002 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 9125 5315 9183 5321
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 9916 5324 10425 5352
rect 9916 5312 9922 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1596 5216 1624 5312
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 7742 5284 7748 5296
rect 4387 5256 7748 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 7742 5244 7748 5256
rect 7800 5284 7806 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7800 5256 7849 5284
rect 7800 5244 7806 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 7837 5247 7895 5253
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1596 5188 1777 5216
rect 1397 5179 1455 5185
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4304 5188 4629 5216
rect 4304 5176 4310 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5721 5179 5779 5185
rect 5920 5188 6009 5216
rect 4172 5148 4200 5176
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 4172 5120 4445 5148
rect 4433 5117 4445 5120
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 5368 5080 5396 5179
rect 4120 5052 5396 5080
rect 4120 5040 4126 5052
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 3142 5012 3148 5024
rect 1995 4984 3148 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 5166 4972 5172 5024
rect 5224 4972 5230 5024
rect 5736 5012 5764 5179
rect 5920 5089 5948 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6236 5188 6469 5216
rect 6236 5176 6242 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 7466 5216 7472 5228
rect 7331 5188 7472 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 7576 5188 9781 5216
rect 6270 5108 6276 5160
rect 6328 5148 6334 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6328 5120 7113 5148
rect 6328 5108 6334 5120
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7576 5148 7604 5188
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 7101 5111 7159 5117
rect 7484 5120 7604 5148
rect 7745 5151 7803 5157
rect 7484 5092 7512 5120
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8018 5148 8024 5160
rect 7791 5120 8024 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 10244 5148 10272 5179
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10244 5120 10824 5148
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5049 5963 5083
rect 6549 5083 6607 5089
rect 5905 5043 5963 5049
rect 6012 5052 6316 5080
rect 6012 5012 6040 5052
rect 5736 4984 6040 5012
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 6288 5012 6316 5052
rect 6549 5049 6561 5083
rect 6595 5080 6607 5083
rect 7374 5080 7380 5092
rect 6595 5052 7380 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 7374 5040 7380 5052
rect 7432 5040 7438 5092
rect 7466 5040 7472 5092
rect 7524 5040 7530 5092
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 7616 5052 10057 5080
rect 7616 5040 7622 5052
rect 10045 5049 10057 5052
rect 10091 5049 10103 5083
rect 10045 5043 10103 5049
rect 10796 5024 10824 5120
rect 6730 5012 6736 5024
rect 6288 4984 6736 5012
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 6822 4972 6828 5024
rect 6880 4972 6886 5024
rect 9950 4972 9956 5024
rect 10008 4972 10014 5024
rect 10778 4972 10784 5024
rect 10836 4972 10842 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 4982 4808 4988 4820
rect 4479 4780 4988 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 6178 4768 6184 4820
rect 6236 4768 6242 4820
rect 6822 4768 6828 4820
rect 6880 4768 6886 4820
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 8018 4808 8024 4820
rect 7699 4780 8024 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3375 4712 4844 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 4816 4681 4844 4712
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3559 4644 3985 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 3973 4635 4031 4641
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4641 4859 4675
rect 6196 4672 6224 4768
rect 6840 4740 6868 4768
rect 6840 4712 7972 4740
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 6196 4644 6469 4672
rect 4801 4635 4859 4641
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 6972 4644 7205 4672
rect 6972 4632 6978 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7944 4681 7972 4712
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 9824 4712 10057 4740
rect 9824 4700 9830 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7432 4644 7757 4672
rect 7432 4632 7438 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9398 4672 9404 4684
rect 8435 4644 9404 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 9398 4632 9404 4644
rect 9456 4672 9462 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9456 4644 9689 4672
rect 9456 4632 9462 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3694 4604 3700 4616
rect 3651 4576 3700 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 3160 4536 3188 4567
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 7668 4576 8677 4604
rect 4154 4536 4160 4548
rect 3160 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 6748 4536 6776 4564
rect 7668 4536 7696 4576
rect 8665 4573 8677 4576
rect 8711 4604 8723 4607
rect 8754 4604 8760 4616
rect 8711 4576 8760 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8754 4564 8760 4576
rect 8812 4604 8818 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 8812 4576 9505 4604
rect 8812 4564 8818 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 6748 4508 7696 4536
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8573 4539 8631 4545
rect 8573 4536 8585 4539
rect 7800 4508 8585 4536
rect 7800 4496 7806 4508
rect 8573 4505 8585 4508
rect 8619 4505 8631 4539
rect 8573 4499 8631 4505
rect 9122 4496 9128 4548
rect 9180 4536 9186 4548
rect 9876 4536 9904 4567
rect 9180 4508 9904 4536
rect 9180 4496 9186 4508
rect 6914 4428 6920 4480
rect 6972 4428 6978 4480
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 7984 4440 8953 4468
rect 7984 4428 7990 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 8941 4431 8999 4437
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 3878 4224 3884 4276
rect 3936 4224 3942 4276
rect 4154 4224 4160 4276
rect 4212 4224 4218 4276
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 4614 4264 4620 4276
rect 4571 4236 4620 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6822 4264 6828 4276
rect 6236 4236 6828 4264
rect 6236 4224 6242 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7193 4267 7251 4273
rect 7193 4264 7205 4267
rect 6972 4236 7205 4264
rect 6972 4224 6978 4236
rect 7193 4233 7205 4236
rect 7239 4233 7251 4267
rect 9950 4264 9956 4276
rect 7193 4227 7251 4233
rect 9876 4236 9956 4264
rect 3896 4196 3924 4224
rect 7208 4196 7236 4227
rect 9766 4196 9772 4208
rect 3896 4168 4108 4196
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 992 4100 1409 4128
rect 992 4088 998 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 4080 4128 4108 4168
rect 4448 4168 5948 4196
rect 7208 4168 7696 4196
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4080 4100 4353 4128
rect 1397 4091 1455 4097
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 1762 4060 1768 4072
rect 1596 4032 1768 4060
rect 1596 4001 1624 4032
rect 1762 4020 1768 4032
rect 1820 4060 1826 4072
rect 4448 4060 4476 4168
rect 5920 4137 5948 4168
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4663 4100 4905 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4128 6055 4131
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6043 4100 6561 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 6549 4097 6561 4100
rect 6595 4128 6607 4131
rect 7006 4128 7012 4140
rect 6595 4100 7012 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 1820 4032 4476 4060
rect 1820 4020 1826 4032
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3961 1639 3995
rect 1581 3955 1639 3961
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 4709 3995 4767 4001
rect 4709 3992 4721 3995
rect 1912 3964 4721 3992
rect 1912 3952 1918 3964
rect 4709 3961 4721 3964
rect 4755 3961 4767 3995
rect 4709 3955 4767 3961
rect 4908 3924 4936 4091
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7668 4137 7696 4168
rect 9600 4168 9772 4196
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8570 4128 8576 4140
rect 8435 4100 8576 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 9306 4128 9312 4140
rect 8711 4100 9312 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9600 4137 9628 4168
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 9876 4205 9904 4236
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 9861 4199 9919 4205
rect 9861 4165 9873 4199
rect 9907 4165 9919 4199
rect 9861 4159 9919 4165
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9585 4091 9643 4097
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4060 6791 4063
rect 7760 4060 7788 4088
rect 6779 4032 7788 4060
rect 7837 4063 7895 4069
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 7469 3995 7527 4001
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 7852 3992 7880 4023
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8812 4032 8953 4060
rect 8812 4020 8818 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 7515 3964 7880 3992
rect 8849 3995 8907 4001
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 9140 3992 9168 4023
rect 8895 3964 9168 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 10318 3952 10324 4004
rect 10376 3952 10382 4004
rect 7374 3924 7380 3936
rect 4908 3896 7380 3924
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 8294 3884 8300 3936
rect 8352 3884 8358 3936
rect 8573 3927 8631 3933
rect 8573 3893 8585 3927
rect 8619 3924 8631 3927
rect 9030 3924 9036 3936
rect 8619 3896 9036 3924
rect 8619 3893 8631 3896
rect 8573 3887 8631 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3786 3720 3792 3732
rect 3099 3692 3792 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5583 3692 5917 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5905 3689 5917 3692
rect 5951 3720 5963 3723
rect 5951 3692 7880 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 6362 3544 6368 3596
rect 6420 3544 6426 3596
rect 7852 3593 7880 3692
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8662 3720 8668 3732
rect 8352 3692 8668 3720
rect 8352 3680 8358 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 8754 3680 8760 3732
rect 8812 3680 8818 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 10100 3692 10333 3720
rect 10100 3680 10106 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10321 3683 10379 3689
rect 8772 3593 8800 3680
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3553 8815 3587
rect 8757 3547 8815 3553
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2590 3516 2596 3528
rect 1636 3488 2596 3516
rect 1636 3476 1642 3488
rect 2590 3476 2596 3488
rect 2648 3516 2654 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2648 3488 2697 3516
rect 2648 3476 2654 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 2976 3448 3004 3479
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5626 3516 5632 3528
rect 5123 3488 5632 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6178 3516 6184 3528
rect 6135 3488 6184 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6270 3476 6276 3528
rect 6328 3476 6334 3528
rect 6632 3519 6690 3525
rect 6632 3485 6644 3519
rect 6678 3516 6690 3519
rect 7926 3516 7932 3528
rect 6678 3488 7932 3516
rect 6678 3485 6690 3488
rect 6632 3479 6690 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 2516 3420 3004 3448
rect 2516 3392 2544 3420
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 9214 3457 9220 3460
rect 5592 3420 7880 3448
rect 5592 3408 5598 3420
rect 7852 3392 7880 3420
rect 9208 3411 9220 3457
rect 9214 3408 9220 3411
rect 9272 3408 9278 3460
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 2866 3340 2872 3392
rect 2924 3340 2930 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 7466 3380 7472 3392
rect 5500 3352 7472 3380
rect 5500 3340 5506 3352
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 7834 3340 7840 3392
rect 7892 3340 7898 3392
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 10042 3380 10048 3392
rect 7984 3352 10048 3380
rect 7984 3340 7990 3352
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1762 3136 1768 3188
rect 1820 3136 1826 3188
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4948 3148 5273 3176
rect 4948 3136 4954 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 5810 3176 5816 3188
rect 5684 3148 5816 3176
rect 5684 3136 5690 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6178 3176 6184 3188
rect 5951 3148 6184 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6733 3179 6791 3185
rect 6733 3176 6745 3179
rect 6328 3148 6745 3176
rect 6328 3136 6334 3148
rect 6733 3145 6745 3148
rect 6779 3145 6791 3179
rect 6733 3139 6791 3145
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 7926 3136 7932 3188
rect 7984 3136 7990 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 8076 3148 8125 3176
rect 8076 3136 8082 3148
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 8113 3139 8171 3145
rect 9125 3179 9183 3185
rect 9125 3145 9137 3179
rect 9171 3176 9183 3179
rect 9214 3176 9220 3188
rect 9171 3148 9220 3176
rect 9171 3145 9183 3148
rect 9125 3139 9183 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 1394 3000 1400 3052
rect 1452 3000 1458 3052
rect 1780 3049 1808 3136
rect 5552 3108 5580 3136
rect 5092 3080 5580 3108
rect 5644 3080 6868 3108
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 5092 3049 5120 3080
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3040 5503 3043
rect 5644 3040 5672 3080
rect 5491 3012 5672 3040
rect 5721 3043 5779 3049
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 6181 3043 6239 3049
rect 5767 3012 6040 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 2516 2972 2544 3000
rect 1596 2944 2544 2972
rect 2608 2972 2636 3000
rect 5184 2972 5212 3003
rect 2608 2944 5212 2972
rect 6012 2972 6040 3012
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6227 3012 6561 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6564 2972 6592 3003
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 6730 2972 6736 2984
rect 6012 2944 6408 2972
rect 6564 2944 6736 2972
rect 1596 2913 1624 2944
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2873 1639 2907
rect 1581 2867 1639 2873
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 2317 2907 2375 2913
rect 2317 2904 2329 2907
rect 1912 2876 2329 2904
rect 1912 2864 1918 2876
rect 2317 2873 2329 2876
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 2746 2876 5764 2904
rect 1946 2796 1952 2848
rect 2004 2796 2010 2848
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2746 2836 2774 2876
rect 2271 2808 2774 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 4893 2839 4951 2845
rect 4893 2836 4905 2839
rect 4580 2808 4905 2836
rect 4580 2796 4586 2808
rect 4893 2805 4905 2808
rect 4939 2805 4951 2839
rect 4893 2799 4951 2805
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5500 2808 5641 2836
rect 5500 2796 5506 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 5736 2836 5764 2876
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6380 2913 6408 2944
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 6840 2972 6868 3080
rect 6932 3049 6960 3136
rect 7944 3108 7972 3136
rect 7484 3080 7972 3108
rect 8128 3080 9444 3108
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7484 2972 7512 3080
rect 8128 3052 8156 3080
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7742 3040 7748 3052
rect 7699 3012 7748 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 6840 2944 7512 2972
rect 6089 2907 6147 2913
rect 6089 2904 6101 2907
rect 5868 2876 6101 2904
rect 5868 2864 5874 2876
rect 6089 2873 6101 2876
rect 6135 2873 6147 2907
rect 6089 2867 6147 2873
rect 6365 2907 6423 2913
rect 6365 2873 6377 2907
rect 6411 2873 6423 2907
rect 6365 2867 6423 2873
rect 6472 2876 7512 2904
rect 6472 2836 6500 2876
rect 7484 2848 7512 2876
rect 5736 2808 6500 2836
rect 5629 2799 5687 2805
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7101 2839 7159 2845
rect 7101 2836 7113 2839
rect 6972 2808 7113 2836
rect 6972 2796 6978 2808
rect 7101 2805 7113 2808
rect 7147 2805 7159 2839
rect 7101 2799 7159 2805
rect 7466 2796 7472 2848
rect 7524 2796 7530 2848
rect 7668 2836 7696 3003
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 7852 3012 7941 3040
rect 7852 2913 7880 3012
rect 7929 3009 7941 3012
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 8110 3000 8116 3052
rect 8168 3000 8174 3052
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8251 3012 8285 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8220 2972 8248 3003
rect 8662 3000 8668 3052
rect 8720 3000 8726 3052
rect 9416 3049 9444 3080
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9861 3111 9919 3117
rect 9861 3108 9873 3111
rect 9640 3080 9873 3108
rect 9640 3068 9646 3080
rect 9861 3077 9873 3080
rect 9907 3077 9919 3111
rect 10336 3108 10364 3136
rect 10413 3111 10471 3117
rect 10413 3108 10425 3111
rect 10336 3080 10425 3108
rect 9861 3071 9919 3077
rect 10413 3077 10425 3080
rect 10459 3077 10471 3111
rect 10413 3071 10471 3077
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8220 2944 8493 2972
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2873 7895 2907
rect 7837 2867 7895 2873
rect 8220 2836 8248 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8680 2972 8708 3000
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 8680 2944 9781 2972
rect 8481 2935 8539 2941
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 10134 2932 10140 2984
rect 10192 2932 10198 2984
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 9122 2904 9128 2916
rect 8343 2876 9128 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 9122 2864 9128 2876
rect 9180 2864 9186 2916
rect 9585 2907 9643 2913
rect 9585 2873 9597 2907
rect 9631 2904 9643 2907
rect 10152 2904 10180 2932
rect 9631 2876 10180 2904
rect 9631 2873 9643 2876
rect 9585 2867 9643 2873
rect 9858 2836 9864 2848
rect 7668 2808 9864 2836
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 6454 2632 6460 2644
rect 3292 2604 6460 2632
rect 3292 2592 3298 2604
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7484 2604 9260 2632
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 5721 2567 5779 2573
rect 5721 2564 5733 2567
rect 5592 2536 5733 2564
rect 5592 2524 5598 2536
rect 5721 2533 5733 2536
rect 5767 2533 5779 2567
rect 7374 2564 7380 2576
rect 5721 2527 5779 2533
rect 5920 2536 7380 2564
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 1854 2428 1860 2440
rect 1811 2400 1860 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 2004 2400 2053 2428
rect 2004 2388 2010 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2924 2400 3065 2428
rect 2924 2388 2930 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3200 2400 4077 2428
rect 3200 2388 3206 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5224 2400 5365 2428
rect 5224 2388 5230 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 842 2320 848 2372
rect 900 2360 906 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 900 2332 1409 2360
rect 900 2320 906 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 4982 2320 4988 2372
rect 5040 2320 5046 2372
rect 5736 2360 5764 2527
rect 5920 2437 5948 2536
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 7484 2496 7512 2604
rect 7926 2564 7932 2576
rect 6196 2468 7512 2496
rect 7760 2536 7932 2564
rect 6196 2437 6224 2468
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6454 2388 6460 2440
rect 6512 2388 6518 2440
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6972 2400 7113 2428
rect 6972 2388 6978 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 7760 2437 7788 2536
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9122 2564 9128 2576
rect 8619 2536 9128 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 9232 2564 9260 2604
rect 9306 2592 9312 2644
rect 9364 2632 9370 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9364 2604 9597 2632
rect 9364 2592 9370 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 10042 2564 10048 2576
rect 9232 2536 10048 2564
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 9398 2496 9404 2508
rect 7883 2468 9404 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9769 2431 9827 2437
rect 8803 2400 9720 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 6638 2360 6644 2372
rect 5736 2332 6644 2360
rect 6638 2320 6644 2332
rect 6696 2320 6702 2372
rect 7484 2360 7512 2388
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7484 2332 8125 2360
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 9122 2320 9128 2372
rect 9180 2320 9186 2372
rect 9692 2360 9720 2400
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9858 2428 9864 2440
rect 9815 2400 9864 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10042 2360 10048 2372
rect 9692 2332 10048 2360
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 10134 2320 10140 2372
rect 10192 2320 10198 2372
rect 1854 2252 1860 2304
rect 1912 2292 1918 2304
rect 2133 2295 2191 2301
rect 2133 2292 2145 2295
rect 1912 2264 2145 2292
rect 1912 2252 1918 2264
rect 2133 2261 2145 2264
rect 2179 2261 2191 2295
rect 2133 2255 2191 2261
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 3145 2295 3203 2301
rect 3145 2292 3157 2295
rect 2924 2264 3157 2292
rect 2924 2252 2930 2264
rect 3145 2261 3157 2264
rect 3191 2261 3203 2295
rect 3145 2255 3203 2261
rect 4154 2252 4160 2304
rect 4212 2252 4218 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 6362 2292 6368 2304
rect 6135 2264 6368 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 6362 2252 6368 2264
rect 6420 2252 6426 2304
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 6972 2264 7205 2292
rect 6972 2252 6978 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 7984 2264 8217 2292
rect 7984 2252 7990 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8996 2264 9229 2292
rect 8996 2252 9002 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10229 2295 10287 2301
rect 10229 2292 10241 2295
rect 10008 2264 10241 2292
rect 10008 2252 10014 2264
rect 10229 2261 10241 2264
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 6362 2048 6368 2100
rect 6420 2088 6426 2100
rect 10134 2088 10140 2100
rect 6420 2060 10140 2088
rect 6420 2048 6426 2060
rect 10134 2048 10140 2060
rect 10192 2048 10198 2100
rect 9122 2020 9128 2032
rect 6886 1992 9128 2020
rect 5258 1844 5264 1896
rect 5316 1884 5322 1896
rect 6886 1884 6914 1992
rect 9122 1980 9128 1992
rect 9180 1980 9186 2032
rect 5316 1856 6914 1884
rect 5316 1844 5322 1856
rect 5902 1368 5908 1420
rect 5960 1408 5966 1420
rect 6546 1408 6552 1420
rect 5960 1380 6552 1408
rect 5960 1368 5966 1380
rect 6546 1368 6552 1380
rect 6604 1368 6610 1420
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 848 9596 900 9648
rect 1860 9596 1912 9648
rect 2872 9596 2924 9648
rect 3884 9596 3936 9648
rect 4896 9596 4948 9648
rect 6184 9596 6236 9648
rect 6920 9596 6972 9648
rect 7932 9596 7984 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 9588 9664 9640 9716
rect 8944 9596 8996 9648
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10600 9528 10652 9580
rect 8944 9460 8996 9512
rect 9956 9392 10008 9444
rect 9036 9324 9088 9376
rect 9220 9324 9272 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 7380 9120 7432 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 9220 9120 9272 9172
rect 9312 9120 9364 9172
rect 940 8916 992 8968
rect 2780 8984 2832 9036
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 5632 9052 5684 9104
rect 10140 9052 10192 9104
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 11060 8916 11112 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 10048 8848 10100 8900
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2136 8780 2188 8789
rect 5264 8780 5316 8832
rect 5540 8780 5592 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 6920 8780 6972 8832
rect 8668 8780 8720 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 6460 8576 6512 8628
rect 6736 8576 6788 8628
rect 8944 8576 8996 8628
rect 1584 8508 1636 8560
rect 6276 8508 6328 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 5172 8440 5224 8492
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 6552 8440 6604 8492
rect 9312 8440 9364 8492
rect 5632 8372 5684 8424
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 3792 8304 3844 8356
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 8668 8304 8720 8356
rect 10140 8440 10192 8492
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 5632 8032 5684 8084
rect 6644 8032 6696 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8300 8032 8352 8084
rect 4436 7896 4488 7948
rect 5172 7896 5224 7948
rect 5540 7964 5592 8016
rect 6920 7896 6972 7948
rect 5172 7692 5224 7744
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9036 7828 9088 7880
rect 7840 7692 7892 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 6644 7488 6696 7540
rect 6736 7488 6788 7540
rect 9864 7488 9916 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 3792 7352 3844 7404
rect 5080 7395 5132 7404
rect 5080 7361 5114 7395
rect 5114 7361 5132 7395
rect 5080 7352 5132 7361
rect 5908 7352 5960 7404
rect 4068 7148 4120 7200
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 8024 7284 8076 7336
rect 9864 7284 9916 7336
rect 5448 7148 5500 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 6920 7148 6972 7200
rect 9404 7148 9456 7200
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 5080 6944 5132 6996
rect 9404 6987 9456 6996
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 5172 6919 5224 6928
rect 5172 6885 5181 6919
rect 5181 6885 5215 6919
rect 5215 6885 5224 6919
rect 5172 6876 5224 6885
rect 5908 6876 5960 6928
rect 5540 6808 5592 6860
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 7656 6808 7708 6860
rect 3792 6740 3844 6749
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 6460 6740 6512 6792
rect 6920 6740 6972 6792
rect 5632 6604 5684 6656
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10876 6808 10928 6860
rect 7748 6604 7800 6613
rect 8116 6604 8168 6656
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9680 6604 9732 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 2504 6400 2556 6452
rect 5632 6400 5684 6452
rect 5724 6400 5776 6452
rect 6184 6400 6236 6452
rect 940 6264 992 6316
rect 5448 6332 5500 6384
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4068 6196 4120 6248
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5080 6196 5132 6205
rect 7748 6400 7800 6452
rect 8668 6400 8720 6452
rect 9128 6400 9180 6452
rect 9772 6400 9824 6452
rect 8116 6332 8168 6384
rect 8944 6264 8996 6316
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 7472 6128 7524 6180
rect 9680 6196 9732 6248
rect 10324 6196 10376 6248
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 4160 6060 4212 6112
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 4344 6060 4396 6112
rect 4988 6060 5040 6112
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 5816 6060 5868 6112
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 10232 6060 10284 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 4252 5856 4304 5908
rect 4344 5856 4396 5908
rect 4988 5856 5040 5908
rect 5356 5856 5408 5908
rect 6552 5856 6604 5908
rect 5724 5788 5776 5840
rect 8944 5788 8996 5840
rect 3884 5695 3936 5704
rect 3884 5661 3893 5695
rect 3893 5661 3927 5695
rect 3927 5661 3936 5695
rect 3884 5652 3936 5661
rect 4252 5652 4304 5704
rect 4988 5652 5040 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 7564 5720 7616 5772
rect 5816 5652 5868 5661
rect 5080 5584 5132 5636
rect 5448 5584 5500 5636
rect 6460 5627 6512 5636
rect 6460 5593 6469 5627
rect 6469 5593 6503 5627
rect 6503 5593 6512 5627
rect 6460 5584 6512 5593
rect 8852 5584 8904 5636
rect 10232 5584 10284 5636
rect 4252 5516 4304 5568
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8668 5516 8720 5568
rect 8760 5516 8812 5568
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 1584 5312 1636 5364
rect 3792 5312 3844 5364
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 8944 5312 8996 5364
rect 9864 5312 9916 5364
rect 940 5176 992 5228
rect 7748 5244 7800 5296
rect 4160 5176 4212 5228
rect 4252 5176 4304 5228
rect 4068 5040 4120 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 3148 4972 3200 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 6184 5176 6236 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7472 5176 7524 5228
rect 6276 5108 6328 5160
rect 8024 5108 8076 5160
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 7380 5040 7432 5092
rect 7472 5040 7524 5092
rect 7564 5040 7616 5092
rect 6736 4972 6788 5024
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 10784 4972 10836 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 6184 4768 6236 4820
rect 6828 4768 6880 4820
rect 8024 4768 8076 4820
rect 6920 4632 6972 4684
rect 7380 4632 7432 4684
rect 9772 4700 9824 4752
rect 9404 4632 9456 4684
rect 3700 4564 3752 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 6736 4564 6788 4616
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 4160 4496 4212 4548
rect 8760 4564 8812 4616
rect 7748 4496 7800 4548
rect 9128 4496 9180 4548
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 7932 4428 7984 4480
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 3884 4224 3936 4276
rect 4160 4267 4212 4276
rect 4160 4233 4169 4267
rect 4169 4233 4203 4267
rect 4203 4233 4212 4267
rect 4160 4224 4212 4233
rect 4620 4224 4672 4276
rect 6184 4224 6236 4276
rect 6828 4224 6880 4276
rect 6920 4224 6972 4276
rect 9772 4199 9824 4208
rect 940 4088 992 4140
rect 1768 4020 1820 4072
rect 1860 3952 1912 4004
rect 7012 4088 7064 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7748 4088 7800 4140
rect 8576 4088 8628 4140
rect 9312 4088 9364 4140
rect 9772 4165 9781 4199
rect 9781 4165 9815 4199
rect 9815 4165 9824 4199
rect 9772 4156 9824 4165
rect 9956 4224 10008 4276
rect 8760 4020 8812 4072
rect 10324 3995 10376 4004
rect 10324 3961 10333 3995
rect 10333 3961 10367 3995
rect 10367 3961 10376 3995
rect 10324 3952 10376 3961
rect 7380 3884 7432 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8300 3884 8352 3893
rect 9036 3884 9088 3936
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 3792 3680 3844 3732
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 8668 3680 8720 3732
rect 8760 3680 8812 3732
rect 10048 3680 10100 3732
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 1584 3476 1636 3528
rect 2596 3476 2648 3528
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 5632 3476 5684 3528
rect 6184 3476 6236 3528
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 7932 3476 7984 3528
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 5540 3408 5592 3460
rect 9220 3451 9272 3460
rect 9220 3417 9254 3451
rect 9254 3417 9272 3451
rect 9220 3408 9272 3417
rect 2504 3340 2556 3392
rect 2872 3383 2924 3392
rect 2872 3349 2881 3383
rect 2881 3349 2915 3383
rect 2915 3349 2924 3383
rect 2872 3340 2924 3349
rect 5448 3340 5500 3392
rect 7472 3340 7524 3392
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 7840 3340 7892 3392
rect 7932 3340 7984 3392
rect 10048 3340 10100 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 1768 3136 1820 3188
rect 4896 3136 4948 3188
rect 5540 3136 5592 3188
rect 5632 3136 5684 3188
rect 5816 3136 5868 3188
rect 6184 3136 6236 3188
rect 6276 3136 6328 3188
rect 6920 3136 6972 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 7932 3136 7984 3188
rect 8024 3136 8076 3188
rect 9220 3136 9272 3188
rect 10324 3136 10376 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2596 3000 2648 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 1860 2864 1912 2916
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 4528 2796 4580 2848
rect 5448 2796 5500 2848
rect 5816 2864 5868 2916
rect 6736 2932 6788 2984
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 6920 2796 6972 2848
rect 7472 2796 7524 2848
rect 7748 3000 7800 3052
rect 8116 3000 8168 3052
rect 8668 3000 8720 3052
rect 9588 3068 9640 3120
rect 10140 2932 10192 2984
rect 9128 2864 9180 2916
rect 9864 2796 9916 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 3240 2592 3292 2644
rect 6460 2592 6512 2644
rect 5540 2524 5592 2576
rect 1860 2388 1912 2440
rect 1952 2388 2004 2440
rect 2872 2388 2924 2440
rect 3148 2388 3200 2440
rect 5172 2388 5224 2440
rect 848 2320 900 2372
rect 4988 2363 5040 2372
rect 4988 2329 4997 2363
rect 4997 2329 5031 2363
rect 5031 2329 5040 2363
rect 4988 2320 5040 2329
rect 7380 2524 7432 2576
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 6920 2388 6972 2440
rect 7472 2388 7524 2440
rect 7932 2524 7984 2576
rect 9128 2524 9180 2576
rect 9312 2592 9364 2644
rect 10048 2524 10100 2576
rect 9404 2456 9456 2508
rect 6644 2320 6696 2372
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 9864 2388 9916 2440
rect 10048 2320 10100 2372
rect 10140 2363 10192 2372
rect 10140 2329 10149 2363
rect 10149 2329 10183 2363
rect 10183 2329 10192 2363
rect 10140 2320 10192 2329
rect 1860 2252 1912 2304
rect 2872 2252 2924 2304
rect 4160 2295 4212 2304
rect 4160 2261 4169 2295
rect 4169 2261 4203 2295
rect 4203 2261 4212 2295
rect 4160 2252 4212 2261
rect 6368 2252 6420 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6920 2252 6972 2304
rect 7932 2252 7984 2304
rect 8944 2252 8996 2304
rect 9956 2252 10008 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 6368 2048 6420 2100
rect 10140 2048 10192 2100
rect 5264 1844 5316 1896
rect 9128 1980 9180 2032
rect 5908 1368 5960 1420
rect 6552 1368 6604 1420
<< metal2 >>
rect 846 11200 902 12000
rect 1858 11200 1914 12000
rect 2870 11200 2926 12000
rect 3882 11200 3938 12000
rect 4894 11200 4950 12000
rect 5906 11200 5962 12000
rect 6012 11206 6224 11234
rect 860 9654 888 11200
rect 1872 9654 1900 11200
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 1950 9752 2006 9761
rect 1950 9687 2006 9696
rect 848 9648 900 9654
rect 848 9590 900 9596
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 952 8974 980 9007
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8566 1624 8774
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 1780 6914 1808 9522
rect 1964 8974 1992 9687
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9466 2360 9522
rect 2332 9438 2544 9466
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 2136 8832 2188 8838
rect 2056 8792 2136 8820
rect 1398 6896 1454 6905
rect 1780 6886 1900 6914
rect 1398 6831 1454 6840
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 5817 980 6258
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 938 5808 994 5817
rect 938 5743 994 5752
rect 1596 5370 1624 6054
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4729 980 5170
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3641 980 4082
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 1596 3534 1624 4966
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1780 3194 1808 4014
rect 1872 4010 1900 6886
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 2056 3058 2084 8792
rect 2136 8774 2188 8780
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2516 6458 2544 9438
rect 2792 9042 2820 10911
rect 2884 9654 2912 11200
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3896 9654 3924 11200
rect 4908 9654 4936 11200
rect 5920 11098 5948 11200
rect 6012 11098 6040 11206
rect 5920 11070 6040 11098
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6196 9654 6224 11206
rect 6918 11200 6974 12000
rect 7930 11200 7986 12000
rect 8942 11200 8998 12000
rect 9310 11248 9366 11257
rect 6932 9654 6960 11200
rect 7944 9654 7972 11200
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8956 9654 8984 11200
rect 9954 11200 10010 12000
rect 10966 11200 11022 12000
rect 9310 11183 9366 11192
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 3344 9178 3372 9522
rect 4356 9178 4384 9522
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3804 7410 3832 8298
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3804 5370 3832 6734
rect 4080 6254 4108 7142
rect 4448 6322 4476 7890
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 3058 2544 3334
rect 2608 3058 2636 3470
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1412 2689 1440 2994
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1398 2680 1454 2689
rect 1398 2615 1454 2624
rect 1872 2446 1900 2858
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1964 2446 1992 2790
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2884 2446 2912 3334
rect 3160 2446 3188 4966
rect 3896 4706 3924 5646
rect 4080 5098 4108 6190
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4172 5234 4200 6054
rect 4264 5914 4292 6054
rect 4356 5914 4384 6054
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4448 5794 4476 6258
rect 4264 5766 4476 5794
rect 4264 5710 4292 5766
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5234 4292 5510
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3712 4678 3924 4706
rect 3712 4622 3740 4678
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3804 3738 3832 4558
rect 3896 4282 3924 4678
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4172 4282 4200 4490
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 4540 2854 4568 8910
rect 4908 8634 4936 8910
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 5184 7954 5212 8434
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5092 7002 5120 7346
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5184 6934 5212 7686
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5000 5914 5028 6054
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 5000 4826 5028 5646
rect 5092 5642 5120 6190
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 5092 5370 5120 5578
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4632 4282 4660 4558
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4908 3194 4936 3470
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 848 2372 900 2378
rect 848 2314 900 2320
rect 860 800 888 2314
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 1872 800 1900 2246
rect 2884 800 2912 2246
rect 3252 1465 3280 2586
rect 5184 2446 5212 4966
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4160 2304 4212 2310
rect 3896 2264 4160 2292
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3896 800 3924 2264
rect 4160 2246 4212 2252
rect 5000 1170 5028 2314
rect 5276 1902 5304 8774
rect 5368 5914 5396 9522
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8498 5580 8774
rect 5644 8514 5672 9046
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 6472 8634 6500 8774
rect 6748 8634 6776 9522
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7392 9178 7420 9522
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6276 8560 6328 8566
rect 5540 8492 5592 8498
rect 5644 8486 5764 8514
rect 6276 8502 6328 8508
rect 5540 8434 5592 8440
rect 5552 8022 5580 8434
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5644 8090 5672 8366
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6882 5488 7142
rect 5736 6882 5764 8486
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6934 5948 7346
rect 5460 6866 5580 6882
rect 5460 6860 5592 6866
rect 5460 6854 5540 6860
rect 5540 6802 5592 6808
rect 5644 6854 5764 6882
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5644 6746 5672 6854
rect 5920 6798 5948 6870
rect 5908 6792 5960 6798
rect 5552 6718 5672 6746
rect 5736 6740 5908 6746
rect 5736 6734 5960 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5736 6718 5948 6734
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5460 5642 5488 6326
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5552 3618 5580 6718
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 6458 5672 6598
rect 5736 6458 5764 6718
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 6196 6458 6224 6734
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5736 5846 5764 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5828 5710 5856 6054
rect 5816 5704 5868 5710
rect 6288 5658 6316 8502
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6798 6500 7142
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 5816 5646 5868 5652
rect 6196 5630 6316 5658
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6196 5234 6224 5630
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6196 5114 6224 5170
rect 6288 5166 6316 5510
rect 6104 5086 6224 5114
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6104 4570 6132 5086
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 4826 6224 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6288 4622 6316 5102
rect 6276 4616 6328 4622
rect 6104 4542 6224 4570
rect 6276 4558 6328 4564
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 6196 4282 6224 4542
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 5552 3590 5764 3618
rect 6380 3602 6408 6734
rect 6564 5914 6592 8434
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 8090 6684 8366
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6932 7954 6960 8774
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7576 8090 7604 8366
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6748 7546 6776 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 2854 5488 3334
rect 5552 3194 5580 3402
rect 5644 3194 5672 3470
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5736 2774 5764 3590
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 6196 3194 6224 3470
rect 6288 3194 6316 3470
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 5828 2922 5856 3130
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5552 2746 5764 2774
rect 5552 2582 5580 2746
rect 6472 2650 6500 5578
rect 6656 4978 6684 7482
rect 7024 7342 7052 7822
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 6798 6960 7142
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7668 6866 7696 8910
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 8090 8340 8366
rect 8680 8362 8708 8774
rect 8956 8634 8984 9454
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 9048 7886 9076 9318
rect 9140 9178 9168 9522
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9178 9260 9318
rect 9324 9178 9352 11183
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9600 9722 9628 10095
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9968 9450 9996 11200
rect 10980 10010 11008 11200
rect 10980 9982 11100 10010
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 10152 9110 10180 9522
rect 10140 9104 10192 9110
rect 10612 9081 10640 9522
rect 10140 9046 10192 9052
rect 10598 9072 10654 9081
rect 10598 9007 10654 9016
rect 11072 8974 11100 9982
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9324 7993 9352 8434
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7342 7880 7686
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6458 7788 6598
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 5030 6776 5170
rect 6564 4950 6684 4978
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 6460 2440 6512 2446
rect 6564 2428 6592 4950
rect 6748 4622 6776 4966
rect 6840 4826 6868 4966
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6932 4690 6960 6054
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 7484 5234 7512 6122
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7576 5098 7604 5714
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5302 7788 5510
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 8036 5166 8064 7278
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8128 6390 8156 6598
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8680 6458 8708 6598
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8956 6322 8984 7822
rect 9876 7546 9904 8842
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 7002 9444 7142
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9140 6458 9168 6598
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5846 8984 6258
rect 9692 6254 9720 6598
rect 9784 6458 9812 6734
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 8944 5840 8996 5846
rect 8206 5808 8262 5817
rect 8128 5766 8206 5794
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7392 4690 7420 5034
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6512 2400 6592 2428
rect 6460 2382 6512 2388
rect 6656 2378 6684 2994
rect 6748 2990 6776 4558
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4282 6960 4422
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6840 4162 6868 4218
rect 6840 4134 6960 4162
rect 7024 4146 7052 4558
rect 6932 3194 6960 4134
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7392 3194 7420 3878
rect 7484 3398 7512 5034
rect 8036 4826 8064 5102
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7760 4146 7788 4490
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7576 3890 7604 4082
rect 7576 3862 7788 3890
rect 7760 3398 7788 3862
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7852 3398 7880 3567
rect 7944 3534 7972 4422
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7760 3058 7788 3334
rect 7944 3194 7972 3334
rect 8036 3194 8064 3470
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 6932 2446 6960 2790
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7380 2576 7432 2582
rect 7378 2544 7380 2553
rect 7432 2544 7434 2553
rect 7378 2479 7434 2488
rect 7484 2446 7512 2790
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6380 2106 6408 2246
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 6564 1426 6592 2246
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 6552 1420 6604 1426
rect 6552 1362 6604 1368
rect 4908 1142 5028 1170
rect 4908 800 4936 1142
rect 5920 800 5948 1362
rect 6932 800 6960 2246
rect 846 0 902 800
rect 1858 0 1914 800
rect 2870 0 2926 800
rect 3882 0 3938 800
rect 4894 0 4950 800
rect 5906 0 5962 800
rect 6918 0 6974 800
rect 7576 377 7604 2994
rect 7944 2582 7972 3130
rect 8128 3058 8156 5766
rect 8944 5782 8996 5788
rect 8206 5743 8262 5752
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8680 4162 8708 5510
rect 8772 4622 8800 5510
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8588 4146 8708 4162
rect 8576 4140 8708 4146
rect 8628 4134 8708 4140
rect 8576 4082 8628 4088
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3738 8340 3878
rect 8772 3738 8800 4014
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8680 3058 8708 3674
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8864 2774 8892 5578
rect 8956 5370 8984 5782
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8956 3602 8984 5306
rect 9048 3942 9076 6190
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 4690 9444 6054
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9876 5370 9904 7278
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9140 2922 9168 4490
rect 9784 4214 9812 4694
rect 9968 4282 9996 4966
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9232 3194 9260 3402
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 8864 2746 9168 2774
rect 9140 2582 9168 2746
rect 9324 2650 9352 4082
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 10060 3738 10088 8842
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3398 10088 3674
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9600 2938 9628 3062
rect 10152 2990 10180 8434
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10874 6896 10930 6905
rect 10874 6831 10876 6840
rect 10928 6831 10930 6840
rect 10876 6802 10928 6808
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5642 10272 6054
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10336 5234 10364 6190
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4729 10824 4966
rect 10782 4720 10838 4729
rect 10782 4655 10838 4664
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10336 3194 10364 3946
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 9416 2910 9628 2938
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9416 2514 9444 2910
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9876 2446 9904 2790
rect 10336 2774 10364 3130
rect 10060 2746 10364 2774
rect 10060 2582 10088 2746
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 7944 800 7972 2246
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8956 800 8984 2246
rect 9140 2038 9168 2314
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9968 800 9996 2246
rect 10060 1465 10088 2314
rect 10152 2106 10180 2314
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 10046 1456 10102 1465
rect 10046 1391 10102 1400
rect 7562 368 7618 377
rect 7562 303 7618 312
rect 7930 0 7986 800
rect 8942 0 8998 800
rect 9954 0 10010 800
<< via2 >>
rect 2778 10920 2834 10976
rect 1950 9696 2006 9752
rect 938 9016 994 9072
rect 1398 8200 1454 8256
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 1398 6840 1454 6896
rect 938 5752 994 5808
rect 938 4664 994 4720
rect 938 3576 994 3632
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 9310 11192 9366 11248
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 1398 2624 1454 2680
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 3238 1400 3294 1456
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 9586 10104 9642 10160
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10598 9016 10654 9072
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 9310 7928 9366 7984
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7838 3576 7894 3632
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 7378 2524 7380 2544
rect 7380 2524 7432 2544
rect 7432 2524 7434 2544
rect 7378 2488 7434 2524
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8206 5752 8262 5808
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10874 6860 10930 6896
rect 10874 6840 10876 6860
rect 10876 6840 10928 6860
rect 10928 6840 10930 6860
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10782 4664 10838 4720
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 10046 1400 10102 1456
rect 7562 312 7618 368
<< metal3 >>
rect 0 11250 800 11280
rect 9305 11250 9371 11253
rect 11200 11250 12000 11280
rect 0 11190 1042 11250
rect 0 11160 800 11190
rect 982 10978 1042 11190
rect 9305 11248 12000 11250
rect 9305 11192 9310 11248
rect 9366 11192 12000 11248
rect 9305 11190 12000 11192
rect 9305 11187 9371 11190
rect 11200 11160 12000 11190
rect 2773 10978 2839 10981
rect 982 10976 2839 10978
rect 982 10920 2778 10976
rect 2834 10920 2839 10976
rect 982 10918 2839 10920
rect 2773 10915 2839 10918
rect 0 10162 800 10192
rect 9581 10162 9647 10165
rect 11200 10162 12000 10192
rect 0 10102 1042 10162
rect 0 10072 800 10102
rect 982 9754 1042 10102
rect 9581 10160 12000 10162
rect 9581 10104 9586 10160
rect 9642 10104 12000 10160
rect 9581 10102 12000 10104
rect 9581 10099 9647 10102
rect 11200 10072 12000 10102
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 1945 9754 2011 9757
rect 982 9752 2011 9754
rect 982 9696 1950 9752
rect 2006 9696 2011 9752
rect 982 9694 2011 9696
rect 1945 9691 2011 9694
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 10593 9074 10659 9077
rect 11200 9074 12000 9104
rect 10593 9072 12000 9074
rect 10593 9016 10598 9072
rect 10654 9016 12000 9072
rect 10593 9014 12000 9016
rect 10593 9011 10659 9014
rect 11200 8984 12000 9014
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 1393 8256 1459 8261
rect 1393 8200 1398 8256
rect 1454 8200 1459 8256
rect 1393 8195 1459 8200
rect 0 7986 800 8016
rect 1396 7986 1456 8195
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7926 1456 7986
rect 9305 7986 9371 7989
rect 11200 7986 12000 8016
rect 9305 7984 12000 7986
rect 9305 7928 9310 7984
rect 9366 7928 12000 7984
rect 9305 7926 12000 7928
rect 0 7896 800 7926
rect 9305 7923 9371 7926
rect 11200 7896 12000 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 10869 6898 10935 6901
rect 11200 6898 12000 6928
rect 10869 6896 12000 6898
rect 10869 6840 10874 6896
rect 10930 6840 12000 6896
rect 10869 6838 12000 6840
rect 10869 6835 10935 6838
rect 11200 6808 12000 6838
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 8201 5810 8267 5813
rect 11200 5810 12000 5840
rect 8201 5808 12000 5810
rect 8201 5752 8206 5808
rect 8262 5752 12000 5808
rect 8201 5750 12000 5752
rect 8201 5747 8267 5750
rect 11200 5720 12000 5750
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 10777 4722 10843 4725
rect 11200 4722 12000 4752
rect 10777 4720 12000 4722
rect 10777 4664 10782 4720
rect 10838 4664 12000 4720
rect 10777 4662 12000 4664
rect 10777 4659 10843 4662
rect 11200 4632 12000 4662
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 7833 3634 7899 3637
rect 11200 3634 12000 3664
rect 7833 3632 12000 3634
rect 7833 3576 7838 3632
rect 7894 3576 12000 3632
rect 7833 3574 12000 3576
rect 7833 3571 7899 3574
rect 11200 3544 12000 3574
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 1393 2682 1459 2685
rect 798 2680 1459 2682
rect 798 2624 1398 2680
rect 1454 2624 1459 2680
rect 798 2622 1459 2624
rect 798 2576 858 2622
rect 1393 2619 1459 2622
rect 0 2486 858 2576
rect 7373 2546 7439 2549
rect 11200 2546 12000 2576
rect 7373 2544 12000 2546
rect 7373 2488 7378 2544
rect 7434 2488 12000 2544
rect 7373 2486 12000 2488
rect 0 2456 800 2486
rect 7373 2483 7439 2486
rect 11200 2456 12000 2486
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 0 1458 800 1488
rect 3233 1458 3299 1461
rect 0 1456 3299 1458
rect 0 1400 3238 1456
rect 3294 1400 3299 1456
rect 0 1398 3299 1400
rect 0 1368 800 1398
rect 3233 1395 3299 1398
rect 10041 1458 10107 1461
rect 11200 1458 12000 1488
rect 10041 1456 12000 1458
rect 10041 1400 10046 1456
rect 10102 1400 12000 1456
rect 10041 1398 12000 1400
rect 10041 1395 10107 1398
rect 11200 1368 12000 1398
rect 7557 370 7623 373
rect 11200 370 12000 400
rect 7557 368 12000 370
rect 7557 312 7562 368
rect 7618 312 12000 368
rect 7557 310 12000 312
rect 7557 307 7623 310
rect 11200 280 12000 310
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform -1 0 8740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform -1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform -1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform -1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform -1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1688980957
transform -1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform -1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1688980957
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform -1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1688980957
transform 1 0 4968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1688980957
transform -1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 5520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform -1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1688980957
transform -1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1688980957
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1688980957
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1688980957
transform -1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1688980957
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1688980957
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1688980957
transform 1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _102_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _103_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _104_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _107_
timestamp 1688980957
transform -1 0 10488 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 1688980957
transform -1 0 8832 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _122_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform -1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform -1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1688980957
transform -1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform -1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform -1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _131__42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _132_
timestamp 1688980957
transform 1 0 4600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _133_
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _134_
timestamp 1688980957
transform 1 0 4140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _135_
timestamp 1688980957
transform -1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _136_
timestamp 1688980957
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _137_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _138_
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _139_
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _140_
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _141_
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _142_
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _144_
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _144__43
timestamp 1688980957
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _145_
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _146_
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _147_
timestamp 1688980957
transform -1 0 6348 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _148_
timestamp 1688980957
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _149_
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _150_
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _151_
timestamp 1688980957
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _152_
timestamp 1688980957
transform 1 0 7728 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _153_
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _154_
timestamp 1688980957
transform 1 0 6532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _155__44
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _155_
timestamp 1688980957
transform -1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _156_
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _157_
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _158_
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_48
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_70
timestamp 1688980957
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_95
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_6
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_28
timestamp 1688980957
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_40
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_66
timestamp 1688980957
transform 1 0 7176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_88
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1688980957
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_101
timestamp 1688980957
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_30 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_50
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_67
timestamp 1688980957
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_102
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_46
timestamp 1688980957
transform 1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_54
timestamp 1688980957
transform 1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_10
timestamp 1688980957
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_47
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_64
timestamp 1688980957
transform 1 0 6992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_23
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_52
timestamp 1688980957
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_78
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_102
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_6
timestamp 1688980957
transform 1 0 1656 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_12
timestamp 1688980957
transform 1 0 2208 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_16
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_28
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_56
timestamp 1688980957
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_88
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1688980957
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_77
timestamp 1688980957
transform 1 0 8188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_89
timestamp 1688980957
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_62
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_67
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_74
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_102
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_43
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_66
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_84
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_12
timestamp 1688980957
transform 1 0 2208 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_38
timestamp 1688980957
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_50
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_61
timestamp 1688980957
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_70
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_74
timestamp 1688980957
transform 1 0 7912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 7912 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform -1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform -1 0 3496 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 5520 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 7544 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform -1 0 5520 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 6992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 9016 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
port 0 nsew signal tristate
flabel metal3 s 11200 10072 12000 10192 0 FreeSans 480 0 0 0 ccff_head
port 1 nsew signal input
flabel metal3 s 11200 11160 12000 11280 0 FreeSans 480 0 0 0 ccff_tail
port 2 nsew signal tristate
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 3 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 4 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 5 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 6 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 7 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 8 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 9 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 10 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 11 nsew signal input
flabel metal2 s 846 11200 902 12000 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 12 nsew signal tristate
flabel metal2 s 1858 11200 1914 12000 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 13 nsew signal tristate
flabel metal2 s 2870 11200 2926 12000 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 14 nsew signal tristate
flabel metal2 s 3882 11200 3938 12000 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 15 nsew signal tristate
flabel metal2 s 4894 11200 4950 12000 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 16 nsew signal tristate
flabel metal2 s 5906 11200 5962 12000 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 17 nsew signal tristate
flabel metal2 s 6918 11200 6974 12000 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 18 nsew signal tristate
flabel metal2 s 7930 11200 7986 12000 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 19 nsew signal tristate
flabel metal2 s 8942 11200 8998 12000 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 20 nsew signal tristate
flabel metal3 s 11200 280 12000 400 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 21 nsew signal input
flabel metal3 s 11200 1368 12000 1488 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 22 nsew signal input
flabel metal3 s 11200 2456 12000 2576 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 23 nsew signal input
flabel metal3 s 11200 3544 12000 3664 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 24 nsew signal input
flabel metal3 s 11200 4632 12000 4752 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 25 nsew signal input
flabel metal3 s 11200 5720 12000 5840 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 26 nsew signal input
flabel metal3 s 11200 6808 12000 6928 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 27 nsew signal input
flabel metal3 s 11200 7896 12000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 28 nsew signal input
flabel metal3 s 11200 8984 12000 9104 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 29 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 30 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 31 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 32 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 33 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 34 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 35 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 36 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 37 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 38 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 39 nsew signal input
flabel metal2 s 9954 11200 10010 12000 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 40 nsew signal tristate
flabel metal2 s 10966 11200 11022 12000 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 41 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 5520 7854 5520 7854 0 _000_
rlabel metal2 4186 4386 4186 4386 0 _001_
rlabel metal1 7360 7514 7360 7514 0 _002_
rlabel metal1 6578 6324 6578 6324 0 _003_
rlabel metal1 9844 6290 9844 6290 0 _004_
rlabel metal1 5980 5202 5980 5202 0 _005_
rlabel metal1 7912 3026 7912 3026 0 _006_
rlabel metal1 5888 3026 5888 3026 0 _007_
rlabel metal1 5566 2822 5566 2822 0 _008_
rlabel metal1 8510 4114 8510 4114 0 _009_
rlabel metal1 9476 2618 9476 2618 0 _010_
rlabel metal1 6118 6426 6118 6426 0 _011_
rlabel metal1 3450 5746 3450 5746 0 _012_
rlabel metal1 7314 7854 7314 7854 0 _013_
rlabel metal1 6624 8058 6624 8058 0 _014_
rlabel metal1 4830 4692 4830 4692 0 _015_
rlabel metal2 7590 8228 7590 8228 0 _016_
rlabel metal1 4370 5644 4370 5644 0 _017_
rlabel metal1 6302 7956 6302 7956 0 _018_
rlabel metal1 5474 6290 5474 6290 0 _019_
rlabel metal1 3772 4658 3772 4658 0 _020_
rlabel metal1 4462 5202 4462 5202 0 _021_
rlabel metal2 4922 8772 4922 8772 0 _022_
rlabel metal1 5060 5746 5060 5746 0 _023_
rlabel metal1 5382 8058 5382 8058 0 _024_
rlabel metal1 8050 8058 8050 8058 0 _025_
rlabel metal1 9890 4216 9890 4216 0 _026_
rlabel metal1 9154 4012 9154 4012 0 _027_
rlabel metal1 8096 3162 8096 3162 0 _028_
rlabel metal1 8832 3910 8832 3910 0 _029_
rlabel metal1 6072 3162 6072 3162 0 _030_
rlabel metal1 6348 4658 6348 4658 0 _031_
rlabel metal1 8648 2482 8648 2482 0 _032_
rlabel metal1 8740 2890 8740 2890 0 _033_
rlabel metal1 7866 4012 7866 4012 0 _034_
rlabel metal1 7958 4692 7958 4692 0 _035_
rlabel metal1 5980 2890 5980 2890 0 _036_
rlabel metal1 7268 4046 7268 4046 0 _037_
rlabel metal1 10074 6426 10074 6426 0 _038_
rlabel metal1 7406 5202 7406 5202 0 _039_
rlabel metal1 10166 5338 10166 5338 0 _040_
rlabel metal1 7084 4658 7084 4658 0 _041_
rlabel metal2 9982 1520 9982 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 8602 9622 8602 9622 0 ccff_head
rlabel metal1 9798 9146 9798 9146 0 ccff_tail
rlabel metal3 751 2516 751 2516 0 chanx_left_in[0]
rlabel metal3 820 3604 820 3604 0 chanx_left_in[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_in[2]
rlabel metal3 820 5780 820 5780 0 chanx_left_in[3]
rlabel metal3 1050 6868 1050 6868 0 chanx_left_in[4]
rlabel metal3 1050 7956 1050 7956 0 chanx_left_in[5]
rlabel metal3 820 9044 820 9044 0 chanx_left_in[6]
rlabel metal3 843 10132 843 10132 0 chanx_left_in[7]
rlabel metal3 843 11220 843 11220 0 chanx_left_in[8]
rlabel metal1 1150 9622 1150 9622 0 chanx_left_out[0]
rlabel metal1 1932 9622 1932 9622 0 chanx_left_out[1]
rlabel metal1 2944 9622 2944 9622 0 chanx_left_out[2]
rlabel metal1 3956 9622 3956 9622 0 chanx_left_out[3]
rlabel metal1 4968 9622 4968 9622 0 chanx_left_out[4]
rlabel metal1 6302 9622 6302 9622 0 chanx_left_out[5]
rlabel metal1 6992 9622 6992 9622 0 chanx_left_out[6]
rlabel metal1 8004 9622 8004 9622 0 chanx_left_out[7]
rlabel metal1 9246 9622 9246 9622 0 chanx_left_out[8]
rlabel metal3 9438 340 9438 340 0 chanx_right_in[0]
rlabel metal1 9246 2414 9246 2414 0 chanx_right_in[1]
rlabel metal1 5934 2482 5934 2482 0 chanx_right_in[2]
rlabel metal1 5106 3060 5106 3060 0 chanx_right_in[3]
rlabel metal1 10258 5168 10258 5168 0 chanx_right_in[4]
rlabel metal1 9430 3060 9430 3060 0 chanx_right_in[5]
rlabel metal1 10534 6800 10534 6800 0 chanx_right_in[6]
rlabel metal1 9476 8466 9476 8466 0 chanx_right_in[7]
rlabel metal1 9982 9588 9982 9588 0 chanx_right_in[8]
rlabel metal2 874 1554 874 1554 0 chanx_right_out[0]
rlabel metal2 1886 1520 1886 1520 0 chanx_right_out[1]
rlabel metal2 2898 1520 2898 1520 0 chanx_right_out[2]
rlabel metal2 3910 1520 3910 1520 0 chanx_right_out[3]
rlabel metal2 4922 959 4922 959 0 chanx_right_out[4]
rlabel metal2 5934 1078 5934 1078 0 chanx_right_out[5]
rlabel metal2 6946 1520 6946 1520 0 chanx_right_out[6]
rlabel metal2 7958 1520 7958 1520 0 chanx_right_out[7]
rlabel metal2 8970 1520 8970 1520 0 chanx_right_out[8]
rlabel metal1 6118 5270 6118 5270 0 clknet_0_prog_clk
rlabel metal2 6394 5168 6394 5168 0 clknet_1_0__leaf_prog_clk
rlabel metal1 8878 6290 8878 6290 0 clknet_1_1__leaf_prog_clk
rlabel metal2 7866 7514 7866 7514 0 mem_bottom_ipin_0.DFF_0_.Q
rlabel metal2 5934 7072 5934 7072 0 mem_bottom_ipin_0.DFF_1_.Q
rlabel metal1 7038 7276 7038 7276 0 mem_bottom_ipin_0.DFF_2_.Q
rlabel metal1 7820 6630 7820 6630 0 mem_bottom_ipin_1.DFF_0_.Q
rlabel metal1 9982 6222 9982 6222 0 mem_bottom_ipin_1.DFF_1_.Q
rlabel metal1 6394 3026 6394 3026 0 mem_top_ipin_0.DFF_0_.Q
rlabel metal1 9844 2414 9844 2414 0 mem_top_ipin_0.DFF_1_.Q
rlabel metal1 3450 3706 3450 3706 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 4600 4250 4600 4250 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 4324 5134 4324 5134 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 4278 5746 4278 5746 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 5152 9010 5152 9010 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal1 6716 7922 6716 7922 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal2 5014 5236 5014 5236 0 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4968 5610 4968 5610 0 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 5566 8636 5566 8636 0 mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 6072 5814 6072 5814 0 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6532 8330 6532 8330 0 mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 8280 8330 8280 8330 0 mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 6808 4114 6808 4114 0 mux_bottom_ipin_1.INVTX1_0_.out
rlabel metal2 6302 5066 6302 5066 0 mux_bottom_ipin_1.INVTX1_1_.out
rlabel metal1 7912 5134 7912 5134 0 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9706 7174 9706 7174 0 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5106 3162 5106 3162 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 6532 3162 6532 3162 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal1 7590 4658 7590 4658 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal1 8786 6222 8786 6222 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal1 7084 4250 7084 4250 0 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6900 3706 6900 3706 0 mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9568 4658 9568 4658 0 mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 8326 3808 8326 3808 0 mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 9798 4454 9798 4454 0 mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 6210 2448 6210 2448 0 mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 9144 7854 9144 7854 0 net1
rlabel metal1 1886 8840 1886 8840 0 net10
rlabel metal1 4922 4012 4922 4012 0 net11
rlabel metal1 8878 2550 8878 2550 0 net12
rlabel metal1 5658 2550 5658 2550 0 net13
rlabel metal1 4738 2822 4738 2822 0 net14
rlabel metal1 5980 5678 5980 5678 0 net15
rlabel metal1 9890 2890 9890 2890 0 net16
rlabel metal1 8602 6800 8602 6800 0 net17
rlabel metal1 9936 8466 9936 8466 0 net18
rlabel metal1 8970 8976 8970 8976 0 net19
rlabel metal1 2530 2992 2530 2992 0 net2
rlabel metal2 6394 2176 6394 2176 0 net20
rlabel metal1 10212 3706 10212 3706 0 net21
rlabel metal2 1886 5439 1886 5439 0 net22
rlabel metal1 2438 6426 2438 6426 0 net23
rlabel metal2 3358 9350 3358 9350 0 net24
rlabel metal2 4370 9350 4370 9350 0 net25
rlabel metal1 5520 5882 5520 5882 0 net26
rlabel metal1 10166 8568 10166 8568 0 net27
rlabel metal1 7452 9146 7452 9146 0 net28
rlabel metal1 9430 8602 9430 8602 0 net29
rlabel metal1 1610 4012 1610 4012 0 net3
rlabel metal2 9154 9350 9154 9350 0 net30
rlabel metal1 1840 2414 1840 2414 0 net31
rlabel metal1 2024 2414 2024 2414 0 net32
rlabel metal1 2990 2414 2990 2414 0 net33
rlabel metal1 3634 2414 3634 2414 0 net34
rlabel metal1 5290 2414 5290 2414 0 net35
rlabel metal2 6532 2414 6532 2414 0 net36
rlabel metal1 7038 2414 7038 2414 0 net37
rlabel metal1 7820 2346 7820 2346 0 net38
rlabel metal1 6095 1870 6095 1870 0 net39
rlabel metal1 2162 3502 2162 3502 0 net4
rlabel metal1 9338 9044 9338 9044 0 net40
rlabel metal1 10166 7514 10166 7514 0 net41
rlabel metal1 6486 8534 6486 8534 0 net42
rlabel metal1 8786 3638 8786 3638 0 net43
rlabel metal1 10028 6766 10028 6766 0 net44
rlabel metal1 8330 6358 8330 6358 0 net45
rlabel metal1 6568 6766 6568 6766 0 net46
rlabel viali 10170 5678 10170 5678 0 net47
rlabel metal1 7309 3502 7309 3502 0 net48
rlabel metal1 9200 3162 9200 3162 0 net49
rlabel metal1 1702 5202 1702 5202 0 net5
rlabel metal1 5515 6698 5515 6698 0 net50
rlabel metal1 5198 6970 5198 6970 0 net51
rlabel metal1 4048 6290 4048 6290 0 net6
rlabel metal2 3818 7854 3818 7854 0 net7
rlabel metal2 1610 8670 1610 8670 0 net8
rlabel metal2 2116 8806 2116 8806 0 net9
rlabel metal3 1970 1428 1970 1428 0 prog_clk
rlabel metal1 10166 9418 10166 9418 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal1 10304 8942 10304 8942 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
