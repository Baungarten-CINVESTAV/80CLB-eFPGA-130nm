magic
tech sky130A
magscale 1 2
timestamp 1710357890
<< obsli1 >>
rect 1104 2159 4876 13617
<< obsm1 >>
rect 1104 2128 5035 13648
<< obsm2 >>
rect 1398 2139 5029 13637
<< metal3 >>
rect 0 13608 800 13728
rect 5200 13064 6000 13184
rect 0 9800 800 9920
rect 5200 7896 6000 8016
rect 0 5992 800 6112
rect 5200 2728 6000 2848
<< obsm3 >>
rect 880 13528 5458 13633
rect 800 13264 5458 13528
rect 800 12984 5120 13264
rect 800 10000 5458 12984
rect 880 9720 5458 10000
rect 800 8096 5458 9720
rect 800 7816 5120 8096
rect 800 6192 5458 7816
rect 880 5912 5458 6192
rect 800 2928 5458 5912
rect 800 2648 5120 2928
rect 800 2143 5458 2648
<< metal4 >>
rect 1415 2128 1735 13648
rect 1886 2128 2206 13648
rect 2358 2128 2678 13648
rect 2829 2128 3149 13648
rect 3301 2128 3621 13648
rect 3772 2128 4092 13648
rect 4244 2128 4564 13648
rect 4715 2128 5035 13648
<< labels >>
rlabel metal3 s 5200 2728 6000 2848 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 5200 7896 6000 8016 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 5200 13064 6000 13184 6 gfpga_pad_GPIO_PAD
port 3 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 left_width_0_height_0_subtile_0__pin_inpad_0_
port 4 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 left_width_0_height_0_subtile_0__pin_outpad_0_
port 5 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 prog_clk
port 6 nsew signal input
rlabel metal4 s 1415 2128 1735 13648 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 2358 2128 2678 13648 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 3301 2128 3621 13648 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 4244 2128 4564 13648 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 1886 2128 2206 13648 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 2829 2128 3149 13648 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 3772 2128 4092 13648 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 4715 2128 5035 13648 6 vss
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 16000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 150518
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/grid_io_right/runs/24_03_13_13_24/results/signoff/grid_io_right.magic.gds
string GDS_START 40140
<< end >>

