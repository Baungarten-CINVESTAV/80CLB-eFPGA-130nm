magic
tech sky130A
magscale 1 2
timestamp 1710357643
<< obsli1 >>
rect 1104 2159 4876 9809
<< obsm1 >>
rect 1026 2128 5035 9840
<< metal2 >>
rect 1030 11200 1086 12000
rect 2962 11200 3018 12000
rect 4894 11200 4950 12000
<< obsm2 >>
rect 1142 11144 2906 11234
rect 3074 11144 4838 11234
rect 5006 11144 5029 11234
rect 1032 2139 5029 11144
<< metal3 >>
rect 0 8712 800 8832
rect 5200 8712 6000 8832
rect 5200 2728 6000 2848
<< obsm3 >>
rect 800 8912 5458 9825
rect 880 8632 5120 8912
rect 800 2928 5458 8632
rect 800 2648 5120 2928
rect 800 2143 5458 2648
<< metal4 >>
rect 1415 2128 1735 9840
rect 1886 2128 2206 9840
rect 2358 2128 2678 9840
rect 2829 2128 3149 9840
rect 3301 2128 3621 9840
rect 3772 2128 4092 9840
rect 4244 2128 4564 9840
rect 4715 2128 5035 9840
<< labels >>
rlabel metal3 s 5200 2728 6000 2848 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 5200 8712 6000 8832 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 4894 11200 4950 12000 6 gfpga_pad_GPIO_PAD
port 3 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 prog_clk
port 4 nsew signal input
rlabel metal2 s 1030 11200 1086 12000 6 top_width_0_height_0_subtile_0__pin_inpad_0_
port 5 nsew signal output
rlabel metal2 s 2962 11200 3018 12000 6 top_width_0_height_0_subtile_0__pin_outpad_0_
port 6 nsew signal input
rlabel metal4 s 1415 2128 1735 9840 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 2358 2128 2678 9840 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 3301 2128 3621 9840 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 4244 2128 4564 9840 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 1886 2128 2206 9840 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 2829 2128 3149 9840 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 3772 2128 4092 9840 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 4715 2128 5035 9840 6 vss
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 123200
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/grid_io_bottom/runs/24_03_13_13_20/results/signoff/grid_io_bottom.magic.gds
string GDS_START 44630
<< end >>

