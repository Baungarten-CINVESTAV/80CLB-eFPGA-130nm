VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__10_
  CLASS BLOCK ;
  FOREIGN sb_1__10_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 100.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 88.440 80.000 89.040 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 76.000 92.520 80.000 93.120 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 6.840 80.000 7.440 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 76.000 10.920 80.000 11.520 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 76.000 15.000 80.000 15.600 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 76.000 19.080 80.000 19.680 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 23.160 80.000 23.760 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 76.000 27.240 80.000 27.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 31.320 80.000 31.920 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 35.400 80.000 36.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 39.480 80.000 40.080 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 43.560 80.000 44.160 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 76.000 47.640 80.000 48.240 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 51.720 80.000 52.320 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 55.800 80.000 56.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 59.880 80.000 60.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 63.960 80.000 64.560 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 76.000 68.040 80.000 68.640 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 72.120 80.000 72.720 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 76.200 80.000 76.800 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END chany_bottom_out[8]
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 80.280 80.000 80.880 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.000 84.360 80.000 84.960 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.285 10.640 14.885 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.420 10.640 32.020 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.555 10.640 49.155 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.690 10.640 66.290 87.280 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.850 10.640 23.450 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.985 10.640 40.585 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.120 10.640 57.720 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.255 10.640 74.855 87.280 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 87.125 ;
      LAYER met1 ;
        RECT 1.910 6.160 75.370 87.280 ;
      LAYER met2 ;
        RECT 1.940 4.280 75.350 93.005 ;
        RECT 1.940 3.555 2.570 4.280 ;
        RECT 3.410 3.555 6.250 4.280 ;
        RECT 7.090 3.555 9.930 4.280 ;
        RECT 10.770 3.555 13.610 4.280 ;
        RECT 14.450 3.555 17.290 4.280 ;
        RECT 18.130 3.555 20.970 4.280 ;
        RECT 21.810 3.555 24.650 4.280 ;
        RECT 25.490 3.555 28.330 4.280 ;
        RECT 29.170 3.555 32.010 4.280 ;
        RECT 32.850 3.555 35.690 4.280 ;
        RECT 36.530 3.555 39.370 4.280 ;
        RECT 40.210 3.555 43.050 4.280 ;
        RECT 43.890 3.555 46.730 4.280 ;
        RECT 47.570 3.555 50.410 4.280 ;
        RECT 51.250 3.555 54.090 4.280 ;
        RECT 54.930 3.555 57.770 4.280 ;
        RECT 58.610 3.555 61.450 4.280 ;
        RECT 62.290 3.555 65.130 4.280 ;
        RECT 65.970 3.555 68.810 4.280 ;
        RECT 69.650 3.555 72.490 4.280 ;
        RECT 73.330 3.555 75.350 4.280 ;
      LAYER met3 ;
        RECT 4.400 92.120 75.600 92.985 ;
        RECT 2.825 89.440 76.050 92.120 ;
        RECT 4.400 88.040 75.600 89.440 ;
        RECT 2.825 85.360 76.050 88.040 ;
        RECT 4.400 83.960 75.600 85.360 ;
        RECT 2.825 81.280 76.050 83.960 ;
        RECT 4.400 79.880 75.600 81.280 ;
        RECT 2.825 77.200 76.050 79.880 ;
        RECT 4.400 75.800 75.600 77.200 ;
        RECT 2.825 73.120 76.050 75.800 ;
        RECT 4.400 71.720 75.600 73.120 ;
        RECT 2.825 69.040 76.050 71.720 ;
        RECT 4.400 67.640 75.600 69.040 ;
        RECT 2.825 64.960 76.050 67.640 ;
        RECT 4.400 63.560 75.600 64.960 ;
        RECT 2.825 60.880 76.050 63.560 ;
        RECT 4.400 59.480 75.600 60.880 ;
        RECT 2.825 56.800 76.050 59.480 ;
        RECT 4.400 55.400 75.600 56.800 ;
        RECT 2.825 52.720 76.050 55.400 ;
        RECT 4.400 51.320 75.600 52.720 ;
        RECT 2.825 48.640 76.050 51.320 ;
        RECT 4.400 47.240 75.600 48.640 ;
        RECT 2.825 44.560 76.050 47.240 ;
        RECT 4.400 43.160 75.600 44.560 ;
        RECT 2.825 40.480 76.050 43.160 ;
        RECT 4.400 39.080 75.600 40.480 ;
        RECT 2.825 36.400 76.050 39.080 ;
        RECT 4.400 35.000 75.600 36.400 ;
        RECT 2.825 32.320 76.050 35.000 ;
        RECT 4.400 30.920 75.600 32.320 ;
        RECT 2.825 28.240 76.050 30.920 ;
        RECT 4.400 26.840 75.600 28.240 ;
        RECT 2.825 24.160 76.050 26.840 ;
        RECT 4.400 22.760 75.600 24.160 ;
        RECT 2.825 20.080 76.050 22.760 ;
        RECT 4.400 18.680 75.600 20.080 ;
        RECT 2.825 16.000 76.050 18.680 ;
        RECT 4.400 14.600 75.600 16.000 ;
        RECT 2.825 11.920 76.050 14.600 ;
        RECT 4.400 10.520 75.600 11.920 ;
        RECT 2.825 7.840 76.050 10.520 ;
        RECT 2.825 6.440 75.600 7.840 ;
        RECT 2.825 3.575 76.050 6.440 ;
      LAYER met4 ;
        RECT 3.975 10.240 12.885 72.585 ;
        RECT 15.285 10.240 21.450 72.585 ;
        RECT 23.850 10.240 30.020 72.585 ;
        RECT 32.420 10.240 38.585 72.585 ;
        RECT 40.985 10.240 47.155 72.585 ;
        RECT 49.555 10.240 55.720 72.585 ;
        RECT 58.120 10.240 64.105 72.585 ;
        RECT 3.975 3.575 64.105 10.240 ;
  END
END sb_1__10_
END LIBRARY

