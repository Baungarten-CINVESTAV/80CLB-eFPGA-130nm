magic
tech sky130A
magscale 1 2
timestamp 1710358025
<< viali >>
rect 3157 8585 3191 8619
rect 3433 8449 3467 8483
rect 4537 8449 4571 8483
rect 4353 8313 4387 8347
rect 3341 7497 3375 7531
rect 3525 7361 3559 7395
rect 4537 7157 4571 7191
rect 4537 4573 4571 4607
rect 4353 4437 4387 4471
rect 4537 4233 4571 4267
rect 3157 4097 3191 4131
rect 3424 4097 3458 4131
rect 4353 2601 4387 2635
rect 4537 2397 4571 2431
<< metal1 >>
rect 1104 8730 5035 8752
rect 1104 8678 1892 8730
rect 1944 8678 1956 8730
rect 2008 8678 2020 8730
rect 2072 8678 2084 8730
rect 2136 8678 2148 8730
rect 2200 8678 2835 8730
rect 2887 8678 2899 8730
rect 2951 8678 2963 8730
rect 3015 8678 3027 8730
rect 3079 8678 3091 8730
rect 3143 8678 3778 8730
rect 3830 8678 3842 8730
rect 3894 8678 3906 8730
rect 3958 8678 3970 8730
rect 4022 8678 4034 8730
rect 4086 8678 4721 8730
rect 4773 8678 4785 8730
rect 4837 8678 4849 8730
rect 4901 8678 4913 8730
rect 4965 8678 4977 8730
rect 5029 8678 5035 8730
rect 1104 8656 5035 8678
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8616 3203 8619
rect 3234 8616 3240 8628
rect 3191 8588 3240 8616
rect 3191 8585 3203 8588
rect 3145 8579 3203 8585
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 5074 8508 5080 8560
rect 5132 8508 5138 8560
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3200 8452 3433 8480
rect 3200 8440 3206 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 5092 8480 5120 8508
rect 4571 8452 5120 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4341 8347 4399 8353
rect 4341 8344 4353 8347
rect 3752 8316 4353 8344
rect 3752 8304 3758 8316
rect 4341 8313 4353 8316
rect 4387 8313 4399 8347
rect 4341 8307 4399 8313
rect 1104 8186 4876 8208
rect 1104 8134 1421 8186
rect 1473 8134 1485 8186
rect 1537 8134 1549 8186
rect 1601 8134 1613 8186
rect 1665 8134 1677 8186
rect 1729 8134 2364 8186
rect 2416 8134 2428 8186
rect 2480 8134 2492 8186
rect 2544 8134 2556 8186
rect 2608 8134 2620 8186
rect 2672 8134 3307 8186
rect 3359 8134 3371 8186
rect 3423 8134 3435 8186
rect 3487 8134 3499 8186
rect 3551 8134 3563 8186
rect 3615 8134 4250 8186
rect 4302 8134 4314 8186
rect 4366 8134 4378 8186
rect 4430 8134 4442 8186
rect 4494 8134 4506 8186
rect 4558 8134 4876 8186
rect 1104 8112 4876 8134
rect 1104 7642 5035 7664
rect 1104 7590 1892 7642
rect 1944 7590 1956 7642
rect 2008 7590 2020 7642
rect 2072 7590 2084 7642
rect 2136 7590 2148 7642
rect 2200 7590 2835 7642
rect 2887 7590 2899 7642
rect 2951 7590 2963 7642
rect 3015 7590 3027 7642
rect 3079 7590 3091 7642
rect 3143 7590 3778 7642
rect 3830 7590 3842 7642
rect 3894 7590 3906 7642
rect 3958 7590 3970 7642
rect 4022 7590 4034 7642
rect 4086 7590 4721 7642
rect 4773 7590 4785 7642
rect 4837 7590 4849 7642
rect 4901 7590 4913 7642
rect 4965 7590 4977 7642
rect 5029 7590 5035 7642
rect 1104 7568 5035 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 3292 7500 3341 7528
rect 3292 7488 3298 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 3602 7488 3608 7540
rect 3660 7488 3666 7540
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3620 7392 3648 7488
rect 3559 7364 3648 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4890 7188 4896 7200
rect 4571 7160 4896 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 1104 7098 4876 7120
rect 1104 7046 1421 7098
rect 1473 7046 1485 7098
rect 1537 7046 1549 7098
rect 1601 7046 1613 7098
rect 1665 7046 1677 7098
rect 1729 7046 2364 7098
rect 2416 7046 2428 7098
rect 2480 7046 2492 7098
rect 2544 7046 2556 7098
rect 2608 7046 2620 7098
rect 2672 7046 3307 7098
rect 3359 7046 3371 7098
rect 3423 7046 3435 7098
rect 3487 7046 3499 7098
rect 3551 7046 3563 7098
rect 3615 7046 4250 7098
rect 4302 7046 4314 7098
rect 4366 7046 4378 7098
rect 4430 7046 4442 7098
rect 4494 7046 4506 7098
rect 4558 7046 4876 7098
rect 1104 7024 4876 7046
rect 1104 6554 5035 6576
rect 1104 6502 1892 6554
rect 1944 6502 1956 6554
rect 2008 6502 2020 6554
rect 2072 6502 2084 6554
rect 2136 6502 2148 6554
rect 2200 6502 2835 6554
rect 2887 6502 2899 6554
rect 2951 6502 2963 6554
rect 3015 6502 3027 6554
rect 3079 6502 3091 6554
rect 3143 6502 3778 6554
rect 3830 6502 3842 6554
rect 3894 6502 3906 6554
rect 3958 6502 3970 6554
rect 4022 6502 4034 6554
rect 4086 6502 4721 6554
rect 4773 6502 4785 6554
rect 4837 6502 4849 6554
rect 4901 6502 4913 6554
rect 4965 6502 4977 6554
rect 5029 6502 5035 6554
rect 1104 6480 5035 6502
rect 1104 6010 4876 6032
rect 1104 5958 1421 6010
rect 1473 5958 1485 6010
rect 1537 5958 1549 6010
rect 1601 5958 1613 6010
rect 1665 5958 1677 6010
rect 1729 5958 2364 6010
rect 2416 5958 2428 6010
rect 2480 5958 2492 6010
rect 2544 5958 2556 6010
rect 2608 5958 2620 6010
rect 2672 5958 3307 6010
rect 3359 5958 3371 6010
rect 3423 5958 3435 6010
rect 3487 5958 3499 6010
rect 3551 5958 3563 6010
rect 3615 5958 4250 6010
rect 4302 5958 4314 6010
rect 4366 5958 4378 6010
rect 4430 5958 4442 6010
rect 4494 5958 4506 6010
rect 4558 5958 4876 6010
rect 1104 5936 4876 5958
rect 1104 5466 5035 5488
rect 1104 5414 1892 5466
rect 1944 5414 1956 5466
rect 2008 5414 2020 5466
rect 2072 5414 2084 5466
rect 2136 5414 2148 5466
rect 2200 5414 2835 5466
rect 2887 5414 2899 5466
rect 2951 5414 2963 5466
rect 3015 5414 3027 5466
rect 3079 5414 3091 5466
rect 3143 5414 3778 5466
rect 3830 5414 3842 5466
rect 3894 5414 3906 5466
rect 3958 5414 3970 5466
rect 4022 5414 4034 5466
rect 4086 5414 4721 5466
rect 4773 5414 4785 5466
rect 4837 5414 4849 5466
rect 4901 5414 4913 5466
rect 4965 5414 4977 5466
rect 5029 5414 5035 5466
rect 1104 5392 5035 5414
rect 1104 4922 4876 4944
rect 1104 4870 1421 4922
rect 1473 4870 1485 4922
rect 1537 4870 1549 4922
rect 1601 4870 1613 4922
rect 1665 4870 1677 4922
rect 1729 4870 2364 4922
rect 2416 4870 2428 4922
rect 2480 4870 2492 4922
rect 2544 4870 2556 4922
rect 2608 4870 2620 4922
rect 2672 4870 3307 4922
rect 3359 4870 3371 4922
rect 3423 4870 3435 4922
rect 3487 4870 3499 4922
rect 3551 4870 3563 4922
rect 3615 4870 4250 4922
rect 4302 4870 4314 4922
rect 4366 4870 4378 4922
rect 4430 4870 4442 4922
rect 4494 4870 4506 4922
rect 4558 4870 4876 4922
rect 1104 4848 4876 4870
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 4338 4428 4344 4480
rect 4396 4428 4402 4480
rect 1104 4378 5035 4400
rect 1104 4326 1892 4378
rect 1944 4326 1956 4378
rect 2008 4326 2020 4378
rect 2072 4326 2084 4378
rect 2136 4326 2148 4378
rect 2200 4326 2835 4378
rect 2887 4326 2899 4378
rect 2951 4326 2963 4378
rect 3015 4326 3027 4378
rect 3079 4326 3091 4378
rect 3143 4326 3778 4378
rect 3830 4326 3842 4378
rect 3894 4326 3906 4378
rect 3958 4326 3970 4378
rect 4022 4326 4034 4378
rect 4086 4326 4721 4378
rect 4773 4326 4785 4378
rect 4837 4326 4849 4378
rect 4901 4326 4913 4378
rect 4965 4326 4977 4378
rect 5029 4326 5035 4378
rect 1104 4304 5035 4326
rect 4522 4224 4528 4276
rect 4580 4224 4586 4276
rect 3602 4196 3608 4208
rect 3344 4168 3608 4196
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3344 4128 3372 4168
rect 3602 4156 3608 4168
rect 3660 4156 3666 4208
rect 3191 4100 3372 4128
rect 3412 4131 3470 4137
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3412 4097 3424 4131
rect 3458 4128 3470 4131
rect 4154 4128 4160 4140
rect 3458 4100 4160 4128
rect 3458 4097 3470 4100
rect 3412 4091 3470 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 1104 3834 4876 3856
rect 1104 3782 1421 3834
rect 1473 3782 1485 3834
rect 1537 3782 1549 3834
rect 1601 3782 1613 3834
rect 1665 3782 1677 3834
rect 1729 3782 2364 3834
rect 2416 3782 2428 3834
rect 2480 3782 2492 3834
rect 2544 3782 2556 3834
rect 2608 3782 2620 3834
rect 2672 3782 3307 3834
rect 3359 3782 3371 3834
rect 3423 3782 3435 3834
rect 3487 3782 3499 3834
rect 3551 3782 3563 3834
rect 3615 3782 4250 3834
rect 4302 3782 4314 3834
rect 4366 3782 4378 3834
rect 4430 3782 4442 3834
rect 4494 3782 4506 3834
rect 4558 3782 4876 3834
rect 1104 3760 4876 3782
rect 1104 3290 5035 3312
rect 1104 3238 1892 3290
rect 1944 3238 1956 3290
rect 2008 3238 2020 3290
rect 2072 3238 2084 3290
rect 2136 3238 2148 3290
rect 2200 3238 2835 3290
rect 2887 3238 2899 3290
rect 2951 3238 2963 3290
rect 3015 3238 3027 3290
rect 3079 3238 3091 3290
rect 3143 3238 3778 3290
rect 3830 3238 3842 3290
rect 3894 3238 3906 3290
rect 3958 3238 3970 3290
rect 4022 3238 4034 3290
rect 4086 3238 4721 3290
rect 4773 3238 4785 3290
rect 4837 3238 4849 3290
rect 4901 3238 4913 3290
rect 4965 3238 4977 3290
rect 5029 3238 5035 3290
rect 1104 3216 5035 3238
rect 1104 2746 4876 2768
rect 1104 2694 1421 2746
rect 1473 2694 1485 2746
rect 1537 2694 1549 2746
rect 1601 2694 1613 2746
rect 1665 2694 1677 2746
rect 1729 2694 2364 2746
rect 2416 2694 2428 2746
rect 2480 2694 2492 2746
rect 2544 2694 2556 2746
rect 2608 2694 2620 2746
rect 2672 2694 3307 2746
rect 3359 2694 3371 2746
rect 3423 2694 3435 2746
rect 3487 2694 3499 2746
rect 3551 2694 3563 2746
rect 3615 2694 4250 2746
rect 4302 2694 4314 2746
rect 4366 2694 4378 2746
rect 4430 2694 4442 2746
rect 4494 2694 4506 2746
rect 4558 2694 4876 2746
rect 1104 2672 4876 2694
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4341 2635 4399 2641
rect 4341 2632 4353 2635
rect 4212 2604 4353 2632
rect 4212 2592 4218 2604
rect 4341 2601 4353 2604
rect 4387 2601 4399 2635
rect 4341 2595 4399 2601
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4571 2400 5120 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 5092 2372 5120 2400
rect 5074 2320 5080 2372
rect 5132 2320 5138 2372
rect 1104 2202 5035 2224
rect 1104 2150 1892 2202
rect 1944 2150 1956 2202
rect 2008 2150 2020 2202
rect 2072 2150 2084 2202
rect 2136 2150 2148 2202
rect 2200 2150 2835 2202
rect 2887 2150 2899 2202
rect 2951 2150 2963 2202
rect 3015 2150 3027 2202
rect 3079 2150 3091 2202
rect 3143 2150 3778 2202
rect 3830 2150 3842 2202
rect 3894 2150 3906 2202
rect 3958 2150 3970 2202
rect 4022 2150 4034 2202
rect 4086 2150 4721 2202
rect 4773 2150 4785 2202
rect 4837 2150 4849 2202
rect 4901 2150 4913 2202
rect 4965 2150 4977 2202
rect 5029 2150 5035 2202
rect 1104 2128 5035 2150
<< via1 >>
rect 1892 8678 1944 8730
rect 1956 8678 2008 8730
rect 2020 8678 2072 8730
rect 2084 8678 2136 8730
rect 2148 8678 2200 8730
rect 2835 8678 2887 8730
rect 2899 8678 2951 8730
rect 2963 8678 3015 8730
rect 3027 8678 3079 8730
rect 3091 8678 3143 8730
rect 3778 8678 3830 8730
rect 3842 8678 3894 8730
rect 3906 8678 3958 8730
rect 3970 8678 4022 8730
rect 4034 8678 4086 8730
rect 4721 8678 4773 8730
rect 4785 8678 4837 8730
rect 4849 8678 4901 8730
rect 4913 8678 4965 8730
rect 4977 8678 5029 8730
rect 3240 8576 3292 8628
rect 5080 8508 5132 8560
rect 3148 8440 3200 8492
rect 3700 8304 3752 8356
rect 1421 8134 1473 8186
rect 1485 8134 1537 8186
rect 1549 8134 1601 8186
rect 1613 8134 1665 8186
rect 1677 8134 1729 8186
rect 2364 8134 2416 8186
rect 2428 8134 2480 8186
rect 2492 8134 2544 8186
rect 2556 8134 2608 8186
rect 2620 8134 2672 8186
rect 3307 8134 3359 8186
rect 3371 8134 3423 8186
rect 3435 8134 3487 8186
rect 3499 8134 3551 8186
rect 3563 8134 3615 8186
rect 4250 8134 4302 8186
rect 4314 8134 4366 8186
rect 4378 8134 4430 8186
rect 4442 8134 4494 8186
rect 4506 8134 4558 8186
rect 1892 7590 1944 7642
rect 1956 7590 2008 7642
rect 2020 7590 2072 7642
rect 2084 7590 2136 7642
rect 2148 7590 2200 7642
rect 2835 7590 2887 7642
rect 2899 7590 2951 7642
rect 2963 7590 3015 7642
rect 3027 7590 3079 7642
rect 3091 7590 3143 7642
rect 3778 7590 3830 7642
rect 3842 7590 3894 7642
rect 3906 7590 3958 7642
rect 3970 7590 4022 7642
rect 4034 7590 4086 7642
rect 4721 7590 4773 7642
rect 4785 7590 4837 7642
rect 4849 7590 4901 7642
rect 4913 7590 4965 7642
rect 4977 7590 5029 7642
rect 3240 7488 3292 7540
rect 3608 7488 3660 7540
rect 4896 7148 4948 7200
rect 1421 7046 1473 7098
rect 1485 7046 1537 7098
rect 1549 7046 1601 7098
rect 1613 7046 1665 7098
rect 1677 7046 1729 7098
rect 2364 7046 2416 7098
rect 2428 7046 2480 7098
rect 2492 7046 2544 7098
rect 2556 7046 2608 7098
rect 2620 7046 2672 7098
rect 3307 7046 3359 7098
rect 3371 7046 3423 7098
rect 3435 7046 3487 7098
rect 3499 7046 3551 7098
rect 3563 7046 3615 7098
rect 4250 7046 4302 7098
rect 4314 7046 4366 7098
rect 4378 7046 4430 7098
rect 4442 7046 4494 7098
rect 4506 7046 4558 7098
rect 1892 6502 1944 6554
rect 1956 6502 2008 6554
rect 2020 6502 2072 6554
rect 2084 6502 2136 6554
rect 2148 6502 2200 6554
rect 2835 6502 2887 6554
rect 2899 6502 2951 6554
rect 2963 6502 3015 6554
rect 3027 6502 3079 6554
rect 3091 6502 3143 6554
rect 3778 6502 3830 6554
rect 3842 6502 3894 6554
rect 3906 6502 3958 6554
rect 3970 6502 4022 6554
rect 4034 6502 4086 6554
rect 4721 6502 4773 6554
rect 4785 6502 4837 6554
rect 4849 6502 4901 6554
rect 4913 6502 4965 6554
rect 4977 6502 5029 6554
rect 1421 5958 1473 6010
rect 1485 5958 1537 6010
rect 1549 5958 1601 6010
rect 1613 5958 1665 6010
rect 1677 5958 1729 6010
rect 2364 5958 2416 6010
rect 2428 5958 2480 6010
rect 2492 5958 2544 6010
rect 2556 5958 2608 6010
rect 2620 5958 2672 6010
rect 3307 5958 3359 6010
rect 3371 5958 3423 6010
rect 3435 5958 3487 6010
rect 3499 5958 3551 6010
rect 3563 5958 3615 6010
rect 4250 5958 4302 6010
rect 4314 5958 4366 6010
rect 4378 5958 4430 6010
rect 4442 5958 4494 6010
rect 4506 5958 4558 6010
rect 1892 5414 1944 5466
rect 1956 5414 2008 5466
rect 2020 5414 2072 5466
rect 2084 5414 2136 5466
rect 2148 5414 2200 5466
rect 2835 5414 2887 5466
rect 2899 5414 2951 5466
rect 2963 5414 3015 5466
rect 3027 5414 3079 5466
rect 3091 5414 3143 5466
rect 3778 5414 3830 5466
rect 3842 5414 3894 5466
rect 3906 5414 3958 5466
rect 3970 5414 4022 5466
rect 4034 5414 4086 5466
rect 4721 5414 4773 5466
rect 4785 5414 4837 5466
rect 4849 5414 4901 5466
rect 4913 5414 4965 5466
rect 4977 5414 5029 5466
rect 1421 4870 1473 4922
rect 1485 4870 1537 4922
rect 1549 4870 1601 4922
rect 1613 4870 1665 4922
rect 1677 4870 1729 4922
rect 2364 4870 2416 4922
rect 2428 4870 2480 4922
rect 2492 4870 2544 4922
rect 2556 4870 2608 4922
rect 2620 4870 2672 4922
rect 3307 4870 3359 4922
rect 3371 4870 3423 4922
rect 3435 4870 3487 4922
rect 3499 4870 3551 4922
rect 3563 4870 3615 4922
rect 4250 4870 4302 4922
rect 4314 4870 4366 4922
rect 4378 4870 4430 4922
rect 4442 4870 4494 4922
rect 4506 4870 4558 4922
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 1892 4326 1944 4378
rect 1956 4326 2008 4378
rect 2020 4326 2072 4378
rect 2084 4326 2136 4378
rect 2148 4326 2200 4378
rect 2835 4326 2887 4378
rect 2899 4326 2951 4378
rect 2963 4326 3015 4378
rect 3027 4326 3079 4378
rect 3091 4326 3143 4378
rect 3778 4326 3830 4378
rect 3842 4326 3894 4378
rect 3906 4326 3958 4378
rect 3970 4326 4022 4378
rect 4034 4326 4086 4378
rect 4721 4326 4773 4378
rect 4785 4326 4837 4378
rect 4849 4326 4901 4378
rect 4913 4326 4965 4378
rect 4977 4326 5029 4378
rect 4528 4267 4580 4276
rect 4528 4233 4537 4267
rect 4537 4233 4571 4267
rect 4571 4233 4580 4267
rect 4528 4224 4580 4233
rect 3608 4156 3660 4208
rect 4160 4088 4212 4140
rect 1421 3782 1473 3834
rect 1485 3782 1537 3834
rect 1549 3782 1601 3834
rect 1613 3782 1665 3834
rect 1677 3782 1729 3834
rect 2364 3782 2416 3834
rect 2428 3782 2480 3834
rect 2492 3782 2544 3834
rect 2556 3782 2608 3834
rect 2620 3782 2672 3834
rect 3307 3782 3359 3834
rect 3371 3782 3423 3834
rect 3435 3782 3487 3834
rect 3499 3782 3551 3834
rect 3563 3782 3615 3834
rect 4250 3782 4302 3834
rect 4314 3782 4366 3834
rect 4378 3782 4430 3834
rect 4442 3782 4494 3834
rect 4506 3782 4558 3834
rect 1892 3238 1944 3290
rect 1956 3238 2008 3290
rect 2020 3238 2072 3290
rect 2084 3238 2136 3290
rect 2148 3238 2200 3290
rect 2835 3238 2887 3290
rect 2899 3238 2951 3290
rect 2963 3238 3015 3290
rect 3027 3238 3079 3290
rect 3091 3238 3143 3290
rect 3778 3238 3830 3290
rect 3842 3238 3894 3290
rect 3906 3238 3958 3290
rect 3970 3238 4022 3290
rect 4034 3238 4086 3290
rect 4721 3238 4773 3290
rect 4785 3238 4837 3290
rect 4849 3238 4901 3290
rect 4913 3238 4965 3290
rect 4977 3238 5029 3290
rect 1421 2694 1473 2746
rect 1485 2694 1537 2746
rect 1549 2694 1601 2746
rect 1613 2694 1665 2746
rect 1677 2694 1729 2746
rect 2364 2694 2416 2746
rect 2428 2694 2480 2746
rect 2492 2694 2544 2746
rect 2556 2694 2608 2746
rect 2620 2694 2672 2746
rect 3307 2694 3359 2746
rect 3371 2694 3423 2746
rect 3435 2694 3487 2746
rect 3499 2694 3551 2746
rect 3563 2694 3615 2746
rect 4250 2694 4302 2746
rect 4314 2694 4366 2746
rect 4378 2694 4430 2746
rect 4442 2694 4494 2746
rect 4506 2694 4558 2746
rect 4160 2592 4212 2644
rect 5080 2320 5132 2372
rect 1892 2150 1944 2202
rect 1956 2150 2008 2202
rect 2020 2150 2072 2202
rect 2084 2150 2136 2202
rect 2148 2150 2200 2202
rect 2835 2150 2887 2202
rect 2899 2150 2951 2202
rect 2963 2150 3015 2202
rect 3027 2150 3079 2202
rect 3091 2150 3143 2202
rect 3778 2150 3830 2202
rect 3842 2150 3894 2202
rect 3906 2150 3958 2202
rect 3970 2150 4022 2202
rect 4034 2150 4086 2202
rect 4721 2150 4773 2202
rect 4785 2150 4837 2202
rect 4849 2150 4901 2202
rect 4913 2150 4965 2202
rect 4977 2150 5029 2202
<< metal2 >>
rect 2962 10200 3018 11000
rect 3068 10254 3280 10282
rect 2976 10146 3004 10200
rect 3068 10146 3096 10254
rect 2976 10118 3096 10146
rect 1892 8732 2200 8741
rect 1892 8730 1898 8732
rect 1954 8730 1978 8732
rect 2034 8730 2058 8732
rect 2114 8730 2138 8732
rect 2194 8730 2200 8732
rect 1954 8678 1956 8730
rect 2136 8678 2138 8730
rect 1892 8676 1898 8678
rect 1954 8676 1978 8678
rect 2034 8676 2058 8678
rect 2114 8676 2138 8678
rect 2194 8676 2200 8678
rect 1892 8667 2200 8676
rect 2835 8732 3143 8741
rect 2835 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3081 8732
rect 3137 8730 3143 8732
rect 2897 8678 2899 8730
rect 3079 8678 3081 8730
rect 2835 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3081 8678
rect 3137 8676 3143 8678
rect 2835 8667 3143 8676
rect 3252 8634 3280 10254
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 3778 8732 4086 8741
rect 3778 8730 3784 8732
rect 3840 8730 3864 8732
rect 3920 8730 3944 8732
rect 4000 8730 4024 8732
rect 4080 8730 4086 8732
rect 3840 8678 3842 8730
rect 4022 8678 4024 8730
rect 3778 8676 3784 8678
rect 3840 8676 3864 8678
rect 3920 8676 3944 8678
rect 4000 8676 4024 8678
rect 4080 8676 4086 8678
rect 3778 8667 4086 8676
rect 4721 8732 5029 8741
rect 4721 8730 4727 8732
rect 4783 8730 4807 8732
rect 4863 8730 4887 8732
rect 4943 8730 4967 8732
rect 5023 8730 5029 8732
rect 4783 8678 4785 8730
rect 4965 8678 4967 8730
rect 4721 8676 4727 8678
rect 4783 8676 4807 8678
rect 4863 8676 4887 8678
rect 4943 8676 4967 8678
rect 5023 8676 5029 8678
rect 4721 8667 5029 8676
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 5092 8566 5120 9551
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 1421 8188 1729 8197
rect 1421 8186 1427 8188
rect 1483 8186 1507 8188
rect 1563 8186 1587 8188
rect 1643 8186 1667 8188
rect 1723 8186 1729 8188
rect 1483 8134 1485 8186
rect 1665 8134 1667 8186
rect 1421 8132 1427 8134
rect 1483 8132 1507 8134
rect 1563 8132 1587 8134
rect 1643 8132 1667 8134
rect 1723 8132 1729 8134
rect 1421 8123 1729 8132
rect 2364 8188 2672 8197
rect 2364 8186 2370 8188
rect 2426 8186 2450 8188
rect 2506 8186 2530 8188
rect 2586 8186 2610 8188
rect 2666 8186 2672 8188
rect 2426 8134 2428 8186
rect 2608 8134 2610 8186
rect 2364 8132 2370 8134
rect 2426 8132 2450 8134
rect 2506 8132 2530 8134
rect 2586 8132 2610 8134
rect 2666 8132 2672 8134
rect 2364 8123 2672 8132
rect 3160 7834 3188 8434
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3307 8188 3615 8197
rect 3307 8186 3313 8188
rect 3369 8186 3393 8188
rect 3449 8186 3473 8188
rect 3529 8186 3553 8188
rect 3609 8186 3615 8188
rect 3369 8134 3371 8186
rect 3551 8134 3553 8186
rect 3307 8132 3313 8134
rect 3369 8132 3393 8134
rect 3449 8132 3473 8134
rect 3529 8132 3553 8134
rect 3609 8132 3615 8134
rect 3307 8123 3615 8132
rect 3712 7970 3740 8298
rect 4250 8188 4558 8197
rect 4250 8186 4256 8188
rect 4312 8186 4336 8188
rect 4392 8186 4416 8188
rect 4472 8186 4496 8188
rect 4552 8186 4558 8188
rect 4312 8134 4314 8186
rect 4494 8134 4496 8186
rect 4250 8132 4256 8134
rect 4312 8132 4336 8134
rect 4392 8132 4416 8134
rect 4472 8132 4496 8134
rect 4552 8132 4558 8134
rect 4250 8123 4558 8132
rect 3620 7942 3740 7970
rect 3160 7806 3280 7834
rect 1892 7644 2200 7653
rect 1892 7642 1898 7644
rect 1954 7642 1978 7644
rect 2034 7642 2058 7644
rect 2114 7642 2138 7644
rect 2194 7642 2200 7644
rect 1954 7590 1956 7642
rect 2136 7590 2138 7642
rect 1892 7588 1898 7590
rect 1954 7588 1978 7590
rect 2034 7588 2058 7590
rect 2114 7588 2138 7590
rect 2194 7588 2200 7590
rect 1892 7579 2200 7588
rect 2835 7644 3143 7653
rect 2835 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3081 7644
rect 3137 7642 3143 7644
rect 2897 7590 2899 7642
rect 3079 7590 3081 7642
rect 2835 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3081 7590
rect 3137 7588 3143 7590
rect 2835 7579 3143 7588
rect 3252 7546 3280 7806
rect 3620 7546 3648 7942
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 1421 7100 1729 7109
rect 1421 7098 1427 7100
rect 1483 7098 1507 7100
rect 1563 7098 1587 7100
rect 1643 7098 1667 7100
rect 1723 7098 1729 7100
rect 1483 7046 1485 7098
rect 1665 7046 1667 7098
rect 1421 7044 1427 7046
rect 1483 7044 1507 7046
rect 1563 7044 1587 7046
rect 1643 7044 1667 7046
rect 1723 7044 1729 7046
rect 1421 7035 1729 7044
rect 2364 7100 2672 7109
rect 2364 7098 2370 7100
rect 2426 7098 2450 7100
rect 2506 7098 2530 7100
rect 2586 7098 2610 7100
rect 2666 7098 2672 7100
rect 2426 7046 2428 7098
rect 2608 7046 2610 7098
rect 2364 7044 2370 7046
rect 2426 7044 2450 7046
rect 2506 7044 2530 7046
rect 2586 7044 2610 7046
rect 2666 7044 2672 7046
rect 2364 7035 2672 7044
rect 3307 7100 3615 7109
rect 3307 7098 3313 7100
rect 3369 7098 3393 7100
rect 3449 7098 3473 7100
rect 3529 7098 3553 7100
rect 3609 7098 3615 7100
rect 3369 7046 3371 7098
rect 3551 7046 3553 7098
rect 3307 7044 3313 7046
rect 3369 7044 3393 7046
rect 3449 7044 3473 7046
rect 3529 7044 3553 7046
rect 3609 7044 3615 7046
rect 3307 7035 3615 7044
rect 1892 6556 2200 6565
rect 1892 6554 1898 6556
rect 1954 6554 1978 6556
rect 2034 6554 2058 6556
rect 2114 6554 2138 6556
rect 2194 6554 2200 6556
rect 1954 6502 1956 6554
rect 2136 6502 2138 6554
rect 1892 6500 1898 6502
rect 1954 6500 1978 6502
rect 2034 6500 2058 6502
rect 2114 6500 2138 6502
rect 2194 6500 2200 6502
rect 1892 6491 2200 6500
rect 2835 6556 3143 6565
rect 2835 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3081 6556
rect 3137 6554 3143 6556
rect 2897 6502 2899 6554
rect 3079 6502 3081 6554
rect 2835 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3081 6502
rect 3137 6500 3143 6502
rect 2835 6491 3143 6500
rect 1421 6012 1729 6021
rect 1421 6010 1427 6012
rect 1483 6010 1507 6012
rect 1563 6010 1587 6012
rect 1643 6010 1667 6012
rect 1723 6010 1729 6012
rect 1483 5958 1485 6010
rect 1665 5958 1667 6010
rect 1421 5956 1427 5958
rect 1483 5956 1507 5958
rect 1563 5956 1587 5958
rect 1643 5956 1667 5958
rect 1723 5956 1729 5958
rect 1421 5947 1729 5956
rect 2364 6012 2672 6021
rect 2364 6010 2370 6012
rect 2426 6010 2450 6012
rect 2506 6010 2530 6012
rect 2586 6010 2610 6012
rect 2666 6010 2672 6012
rect 2426 5958 2428 6010
rect 2608 5958 2610 6010
rect 2364 5956 2370 5958
rect 2426 5956 2450 5958
rect 2506 5956 2530 5958
rect 2586 5956 2610 5958
rect 2666 5956 2672 5958
rect 2364 5947 2672 5956
rect 3307 6012 3615 6021
rect 3307 6010 3313 6012
rect 3369 6010 3393 6012
rect 3449 6010 3473 6012
rect 3529 6010 3553 6012
rect 3609 6010 3615 6012
rect 3369 5958 3371 6010
rect 3551 5958 3553 6010
rect 3307 5956 3313 5958
rect 3369 5956 3393 5958
rect 3449 5956 3473 5958
rect 3529 5956 3553 5958
rect 3609 5956 3615 5958
rect 3307 5947 3615 5956
rect 1892 5468 2200 5477
rect 1892 5466 1898 5468
rect 1954 5466 1978 5468
rect 2034 5466 2058 5468
rect 2114 5466 2138 5468
rect 2194 5466 2200 5468
rect 1954 5414 1956 5466
rect 2136 5414 2138 5466
rect 1892 5412 1898 5414
rect 1954 5412 1978 5414
rect 2034 5412 2058 5414
rect 2114 5412 2138 5414
rect 2194 5412 2200 5414
rect 1892 5403 2200 5412
rect 2835 5468 3143 5477
rect 2835 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3081 5468
rect 3137 5466 3143 5468
rect 2897 5414 2899 5466
rect 3079 5414 3081 5466
rect 2835 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3081 5414
rect 3137 5412 3143 5414
rect 2835 5403 3143 5412
rect 1421 4924 1729 4933
rect 1421 4922 1427 4924
rect 1483 4922 1507 4924
rect 1563 4922 1587 4924
rect 1643 4922 1667 4924
rect 1723 4922 1729 4924
rect 1483 4870 1485 4922
rect 1665 4870 1667 4922
rect 1421 4868 1427 4870
rect 1483 4868 1507 4870
rect 1563 4868 1587 4870
rect 1643 4868 1667 4870
rect 1723 4868 1729 4870
rect 1421 4859 1729 4868
rect 2364 4924 2672 4933
rect 2364 4922 2370 4924
rect 2426 4922 2450 4924
rect 2506 4922 2530 4924
rect 2586 4922 2610 4924
rect 2666 4922 2672 4924
rect 2426 4870 2428 4922
rect 2608 4870 2610 4922
rect 2364 4868 2370 4870
rect 2426 4868 2450 4870
rect 2506 4868 2530 4870
rect 2586 4868 2610 4870
rect 2666 4868 2672 4870
rect 2364 4859 2672 4868
rect 3307 4924 3615 4933
rect 3307 4922 3313 4924
rect 3369 4922 3393 4924
rect 3449 4922 3473 4924
rect 3529 4922 3553 4924
rect 3609 4922 3615 4924
rect 3369 4870 3371 4922
rect 3551 4870 3553 4922
rect 3307 4868 3313 4870
rect 3369 4868 3393 4870
rect 3449 4868 3473 4870
rect 3529 4868 3553 4870
rect 3609 4868 3615 4870
rect 3307 4859 3615 4868
rect 3712 4706 3740 7783
rect 3778 7644 4086 7653
rect 3778 7642 3784 7644
rect 3840 7642 3864 7644
rect 3920 7642 3944 7644
rect 4000 7642 4024 7644
rect 4080 7642 4086 7644
rect 3840 7590 3842 7642
rect 4022 7590 4024 7642
rect 3778 7588 3784 7590
rect 3840 7588 3864 7590
rect 3920 7588 3944 7590
rect 4000 7588 4024 7590
rect 4080 7588 4086 7590
rect 3778 7579 4086 7588
rect 4721 7644 5029 7653
rect 4721 7642 4727 7644
rect 4783 7642 4807 7644
rect 4863 7642 4887 7644
rect 4943 7642 4967 7644
rect 5023 7642 5029 7644
rect 4783 7590 4785 7642
rect 4965 7590 4967 7642
rect 4721 7588 4727 7590
rect 4783 7588 4807 7590
rect 4863 7588 4887 7590
rect 4943 7588 4967 7590
rect 5023 7588 5029 7590
rect 4721 7579 5029 7588
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4250 7100 4558 7109
rect 4250 7098 4256 7100
rect 4312 7098 4336 7100
rect 4392 7098 4416 7100
rect 4472 7098 4496 7100
rect 4552 7098 4558 7100
rect 4312 7046 4314 7098
rect 4494 7046 4496 7098
rect 4250 7044 4256 7046
rect 4312 7044 4336 7046
rect 4392 7044 4416 7046
rect 4472 7044 4496 7046
rect 4552 7044 4558 7046
rect 4250 7035 4558 7044
rect 4908 6905 4936 7142
rect 4894 6896 4950 6905
rect 4894 6831 4950 6840
rect 3778 6556 4086 6565
rect 3778 6554 3784 6556
rect 3840 6554 3864 6556
rect 3920 6554 3944 6556
rect 4000 6554 4024 6556
rect 4080 6554 4086 6556
rect 3840 6502 3842 6554
rect 4022 6502 4024 6554
rect 3778 6500 3784 6502
rect 3840 6500 3864 6502
rect 3920 6500 3944 6502
rect 4000 6500 4024 6502
rect 4080 6500 4086 6502
rect 3778 6491 4086 6500
rect 4721 6556 5029 6565
rect 4721 6554 4727 6556
rect 4783 6554 4807 6556
rect 4863 6554 4887 6556
rect 4943 6554 4967 6556
rect 5023 6554 5029 6556
rect 4783 6502 4785 6554
rect 4965 6502 4967 6554
rect 4721 6500 4727 6502
rect 4783 6500 4807 6502
rect 4863 6500 4887 6502
rect 4943 6500 4967 6502
rect 5023 6500 5029 6502
rect 4721 6491 5029 6500
rect 4250 6012 4558 6021
rect 4250 6010 4256 6012
rect 4312 6010 4336 6012
rect 4392 6010 4416 6012
rect 4472 6010 4496 6012
rect 4552 6010 4558 6012
rect 4312 5958 4314 6010
rect 4494 5958 4496 6010
rect 4250 5956 4256 5958
rect 4312 5956 4336 5958
rect 4392 5956 4416 5958
rect 4472 5956 4496 5958
rect 4552 5956 4558 5958
rect 4250 5947 4558 5956
rect 3778 5468 4086 5477
rect 3778 5466 3784 5468
rect 3840 5466 3864 5468
rect 3920 5466 3944 5468
rect 4000 5466 4024 5468
rect 4080 5466 4086 5468
rect 3840 5414 3842 5466
rect 4022 5414 4024 5466
rect 3778 5412 3784 5414
rect 3840 5412 3864 5414
rect 3920 5412 3944 5414
rect 4000 5412 4024 5414
rect 4080 5412 4086 5414
rect 3778 5403 4086 5412
rect 4721 5468 5029 5477
rect 4721 5466 4727 5468
rect 4783 5466 4807 5468
rect 4863 5466 4887 5468
rect 4943 5466 4967 5468
rect 5023 5466 5029 5468
rect 4783 5414 4785 5466
rect 4965 5414 4967 5466
rect 4721 5412 4727 5414
rect 4783 5412 4807 5414
rect 4863 5412 4887 5414
rect 4943 5412 4967 5414
rect 5023 5412 5029 5414
rect 4721 5403 5029 5412
rect 4250 4924 4558 4933
rect 4250 4922 4256 4924
rect 4312 4922 4336 4924
rect 4392 4922 4416 4924
rect 4472 4922 4496 4924
rect 4552 4922 4558 4924
rect 4312 4870 4314 4922
rect 4494 4870 4496 4922
rect 4250 4868 4256 4870
rect 4312 4868 4336 4870
rect 4392 4868 4416 4870
rect 4472 4868 4496 4870
rect 4552 4868 4558 4870
rect 4250 4859 4558 4868
rect 3620 4678 3740 4706
rect 1892 4380 2200 4389
rect 1892 4378 1898 4380
rect 1954 4378 1978 4380
rect 2034 4378 2058 4380
rect 2114 4378 2138 4380
rect 2194 4378 2200 4380
rect 1954 4326 1956 4378
rect 2136 4326 2138 4378
rect 1892 4324 1898 4326
rect 1954 4324 1978 4326
rect 2034 4324 2058 4326
rect 2114 4324 2138 4326
rect 2194 4324 2200 4326
rect 1892 4315 2200 4324
rect 2835 4380 3143 4389
rect 2835 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3081 4380
rect 3137 4378 3143 4380
rect 2897 4326 2899 4378
rect 3079 4326 3081 4378
rect 2835 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3081 4326
rect 3137 4324 3143 4326
rect 2835 4315 3143 4324
rect 3620 4214 3648 4678
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 3778 4380 4086 4389
rect 3778 4378 3784 4380
rect 3840 4378 3864 4380
rect 3920 4378 3944 4380
rect 4000 4378 4024 4380
rect 4080 4378 4086 4380
rect 3840 4326 3842 4378
rect 4022 4326 4024 4378
rect 3778 4324 3784 4326
rect 3840 4324 3864 4326
rect 3920 4324 3944 4326
rect 4000 4324 4024 4326
rect 4080 4324 4086 4326
rect 3778 4315 4086 4324
rect 3608 4208 3660 4214
rect 4356 4185 4384 4422
rect 4540 4282 4568 4558
rect 4721 4380 5029 4389
rect 4721 4378 4727 4380
rect 4783 4378 4807 4380
rect 4863 4378 4887 4380
rect 4943 4378 4967 4380
rect 5023 4378 5029 4380
rect 4783 4326 4785 4378
rect 4965 4326 4967 4378
rect 4721 4324 4727 4326
rect 4783 4324 4807 4326
rect 4863 4324 4887 4326
rect 4943 4324 4967 4326
rect 5023 4324 5029 4326
rect 4721 4315 5029 4324
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 3608 4150 3660 4156
rect 4342 4176 4398 4185
rect 4160 4140 4212 4146
rect 4342 4111 4398 4120
rect 4160 4082 4212 4088
rect 1421 3836 1729 3845
rect 1421 3834 1427 3836
rect 1483 3834 1507 3836
rect 1563 3834 1587 3836
rect 1643 3834 1667 3836
rect 1723 3834 1729 3836
rect 1483 3782 1485 3834
rect 1665 3782 1667 3834
rect 1421 3780 1427 3782
rect 1483 3780 1507 3782
rect 1563 3780 1587 3782
rect 1643 3780 1667 3782
rect 1723 3780 1729 3782
rect 1421 3771 1729 3780
rect 2364 3836 2672 3845
rect 2364 3834 2370 3836
rect 2426 3834 2450 3836
rect 2506 3834 2530 3836
rect 2586 3834 2610 3836
rect 2666 3834 2672 3836
rect 2426 3782 2428 3834
rect 2608 3782 2610 3834
rect 2364 3780 2370 3782
rect 2426 3780 2450 3782
rect 2506 3780 2530 3782
rect 2586 3780 2610 3782
rect 2666 3780 2672 3782
rect 2364 3771 2672 3780
rect 3307 3836 3615 3845
rect 3307 3834 3313 3836
rect 3369 3834 3393 3836
rect 3449 3834 3473 3836
rect 3529 3834 3553 3836
rect 3609 3834 3615 3836
rect 3369 3782 3371 3834
rect 3551 3782 3553 3834
rect 3307 3780 3313 3782
rect 3369 3780 3393 3782
rect 3449 3780 3473 3782
rect 3529 3780 3553 3782
rect 3609 3780 3615 3782
rect 3307 3771 3615 3780
rect 1892 3292 2200 3301
rect 1892 3290 1898 3292
rect 1954 3290 1978 3292
rect 2034 3290 2058 3292
rect 2114 3290 2138 3292
rect 2194 3290 2200 3292
rect 1954 3238 1956 3290
rect 2136 3238 2138 3290
rect 1892 3236 1898 3238
rect 1954 3236 1978 3238
rect 2034 3236 2058 3238
rect 2114 3236 2138 3238
rect 2194 3236 2200 3238
rect 1892 3227 2200 3236
rect 2835 3292 3143 3301
rect 2835 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3081 3292
rect 3137 3290 3143 3292
rect 2897 3238 2899 3290
rect 3079 3238 3081 3290
rect 2835 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3081 3238
rect 3137 3236 3143 3238
rect 2835 3227 3143 3236
rect 3778 3292 4086 3301
rect 3778 3290 3784 3292
rect 3840 3290 3864 3292
rect 3920 3290 3944 3292
rect 4000 3290 4024 3292
rect 4080 3290 4086 3292
rect 3840 3238 3842 3290
rect 4022 3238 4024 3290
rect 3778 3236 3784 3238
rect 3840 3236 3864 3238
rect 3920 3236 3944 3238
rect 4000 3236 4024 3238
rect 4080 3236 4086 3238
rect 3778 3227 4086 3236
rect 1421 2748 1729 2757
rect 1421 2746 1427 2748
rect 1483 2746 1507 2748
rect 1563 2746 1587 2748
rect 1643 2746 1667 2748
rect 1723 2746 1729 2748
rect 1483 2694 1485 2746
rect 1665 2694 1667 2746
rect 1421 2692 1427 2694
rect 1483 2692 1507 2694
rect 1563 2692 1587 2694
rect 1643 2692 1667 2694
rect 1723 2692 1729 2694
rect 1421 2683 1729 2692
rect 2364 2748 2672 2757
rect 2364 2746 2370 2748
rect 2426 2746 2450 2748
rect 2506 2746 2530 2748
rect 2586 2746 2610 2748
rect 2666 2746 2672 2748
rect 2426 2694 2428 2746
rect 2608 2694 2610 2746
rect 2364 2692 2370 2694
rect 2426 2692 2450 2694
rect 2506 2692 2530 2694
rect 2586 2692 2610 2694
rect 2666 2692 2672 2694
rect 2364 2683 2672 2692
rect 3307 2748 3615 2757
rect 3307 2746 3313 2748
rect 3369 2746 3393 2748
rect 3449 2746 3473 2748
rect 3529 2746 3553 2748
rect 3609 2746 3615 2748
rect 3369 2694 3371 2746
rect 3551 2694 3553 2746
rect 3307 2692 3313 2694
rect 3369 2692 3393 2694
rect 3449 2692 3473 2694
rect 3529 2692 3553 2694
rect 3609 2692 3615 2694
rect 3307 2683 3615 2692
rect 4172 2650 4200 4082
rect 4250 3836 4558 3845
rect 4250 3834 4256 3836
rect 4312 3834 4336 3836
rect 4392 3834 4416 3836
rect 4472 3834 4496 3836
rect 4552 3834 4558 3836
rect 4312 3782 4314 3834
rect 4494 3782 4496 3834
rect 4250 3780 4256 3782
rect 4312 3780 4336 3782
rect 4392 3780 4416 3782
rect 4472 3780 4496 3782
rect 4552 3780 4558 3782
rect 4250 3771 4558 3780
rect 4721 3292 5029 3301
rect 4721 3290 4727 3292
rect 4783 3290 4807 3292
rect 4863 3290 4887 3292
rect 4943 3290 4967 3292
rect 5023 3290 5029 3292
rect 4783 3238 4785 3290
rect 4965 3238 4967 3290
rect 4721 3236 4727 3238
rect 4783 3236 4807 3238
rect 4863 3236 4887 3238
rect 4943 3236 4967 3238
rect 5023 3236 5029 3238
rect 4721 3227 5029 3236
rect 4250 2748 4558 2757
rect 4250 2746 4256 2748
rect 4312 2746 4336 2748
rect 4392 2746 4416 2748
rect 4472 2746 4496 2748
rect 4552 2746 4558 2748
rect 4312 2694 4314 2746
rect 4494 2694 4496 2746
rect 4250 2692 4256 2694
rect 4312 2692 4336 2694
rect 4392 2692 4416 2694
rect 4472 2692 4496 2694
rect 4552 2692 4558 2694
rect 4250 2683 4558 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 1892 2204 2200 2213
rect 1892 2202 1898 2204
rect 1954 2202 1978 2204
rect 2034 2202 2058 2204
rect 2114 2202 2138 2204
rect 2194 2202 2200 2204
rect 1954 2150 1956 2202
rect 2136 2150 2138 2202
rect 1892 2148 1898 2150
rect 1954 2148 1978 2150
rect 2034 2148 2058 2150
rect 2114 2148 2138 2150
rect 2194 2148 2200 2150
rect 1892 2139 2200 2148
rect 2835 2204 3143 2213
rect 2835 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3081 2204
rect 3137 2202 3143 2204
rect 2897 2150 2899 2202
rect 3079 2150 3081 2202
rect 2835 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3081 2150
rect 3137 2148 3143 2150
rect 2835 2139 3143 2148
rect 3778 2204 4086 2213
rect 3778 2202 3784 2204
rect 3840 2202 3864 2204
rect 3920 2202 3944 2204
rect 4000 2202 4024 2204
rect 4080 2202 4086 2204
rect 3840 2150 3842 2202
rect 4022 2150 4024 2202
rect 3778 2148 3784 2150
rect 3840 2148 3864 2150
rect 3920 2148 3944 2150
rect 4000 2148 4024 2150
rect 4080 2148 4086 2150
rect 3778 2139 4086 2148
rect 4721 2204 5029 2213
rect 4721 2202 4727 2204
rect 4783 2202 4807 2204
rect 4863 2202 4887 2204
rect 4943 2202 4967 2204
rect 5023 2202 5029 2204
rect 4783 2150 4785 2202
rect 4965 2150 4967 2202
rect 4721 2148 4727 2150
rect 4783 2148 4807 2150
rect 4863 2148 4887 2150
rect 4943 2148 4967 2150
rect 5023 2148 5029 2150
rect 4721 2139 5029 2148
rect 5092 1465 5120 2314
rect 5078 1456 5134 1465
rect 5078 1391 5134 1400
<< via2 >>
rect 1898 8730 1954 8732
rect 1978 8730 2034 8732
rect 2058 8730 2114 8732
rect 2138 8730 2194 8732
rect 1898 8678 1944 8730
rect 1944 8678 1954 8730
rect 1978 8678 2008 8730
rect 2008 8678 2020 8730
rect 2020 8678 2034 8730
rect 2058 8678 2072 8730
rect 2072 8678 2084 8730
rect 2084 8678 2114 8730
rect 2138 8678 2148 8730
rect 2148 8678 2194 8730
rect 1898 8676 1954 8678
rect 1978 8676 2034 8678
rect 2058 8676 2114 8678
rect 2138 8676 2194 8678
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 3081 8730 3137 8732
rect 2841 8678 2887 8730
rect 2887 8678 2897 8730
rect 2921 8678 2951 8730
rect 2951 8678 2963 8730
rect 2963 8678 2977 8730
rect 3001 8678 3015 8730
rect 3015 8678 3027 8730
rect 3027 8678 3057 8730
rect 3081 8678 3091 8730
rect 3091 8678 3137 8730
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 3081 8676 3137 8678
rect 5078 9560 5134 9616
rect 3784 8730 3840 8732
rect 3864 8730 3920 8732
rect 3944 8730 4000 8732
rect 4024 8730 4080 8732
rect 3784 8678 3830 8730
rect 3830 8678 3840 8730
rect 3864 8678 3894 8730
rect 3894 8678 3906 8730
rect 3906 8678 3920 8730
rect 3944 8678 3958 8730
rect 3958 8678 3970 8730
rect 3970 8678 4000 8730
rect 4024 8678 4034 8730
rect 4034 8678 4080 8730
rect 3784 8676 3840 8678
rect 3864 8676 3920 8678
rect 3944 8676 4000 8678
rect 4024 8676 4080 8678
rect 4727 8730 4783 8732
rect 4807 8730 4863 8732
rect 4887 8730 4943 8732
rect 4967 8730 5023 8732
rect 4727 8678 4773 8730
rect 4773 8678 4783 8730
rect 4807 8678 4837 8730
rect 4837 8678 4849 8730
rect 4849 8678 4863 8730
rect 4887 8678 4901 8730
rect 4901 8678 4913 8730
rect 4913 8678 4943 8730
rect 4967 8678 4977 8730
rect 4977 8678 5023 8730
rect 4727 8676 4783 8678
rect 4807 8676 4863 8678
rect 4887 8676 4943 8678
rect 4967 8676 5023 8678
rect 1427 8186 1483 8188
rect 1507 8186 1563 8188
rect 1587 8186 1643 8188
rect 1667 8186 1723 8188
rect 1427 8134 1473 8186
rect 1473 8134 1483 8186
rect 1507 8134 1537 8186
rect 1537 8134 1549 8186
rect 1549 8134 1563 8186
rect 1587 8134 1601 8186
rect 1601 8134 1613 8186
rect 1613 8134 1643 8186
rect 1667 8134 1677 8186
rect 1677 8134 1723 8186
rect 1427 8132 1483 8134
rect 1507 8132 1563 8134
rect 1587 8132 1643 8134
rect 1667 8132 1723 8134
rect 2370 8186 2426 8188
rect 2450 8186 2506 8188
rect 2530 8186 2586 8188
rect 2610 8186 2666 8188
rect 2370 8134 2416 8186
rect 2416 8134 2426 8186
rect 2450 8134 2480 8186
rect 2480 8134 2492 8186
rect 2492 8134 2506 8186
rect 2530 8134 2544 8186
rect 2544 8134 2556 8186
rect 2556 8134 2586 8186
rect 2610 8134 2620 8186
rect 2620 8134 2666 8186
rect 2370 8132 2426 8134
rect 2450 8132 2506 8134
rect 2530 8132 2586 8134
rect 2610 8132 2666 8134
rect 3313 8186 3369 8188
rect 3393 8186 3449 8188
rect 3473 8186 3529 8188
rect 3553 8186 3609 8188
rect 3313 8134 3359 8186
rect 3359 8134 3369 8186
rect 3393 8134 3423 8186
rect 3423 8134 3435 8186
rect 3435 8134 3449 8186
rect 3473 8134 3487 8186
rect 3487 8134 3499 8186
rect 3499 8134 3529 8186
rect 3553 8134 3563 8186
rect 3563 8134 3609 8186
rect 3313 8132 3369 8134
rect 3393 8132 3449 8134
rect 3473 8132 3529 8134
rect 3553 8132 3609 8134
rect 4256 8186 4312 8188
rect 4336 8186 4392 8188
rect 4416 8186 4472 8188
rect 4496 8186 4552 8188
rect 4256 8134 4302 8186
rect 4302 8134 4312 8186
rect 4336 8134 4366 8186
rect 4366 8134 4378 8186
rect 4378 8134 4392 8186
rect 4416 8134 4430 8186
rect 4430 8134 4442 8186
rect 4442 8134 4472 8186
rect 4496 8134 4506 8186
rect 4506 8134 4552 8186
rect 4256 8132 4312 8134
rect 4336 8132 4392 8134
rect 4416 8132 4472 8134
rect 4496 8132 4552 8134
rect 1898 7642 1954 7644
rect 1978 7642 2034 7644
rect 2058 7642 2114 7644
rect 2138 7642 2194 7644
rect 1898 7590 1944 7642
rect 1944 7590 1954 7642
rect 1978 7590 2008 7642
rect 2008 7590 2020 7642
rect 2020 7590 2034 7642
rect 2058 7590 2072 7642
rect 2072 7590 2084 7642
rect 2084 7590 2114 7642
rect 2138 7590 2148 7642
rect 2148 7590 2194 7642
rect 1898 7588 1954 7590
rect 1978 7588 2034 7590
rect 2058 7588 2114 7590
rect 2138 7588 2194 7590
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 3081 7642 3137 7644
rect 2841 7590 2887 7642
rect 2887 7590 2897 7642
rect 2921 7590 2951 7642
rect 2951 7590 2963 7642
rect 2963 7590 2977 7642
rect 3001 7590 3015 7642
rect 3015 7590 3027 7642
rect 3027 7590 3057 7642
rect 3081 7590 3091 7642
rect 3091 7590 3137 7642
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 3081 7588 3137 7590
rect 3698 7792 3754 7848
rect 1427 7098 1483 7100
rect 1507 7098 1563 7100
rect 1587 7098 1643 7100
rect 1667 7098 1723 7100
rect 1427 7046 1473 7098
rect 1473 7046 1483 7098
rect 1507 7046 1537 7098
rect 1537 7046 1549 7098
rect 1549 7046 1563 7098
rect 1587 7046 1601 7098
rect 1601 7046 1613 7098
rect 1613 7046 1643 7098
rect 1667 7046 1677 7098
rect 1677 7046 1723 7098
rect 1427 7044 1483 7046
rect 1507 7044 1563 7046
rect 1587 7044 1643 7046
rect 1667 7044 1723 7046
rect 2370 7098 2426 7100
rect 2450 7098 2506 7100
rect 2530 7098 2586 7100
rect 2610 7098 2666 7100
rect 2370 7046 2416 7098
rect 2416 7046 2426 7098
rect 2450 7046 2480 7098
rect 2480 7046 2492 7098
rect 2492 7046 2506 7098
rect 2530 7046 2544 7098
rect 2544 7046 2556 7098
rect 2556 7046 2586 7098
rect 2610 7046 2620 7098
rect 2620 7046 2666 7098
rect 2370 7044 2426 7046
rect 2450 7044 2506 7046
rect 2530 7044 2586 7046
rect 2610 7044 2666 7046
rect 3313 7098 3369 7100
rect 3393 7098 3449 7100
rect 3473 7098 3529 7100
rect 3553 7098 3609 7100
rect 3313 7046 3359 7098
rect 3359 7046 3369 7098
rect 3393 7046 3423 7098
rect 3423 7046 3435 7098
rect 3435 7046 3449 7098
rect 3473 7046 3487 7098
rect 3487 7046 3499 7098
rect 3499 7046 3529 7098
rect 3553 7046 3563 7098
rect 3563 7046 3609 7098
rect 3313 7044 3369 7046
rect 3393 7044 3449 7046
rect 3473 7044 3529 7046
rect 3553 7044 3609 7046
rect 1898 6554 1954 6556
rect 1978 6554 2034 6556
rect 2058 6554 2114 6556
rect 2138 6554 2194 6556
rect 1898 6502 1944 6554
rect 1944 6502 1954 6554
rect 1978 6502 2008 6554
rect 2008 6502 2020 6554
rect 2020 6502 2034 6554
rect 2058 6502 2072 6554
rect 2072 6502 2084 6554
rect 2084 6502 2114 6554
rect 2138 6502 2148 6554
rect 2148 6502 2194 6554
rect 1898 6500 1954 6502
rect 1978 6500 2034 6502
rect 2058 6500 2114 6502
rect 2138 6500 2194 6502
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 3081 6554 3137 6556
rect 2841 6502 2887 6554
rect 2887 6502 2897 6554
rect 2921 6502 2951 6554
rect 2951 6502 2963 6554
rect 2963 6502 2977 6554
rect 3001 6502 3015 6554
rect 3015 6502 3027 6554
rect 3027 6502 3057 6554
rect 3081 6502 3091 6554
rect 3091 6502 3137 6554
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 3081 6500 3137 6502
rect 1427 6010 1483 6012
rect 1507 6010 1563 6012
rect 1587 6010 1643 6012
rect 1667 6010 1723 6012
rect 1427 5958 1473 6010
rect 1473 5958 1483 6010
rect 1507 5958 1537 6010
rect 1537 5958 1549 6010
rect 1549 5958 1563 6010
rect 1587 5958 1601 6010
rect 1601 5958 1613 6010
rect 1613 5958 1643 6010
rect 1667 5958 1677 6010
rect 1677 5958 1723 6010
rect 1427 5956 1483 5958
rect 1507 5956 1563 5958
rect 1587 5956 1643 5958
rect 1667 5956 1723 5958
rect 2370 6010 2426 6012
rect 2450 6010 2506 6012
rect 2530 6010 2586 6012
rect 2610 6010 2666 6012
rect 2370 5958 2416 6010
rect 2416 5958 2426 6010
rect 2450 5958 2480 6010
rect 2480 5958 2492 6010
rect 2492 5958 2506 6010
rect 2530 5958 2544 6010
rect 2544 5958 2556 6010
rect 2556 5958 2586 6010
rect 2610 5958 2620 6010
rect 2620 5958 2666 6010
rect 2370 5956 2426 5958
rect 2450 5956 2506 5958
rect 2530 5956 2586 5958
rect 2610 5956 2666 5958
rect 3313 6010 3369 6012
rect 3393 6010 3449 6012
rect 3473 6010 3529 6012
rect 3553 6010 3609 6012
rect 3313 5958 3359 6010
rect 3359 5958 3369 6010
rect 3393 5958 3423 6010
rect 3423 5958 3435 6010
rect 3435 5958 3449 6010
rect 3473 5958 3487 6010
rect 3487 5958 3499 6010
rect 3499 5958 3529 6010
rect 3553 5958 3563 6010
rect 3563 5958 3609 6010
rect 3313 5956 3369 5958
rect 3393 5956 3449 5958
rect 3473 5956 3529 5958
rect 3553 5956 3609 5958
rect 1898 5466 1954 5468
rect 1978 5466 2034 5468
rect 2058 5466 2114 5468
rect 2138 5466 2194 5468
rect 1898 5414 1944 5466
rect 1944 5414 1954 5466
rect 1978 5414 2008 5466
rect 2008 5414 2020 5466
rect 2020 5414 2034 5466
rect 2058 5414 2072 5466
rect 2072 5414 2084 5466
rect 2084 5414 2114 5466
rect 2138 5414 2148 5466
rect 2148 5414 2194 5466
rect 1898 5412 1954 5414
rect 1978 5412 2034 5414
rect 2058 5412 2114 5414
rect 2138 5412 2194 5414
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 3081 5466 3137 5468
rect 2841 5414 2887 5466
rect 2887 5414 2897 5466
rect 2921 5414 2951 5466
rect 2951 5414 2963 5466
rect 2963 5414 2977 5466
rect 3001 5414 3015 5466
rect 3015 5414 3027 5466
rect 3027 5414 3057 5466
rect 3081 5414 3091 5466
rect 3091 5414 3137 5466
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 3081 5412 3137 5414
rect 1427 4922 1483 4924
rect 1507 4922 1563 4924
rect 1587 4922 1643 4924
rect 1667 4922 1723 4924
rect 1427 4870 1473 4922
rect 1473 4870 1483 4922
rect 1507 4870 1537 4922
rect 1537 4870 1549 4922
rect 1549 4870 1563 4922
rect 1587 4870 1601 4922
rect 1601 4870 1613 4922
rect 1613 4870 1643 4922
rect 1667 4870 1677 4922
rect 1677 4870 1723 4922
rect 1427 4868 1483 4870
rect 1507 4868 1563 4870
rect 1587 4868 1643 4870
rect 1667 4868 1723 4870
rect 2370 4922 2426 4924
rect 2450 4922 2506 4924
rect 2530 4922 2586 4924
rect 2610 4922 2666 4924
rect 2370 4870 2416 4922
rect 2416 4870 2426 4922
rect 2450 4870 2480 4922
rect 2480 4870 2492 4922
rect 2492 4870 2506 4922
rect 2530 4870 2544 4922
rect 2544 4870 2556 4922
rect 2556 4870 2586 4922
rect 2610 4870 2620 4922
rect 2620 4870 2666 4922
rect 2370 4868 2426 4870
rect 2450 4868 2506 4870
rect 2530 4868 2586 4870
rect 2610 4868 2666 4870
rect 3313 4922 3369 4924
rect 3393 4922 3449 4924
rect 3473 4922 3529 4924
rect 3553 4922 3609 4924
rect 3313 4870 3359 4922
rect 3359 4870 3369 4922
rect 3393 4870 3423 4922
rect 3423 4870 3435 4922
rect 3435 4870 3449 4922
rect 3473 4870 3487 4922
rect 3487 4870 3499 4922
rect 3499 4870 3529 4922
rect 3553 4870 3563 4922
rect 3563 4870 3609 4922
rect 3313 4868 3369 4870
rect 3393 4868 3449 4870
rect 3473 4868 3529 4870
rect 3553 4868 3609 4870
rect 3784 7642 3840 7644
rect 3864 7642 3920 7644
rect 3944 7642 4000 7644
rect 4024 7642 4080 7644
rect 3784 7590 3830 7642
rect 3830 7590 3840 7642
rect 3864 7590 3894 7642
rect 3894 7590 3906 7642
rect 3906 7590 3920 7642
rect 3944 7590 3958 7642
rect 3958 7590 3970 7642
rect 3970 7590 4000 7642
rect 4024 7590 4034 7642
rect 4034 7590 4080 7642
rect 3784 7588 3840 7590
rect 3864 7588 3920 7590
rect 3944 7588 4000 7590
rect 4024 7588 4080 7590
rect 4727 7642 4783 7644
rect 4807 7642 4863 7644
rect 4887 7642 4943 7644
rect 4967 7642 5023 7644
rect 4727 7590 4773 7642
rect 4773 7590 4783 7642
rect 4807 7590 4837 7642
rect 4837 7590 4849 7642
rect 4849 7590 4863 7642
rect 4887 7590 4901 7642
rect 4901 7590 4913 7642
rect 4913 7590 4943 7642
rect 4967 7590 4977 7642
rect 4977 7590 5023 7642
rect 4727 7588 4783 7590
rect 4807 7588 4863 7590
rect 4887 7588 4943 7590
rect 4967 7588 5023 7590
rect 4256 7098 4312 7100
rect 4336 7098 4392 7100
rect 4416 7098 4472 7100
rect 4496 7098 4552 7100
rect 4256 7046 4302 7098
rect 4302 7046 4312 7098
rect 4336 7046 4366 7098
rect 4366 7046 4378 7098
rect 4378 7046 4392 7098
rect 4416 7046 4430 7098
rect 4430 7046 4442 7098
rect 4442 7046 4472 7098
rect 4496 7046 4506 7098
rect 4506 7046 4552 7098
rect 4256 7044 4312 7046
rect 4336 7044 4392 7046
rect 4416 7044 4472 7046
rect 4496 7044 4552 7046
rect 4894 6840 4950 6896
rect 3784 6554 3840 6556
rect 3864 6554 3920 6556
rect 3944 6554 4000 6556
rect 4024 6554 4080 6556
rect 3784 6502 3830 6554
rect 3830 6502 3840 6554
rect 3864 6502 3894 6554
rect 3894 6502 3906 6554
rect 3906 6502 3920 6554
rect 3944 6502 3958 6554
rect 3958 6502 3970 6554
rect 3970 6502 4000 6554
rect 4024 6502 4034 6554
rect 4034 6502 4080 6554
rect 3784 6500 3840 6502
rect 3864 6500 3920 6502
rect 3944 6500 4000 6502
rect 4024 6500 4080 6502
rect 4727 6554 4783 6556
rect 4807 6554 4863 6556
rect 4887 6554 4943 6556
rect 4967 6554 5023 6556
rect 4727 6502 4773 6554
rect 4773 6502 4783 6554
rect 4807 6502 4837 6554
rect 4837 6502 4849 6554
rect 4849 6502 4863 6554
rect 4887 6502 4901 6554
rect 4901 6502 4913 6554
rect 4913 6502 4943 6554
rect 4967 6502 4977 6554
rect 4977 6502 5023 6554
rect 4727 6500 4783 6502
rect 4807 6500 4863 6502
rect 4887 6500 4943 6502
rect 4967 6500 5023 6502
rect 4256 6010 4312 6012
rect 4336 6010 4392 6012
rect 4416 6010 4472 6012
rect 4496 6010 4552 6012
rect 4256 5958 4302 6010
rect 4302 5958 4312 6010
rect 4336 5958 4366 6010
rect 4366 5958 4378 6010
rect 4378 5958 4392 6010
rect 4416 5958 4430 6010
rect 4430 5958 4442 6010
rect 4442 5958 4472 6010
rect 4496 5958 4506 6010
rect 4506 5958 4552 6010
rect 4256 5956 4312 5958
rect 4336 5956 4392 5958
rect 4416 5956 4472 5958
rect 4496 5956 4552 5958
rect 3784 5466 3840 5468
rect 3864 5466 3920 5468
rect 3944 5466 4000 5468
rect 4024 5466 4080 5468
rect 3784 5414 3830 5466
rect 3830 5414 3840 5466
rect 3864 5414 3894 5466
rect 3894 5414 3906 5466
rect 3906 5414 3920 5466
rect 3944 5414 3958 5466
rect 3958 5414 3970 5466
rect 3970 5414 4000 5466
rect 4024 5414 4034 5466
rect 4034 5414 4080 5466
rect 3784 5412 3840 5414
rect 3864 5412 3920 5414
rect 3944 5412 4000 5414
rect 4024 5412 4080 5414
rect 4727 5466 4783 5468
rect 4807 5466 4863 5468
rect 4887 5466 4943 5468
rect 4967 5466 5023 5468
rect 4727 5414 4773 5466
rect 4773 5414 4783 5466
rect 4807 5414 4837 5466
rect 4837 5414 4849 5466
rect 4849 5414 4863 5466
rect 4887 5414 4901 5466
rect 4901 5414 4913 5466
rect 4913 5414 4943 5466
rect 4967 5414 4977 5466
rect 4977 5414 5023 5466
rect 4727 5412 4783 5414
rect 4807 5412 4863 5414
rect 4887 5412 4943 5414
rect 4967 5412 5023 5414
rect 4256 4922 4312 4924
rect 4336 4922 4392 4924
rect 4416 4922 4472 4924
rect 4496 4922 4552 4924
rect 4256 4870 4302 4922
rect 4302 4870 4312 4922
rect 4336 4870 4366 4922
rect 4366 4870 4378 4922
rect 4378 4870 4392 4922
rect 4416 4870 4430 4922
rect 4430 4870 4442 4922
rect 4442 4870 4472 4922
rect 4496 4870 4506 4922
rect 4506 4870 4552 4922
rect 4256 4868 4312 4870
rect 4336 4868 4392 4870
rect 4416 4868 4472 4870
rect 4496 4868 4552 4870
rect 1898 4378 1954 4380
rect 1978 4378 2034 4380
rect 2058 4378 2114 4380
rect 2138 4378 2194 4380
rect 1898 4326 1944 4378
rect 1944 4326 1954 4378
rect 1978 4326 2008 4378
rect 2008 4326 2020 4378
rect 2020 4326 2034 4378
rect 2058 4326 2072 4378
rect 2072 4326 2084 4378
rect 2084 4326 2114 4378
rect 2138 4326 2148 4378
rect 2148 4326 2194 4378
rect 1898 4324 1954 4326
rect 1978 4324 2034 4326
rect 2058 4324 2114 4326
rect 2138 4324 2194 4326
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 3081 4378 3137 4380
rect 2841 4326 2887 4378
rect 2887 4326 2897 4378
rect 2921 4326 2951 4378
rect 2951 4326 2963 4378
rect 2963 4326 2977 4378
rect 3001 4326 3015 4378
rect 3015 4326 3027 4378
rect 3027 4326 3057 4378
rect 3081 4326 3091 4378
rect 3091 4326 3137 4378
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 3081 4324 3137 4326
rect 3784 4378 3840 4380
rect 3864 4378 3920 4380
rect 3944 4378 4000 4380
rect 4024 4378 4080 4380
rect 3784 4326 3830 4378
rect 3830 4326 3840 4378
rect 3864 4326 3894 4378
rect 3894 4326 3906 4378
rect 3906 4326 3920 4378
rect 3944 4326 3958 4378
rect 3958 4326 3970 4378
rect 3970 4326 4000 4378
rect 4024 4326 4034 4378
rect 4034 4326 4080 4378
rect 3784 4324 3840 4326
rect 3864 4324 3920 4326
rect 3944 4324 4000 4326
rect 4024 4324 4080 4326
rect 4727 4378 4783 4380
rect 4807 4378 4863 4380
rect 4887 4378 4943 4380
rect 4967 4378 5023 4380
rect 4727 4326 4773 4378
rect 4773 4326 4783 4378
rect 4807 4326 4837 4378
rect 4837 4326 4849 4378
rect 4849 4326 4863 4378
rect 4887 4326 4901 4378
rect 4901 4326 4913 4378
rect 4913 4326 4943 4378
rect 4967 4326 4977 4378
rect 4977 4326 5023 4378
rect 4727 4324 4783 4326
rect 4807 4324 4863 4326
rect 4887 4324 4943 4326
rect 4967 4324 5023 4326
rect 4342 4120 4398 4176
rect 1427 3834 1483 3836
rect 1507 3834 1563 3836
rect 1587 3834 1643 3836
rect 1667 3834 1723 3836
rect 1427 3782 1473 3834
rect 1473 3782 1483 3834
rect 1507 3782 1537 3834
rect 1537 3782 1549 3834
rect 1549 3782 1563 3834
rect 1587 3782 1601 3834
rect 1601 3782 1613 3834
rect 1613 3782 1643 3834
rect 1667 3782 1677 3834
rect 1677 3782 1723 3834
rect 1427 3780 1483 3782
rect 1507 3780 1563 3782
rect 1587 3780 1643 3782
rect 1667 3780 1723 3782
rect 2370 3834 2426 3836
rect 2450 3834 2506 3836
rect 2530 3834 2586 3836
rect 2610 3834 2666 3836
rect 2370 3782 2416 3834
rect 2416 3782 2426 3834
rect 2450 3782 2480 3834
rect 2480 3782 2492 3834
rect 2492 3782 2506 3834
rect 2530 3782 2544 3834
rect 2544 3782 2556 3834
rect 2556 3782 2586 3834
rect 2610 3782 2620 3834
rect 2620 3782 2666 3834
rect 2370 3780 2426 3782
rect 2450 3780 2506 3782
rect 2530 3780 2586 3782
rect 2610 3780 2666 3782
rect 3313 3834 3369 3836
rect 3393 3834 3449 3836
rect 3473 3834 3529 3836
rect 3553 3834 3609 3836
rect 3313 3782 3359 3834
rect 3359 3782 3369 3834
rect 3393 3782 3423 3834
rect 3423 3782 3435 3834
rect 3435 3782 3449 3834
rect 3473 3782 3487 3834
rect 3487 3782 3499 3834
rect 3499 3782 3529 3834
rect 3553 3782 3563 3834
rect 3563 3782 3609 3834
rect 3313 3780 3369 3782
rect 3393 3780 3449 3782
rect 3473 3780 3529 3782
rect 3553 3780 3609 3782
rect 1898 3290 1954 3292
rect 1978 3290 2034 3292
rect 2058 3290 2114 3292
rect 2138 3290 2194 3292
rect 1898 3238 1944 3290
rect 1944 3238 1954 3290
rect 1978 3238 2008 3290
rect 2008 3238 2020 3290
rect 2020 3238 2034 3290
rect 2058 3238 2072 3290
rect 2072 3238 2084 3290
rect 2084 3238 2114 3290
rect 2138 3238 2148 3290
rect 2148 3238 2194 3290
rect 1898 3236 1954 3238
rect 1978 3236 2034 3238
rect 2058 3236 2114 3238
rect 2138 3236 2194 3238
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 3081 3290 3137 3292
rect 2841 3238 2887 3290
rect 2887 3238 2897 3290
rect 2921 3238 2951 3290
rect 2951 3238 2963 3290
rect 2963 3238 2977 3290
rect 3001 3238 3015 3290
rect 3015 3238 3027 3290
rect 3027 3238 3057 3290
rect 3081 3238 3091 3290
rect 3091 3238 3137 3290
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 3081 3236 3137 3238
rect 3784 3290 3840 3292
rect 3864 3290 3920 3292
rect 3944 3290 4000 3292
rect 4024 3290 4080 3292
rect 3784 3238 3830 3290
rect 3830 3238 3840 3290
rect 3864 3238 3894 3290
rect 3894 3238 3906 3290
rect 3906 3238 3920 3290
rect 3944 3238 3958 3290
rect 3958 3238 3970 3290
rect 3970 3238 4000 3290
rect 4024 3238 4034 3290
rect 4034 3238 4080 3290
rect 3784 3236 3840 3238
rect 3864 3236 3920 3238
rect 3944 3236 4000 3238
rect 4024 3236 4080 3238
rect 1427 2746 1483 2748
rect 1507 2746 1563 2748
rect 1587 2746 1643 2748
rect 1667 2746 1723 2748
rect 1427 2694 1473 2746
rect 1473 2694 1483 2746
rect 1507 2694 1537 2746
rect 1537 2694 1549 2746
rect 1549 2694 1563 2746
rect 1587 2694 1601 2746
rect 1601 2694 1613 2746
rect 1613 2694 1643 2746
rect 1667 2694 1677 2746
rect 1677 2694 1723 2746
rect 1427 2692 1483 2694
rect 1507 2692 1563 2694
rect 1587 2692 1643 2694
rect 1667 2692 1723 2694
rect 2370 2746 2426 2748
rect 2450 2746 2506 2748
rect 2530 2746 2586 2748
rect 2610 2746 2666 2748
rect 2370 2694 2416 2746
rect 2416 2694 2426 2746
rect 2450 2694 2480 2746
rect 2480 2694 2492 2746
rect 2492 2694 2506 2746
rect 2530 2694 2544 2746
rect 2544 2694 2556 2746
rect 2556 2694 2586 2746
rect 2610 2694 2620 2746
rect 2620 2694 2666 2746
rect 2370 2692 2426 2694
rect 2450 2692 2506 2694
rect 2530 2692 2586 2694
rect 2610 2692 2666 2694
rect 3313 2746 3369 2748
rect 3393 2746 3449 2748
rect 3473 2746 3529 2748
rect 3553 2746 3609 2748
rect 3313 2694 3359 2746
rect 3359 2694 3369 2746
rect 3393 2694 3423 2746
rect 3423 2694 3435 2746
rect 3435 2694 3449 2746
rect 3473 2694 3487 2746
rect 3487 2694 3499 2746
rect 3499 2694 3529 2746
rect 3553 2694 3563 2746
rect 3563 2694 3609 2746
rect 3313 2692 3369 2694
rect 3393 2692 3449 2694
rect 3473 2692 3529 2694
rect 3553 2692 3609 2694
rect 4256 3834 4312 3836
rect 4336 3834 4392 3836
rect 4416 3834 4472 3836
rect 4496 3834 4552 3836
rect 4256 3782 4302 3834
rect 4302 3782 4312 3834
rect 4336 3782 4366 3834
rect 4366 3782 4378 3834
rect 4378 3782 4392 3834
rect 4416 3782 4430 3834
rect 4430 3782 4442 3834
rect 4442 3782 4472 3834
rect 4496 3782 4506 3834
rect 4506 3782 4552 3834
rect 4256 3780 4312 3782
rect 4336 3780 4392 3782
rect 4416 3780 4472 3782
rect 4496 3780 4552 3782
rect 4727 3290 4783 3292
rect 4807 3290 4863 3292
rect 4887 3290 4943 3292
rect 4967 3290 5023 3292
rect 4727 3238 4773 3290
rect 4773 3238 4783 3290
rect 4807 3238 4837 3290
rect 4837 3238 4849 3290
rect 4849 3238 4863 3290
rect 4887 3238 4901 3290
rect 4901 3238 4913 3290
rect 4913 3238 4943 3290
rect 4967 3238 4977 3290
rect 4977 3238 5023 3290
rect 4727 3236 4783 3238
rect 4807 3236 4863 3238
rect 4887 3236 4943 3238
rect 4967 3236 5023 3238
rect 4256 2746 4312 2748
rect 4336 2746 4392 2748
rect 4416 2746 4472 2748
rect 4496 2746 4552 2748
rect 4256 2694 4302 2746
rect 4302 2694 4312 2746
rect 4336 2694 4366 2746
rect 4366 2694 4378 2746
rect 4378 2694 4392 2746
rect 4416 2694 4430 2746
rect 4430 2694 4442 2746
rect 4442 2694 4472 2746
rect 4496 2694 4506 2746
rect 4506 2694 4552 2746
rect 4256 2692 4312 2694
rect 4336 2692 4392 2694
rect 4416 2692 4472 2694
rect 4496 2692 4552 2694
rect 1898 2202 1954 2204
rect 1978 2202 2034 2204
rect 2058 2202 2114 2204
rect 2138 2202 2194 2204
rect 1898 2150 1944 2202
rect 1944 2150 1954 2202
rect 1978 2150 2008 2202
rect 2008 2150 2020 2202
rect 2020 2150 2034 2202
rect 2058 2150 2072 2202
rect 2072 2150 2084 2202
rect 2084 2150 2114 2202
rect 2138 2150 2148 2202
rect 2148 2150 2194 2202
rect 1898 2148 1954 2150
rect 1978 2148 2034 2150
rect 2058 2148 2114 2150
rect 2138 2148 2194 2150
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 3081 2202 3137 2204
rect 2841 2150 2887 2202
rect 2887 2150 2897 2202
rect 2921 2150 2951 2202
rect 2951 2150 2963 2202
rect 2963 2150 2977 2202
rect 3001 2150 3015 2202
rect 3015 2150 3027 2202
rect 3027 2150 3057 2202
rect 3081 2150 3091 2202
rect 3091 2150 3137 2202
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 3081 2148 3137 2150
rect 3784 2202 3840 2204
rect 3864 2202 3920 2204
rect 3944 2202 4000 2204
rect 4024 2202 4080 2204
rect 3784 2150 3830 2202
rect 3830 2150 3840 2202
rect 3864 2150 3894 2202
rect 3894 2150 3906 2202
rect 3906 2150 3920 2202
rect 3944 2150 3958 2202
rect 3958 2150 3970 2202
rect 3970 2150 4000 2202
rect 4024 2150 4034 2202
rect 4034 2150 4080 2202
rect 3784 2148 3840 2150
rect 3864 2148 3920 2150
rect 3944 2148 4000 2150
rect 4024 2148 4080 2150
rect 4727 2202 4783 2204
rect 4807 2202 4863 2204
rect 4887 2202 4943 2204
rect 4967 2202 5023 2204
rect 4727 2150 4773 2202
rect 4773 2150 4783 2202
rect 4807 2150 4837 2202
rect 4837 2150 4849 2202
rect 4849 2150 4863 2202
rect 4887 2150 4901 2202
rect 4901 2150 4913 2202
rect 4913 2150 4943 2202
rect 4967 2150 4977 2202
rect 4977 2150 5023 2202
rect 4727 2148 4783 2150
rect 4807 2148 4863 2150
rect 4887 2148 4943 2150
rect 4967 2148 5023 2150
rect 5078 1400 5134 1456
<< metal3 >>
rect 5073 9618 5139 9621
rect 5200 9618 6000 9648
rect 5073 9616 6000 9618
rect 5073 9560 5078 9616
rect 5134 9560 6000 9616
rect 5073 9558 6000 9560
rect 5073 9555 5139 9558
rect 5200 9528 6000 9558
rect 1888 8736 2204 8737
rect 1888 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2204 8736
rect 1888 8671 2204 8672
rect 2831 8736 3147 8737
rect 2831 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3147 8736
rect 2831 8671 3147 8672
rect 3774 8736 4090 8737
rect 3774 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4090 8736
rect 3774 8671 4090 8672
rect 4717 8736 5033 8737
rect 4717 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5033 8736
rect 4717 8671 5033 8672
rect 0 8258 800 8288
rect 0 8198 1226 8258
rect 0 8168 800 8198
rect 1166 7850 1226 8198
rect 1417 8192 1733 8193
rect 1417 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1733 8192
rect 1417 8127 1733 8128
rect 2360 8192 2676 8193
rect 2360 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2676 8192
rect 2360 8127 2676 8128
rect 3303 8192 3619 8193
rect 3303 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3619 8192
rect 3303 8127 3619 8128
rect 4246 8192 4562 8193
rect 4246 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4562 8192
rect 4246 8127 4562 8128
rect 3693 7850 3759 7853
rect 1166 7848 3759 7850
rect 1166 7792 3698 7848
rect 3754 7792 3759 7848
rect 1166 7790 3759 7792
rect 3693 7787 3759 7790
rect 1888 7648 2204 7649
rect 1888 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2204 7648
rect 1888 7583 2204 7584
rect 2831 7648 3147 7649
rect 2831 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3147 7648
rect 2831 7583 3147 7584
rect 3774 7648 4090 7649
rect 3774 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4090 7648
rect 3774 7583 4090 7584
rect 4717 7648 5033 7649
rect 4717 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5033 7648
rect 4717 7583 5033 7584
rect 1417 7104 1733 7105
rect 1417 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1733 7104
rect 1417 7039 1733 7040
rect 2360 7104 2676 7105
rect 2360 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2676 7104
rect 2360 7039 2676 7040
rect 3303 7104 3619 7105
rect 3303 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3619 7104
rect 3303 7039 3619 7040
rect 4246 7104 4562 7105
rect 4246 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4562 7104
rect 4246 7039 4562 7040
rect 4889 6898 4955 6901
rect 5200 6898 6000 6928
rect 4889 6896 6000 6898
rect 4889 6840 4894 6896
rect 4950 6840 6000 6896
rect 4889 6838 6000 6840
rect 4889 6835 4955 6838
rect 5200 6808 6000 6838
rect 1888 6560 2204 6561
rect 1888 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2204 6560
rect 1888 6495 2204 6496
rect 2831 6560 3147 6561
rect 2831 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3147 6560
rect 2831 6495 3147 6496
rect 3774 6560 4090 6561
rect 3774 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4090 6560
rect 3774 6495 4090 6496
rect 4717 6560 5033 6561
rect 4717 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5033 6560
rect 4717 6495 5033 6496
rect 1417 6016 1733 6017
rect 1417 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1733 6016
rect 1417 5951 1733 5952
rect 2360 6016 2676 6017
rect 2360 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2676 6016
rect 2360 5951 2676 5952
rect 3303 6016 3619 6017
rect 3303 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3619 6016
rect 3303 5951 3619 5952
rect 4246 6016 4562 6017
rect 4246 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4562 6016
rect 4246 5951 4562 5952
rect 1888 5472 2204 5473
rect 1888 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2204 5472
rect 1888 5407 2204 5408
rect 2831 5472 3147 5473
rect 2831 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3147 5472
rect 2831 5407 3147 5408
rect 3774 5472 4090 5473
rect 3774 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4090 5472
rect 3774 5407 4090 5408
rect 4717 5472 5033 5473
rect 4717 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5033 5472
rect 4717 5407 5033 5408
rect 1417 4928 1733 4929
rect 1417 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1733 4928
rect 1417 4863 1733 4864
rect 2360 4928 2676 4929
rect 2360 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2676 4928
rect 2360 4863 2676 4864
rect 3303 4928 3619 4929
rect 3303 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3619 4928
rect 3303 4863 3619 4864
rect 4246 4928 4562 4929
rect 4246 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4562 4928
rect 4246 4863 4562 4864
rect 1888 4384 2204 4385
rect 1888 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2204 4384
rect 1888 4319 2204 4320
rect 2831 4384 3147 4385
rect 2831 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3147 4384
rect 2831 4319 3147 4320
rect 3774 4384 4090 4385
rect 3774 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4090 4384
rect 3774 4319 4090 4320
rect 4717 4384 5033 4385
rect 4717 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5033 4384
rect 4717 4319 5033 4320
rect 4337 4178 4403 4181
rect 5200 4178 6000 4208
rect 4337 4176 6000 4178
rect 4337 4120 4342 4176
rect 4398 4120 6000 4176
rect 4337 4118 6000 4120
rect 4337 4115 4403 4118
rect 5200 4088 6000 4118
rect 1417 3840 1733 3841
rect 1417 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1733 3840
rect 1417 3775 1733 3776
rect 2360 3840 2676 3841
rect 2360 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2676 3840
rect 2360 3775 2676 3776
rect 3303 3840 3619 3841
rect 3303 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3619 3840
rect 3303 3775 3619 3776
rect 4246 3840 4562 3841
rect 4246 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4562 3840
rect 4246 3775 4562 3776
rect 1888 3296 2204 3297
rect 1888 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2204 3296
rect 1888 3231 2204 3232
rect 2831 3296 3147 3297
rect 2831 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3147 3296
rect 2831 3231 3147 3232
rect 3774 3296 4090 3297
rect 3774 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4090 3296
rect 3774 3231 4090 3232
rect 4717 3296 5033 3297
rect 4717 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5033 3296
rect 4717 3231 5033 3232
rect 1417 2752 1733 2753
rect 1417 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1733 2752
rect 1417 2687 1733 2688
rect 2360 2752 2676 2753
rect 2360 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2676 2752
rect 2360 2687 2676 2688
rect 3303 2752 3619 2753
rect 3303 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3619 2752
rect 3303 2687 3619 2688
rect 4246 2752 4562 2753
rect 4246 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4562 2752
rect 4246 2687 4562 2688
rect 1888 2208 2204 2209
rect 1888 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2204 2208
rect 1888 2143 2204 2144
rect 2831 2208 3147 2209
rect 2831 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3147 2208
rect 2831 2143 3147 2144
rect 3774 2208 4090 2209
rect 3774 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4090 2208
rect 3774 2143 4090 2144
rect 4717 2208 5033 2209
rect 4717 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5033 2208
rect 4717 2143 5033 2144
rect 5073 1458 5139 1461
rect 5200 1458 6000 1488
rect 5073 1456 6000 1458
rect 5073 1400 5078 1456
rect 5134 1400 6000 1456
rect 5073 1398 6000 1400
rect 5073 1395 5139 1398
rect 5200 1368 6000 1398
<< via3 >>
rect 1894 8732 1958 8736
rect 1894 8676 1898 8732
rect 1898 8676 1954 8732
rect 1954 8676 1958 8732
rect 1894 8672 1958 8676
rect 1974 8732 2038 8736
rect 1974 8676 1978 8732
rect 1978 8676 2034 8732
rect 2034 8676 2038 8732
rect 1974 8672 2038 8676
rect 2054 8732 2118 8736
rect 2054 8676 2058 8732
rect 2058 8676 2114 8732
rect 2114 8676 2118 8732
rect 2054 8672 2118 8676
rect 2134 8732 2198 8736
rect 2134 8676 2138 8732
rect 2138 8676 2194 8732
rect 2194 8676 2198 8732
rect 2134 8672 2198 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 3077 8732 3141 8736
rect 3077 8676 3081 8732
rect 3081 8676 3137 8732
rect 3137 8676 3141 8732
rect 3077 8672 3141 8676
rect 3780 8732 3844 8736
rect 3780 8676 3784 8732
rect 3784 8676 3840 8732
rect 3840 8676 3844 8732
rect 3780 8672 3844 8676
rect 3860 8732 3924 8736
rect 3860 8676 3864 8732
rect 3864 8676 3920 8732
rect 3920 8676 3924 8732
rect 3860 8672 3924 8676
rect 3940 8732 4004 8736
rect 3940 8676 3944 8732
rect 3944 8676 4000 8732
rect 4000 8676 4004 8732
rect 3940 8672 4004 8676
rect 4020 8732 4084 8736
rect 4020 8676 4024 8732
rect 4024 8676 4080 8732
rect 4080 8676 4084 8732
rect 4020 8672 4084 8676
rect 4723 8732 4787 8736
rect 4723 8676 4727 8732
rect 4727 8676 4783 8732
rect 4783 8676 4787 8732
rect 4723 8672 4787 8676
rect 4803 8732 4867 8736
rect 4803 8676 4807 8732
rect 4807 8676 4863 8732
rect 4863 8676 4867 8732
rect 4803 8672 4867 8676
rect 4883 8732 4947 8736
rect 4883 8676 4887 8732
rect 4887 8676 4943 8732
rect 4943 8676 4947 8732
rect 4883 8672 4947 8676
rect 4963 8732 5027 8736
rect 4963 8676 4967 8732
rect 4967 8676 5023 8732
rect 5023 8676 5027 8732
rect 4963 8672 5027 8676
rect 1423 8188 1487 8192
rect 1423 8132 1427 8188
rect 1427 8132 1483 8188
rect 1483 8132 1487 8188
rect 1423 8128 1487 8132
rect 1503 8188 1567 8192
rect 1503 8132 1507 8188
rect 1507 8132 1563 8188
rect 1563 8132 1567 8188
rect 1503 8128 1567 8132
rect 1583 8188 1647 8192
rect 1583 8132 1587 8188
rect 1587 8132 1643 8188
rect 1643 8132 1647 8188
rect 1583 8128 1647 8132
rect 1663 8188 1727 8192
rect 1663 8132 1667 8188
rect 1667 8132 1723 8188
rect 1723 8132 1727 8188
rect 1663 8128 1727 8132
rect 2366 8188 2430 8192
rect 2366 8132 2370 8188
rect 2370 8132 2426 8188
rect 2426 8132 2430 8188
rect 2366 8128 2430 8132
rect 2446 8188 2510 8192
rect 2446 8132 2450 8188
rect 2450 8132 2506 8188
rect 2506 8132 2510 8188
rect 2446 8128 2510 8132
rect 2526 8188 2590 8192
rect 2526 8132 2530 8188
rect 2530 8132 2586 8188
rect 2586 8132 2590 8188
rect 2526 8128 2590 8132
rect 2606 8188 2670 8192
rect 2606 8132 2610 8188
rect 2610 8132 2666 8188
rect 2666 8132 2670 8188
rect 2606 8128 2670 8132
rect 3309 8188 3373 8192
rect 3309 8132 3313 8188
rect 3313 8132 3369 8188
rect 3369 8132 3373 8188
rect 3309 8128 3373 8132
rect 3389 8188 3453 8192
rect 3389 8132 3393 8188
rect 3393 8132 3449 8188
rect 3449 8132 3453 8188
rect 3389 8128 3453 8132
rect 3469 8188 3533 8192
rect 3469 8132 3473 8188
rect 3473 8132 3529 8188
rect 3529 8132 3533 8188
rect 3469 8128 3533 8132
rect 3549 8188 3613 8192
rect 3549 8132 3553 8188
rect 3553 8132 3609 8188
rect 3609 8132 3613 8188
rect 3549 8128 3613 8132
rect 4252 8188 4316 8192
rect 4252 8132 4256 8188
rect 4256 8132 4312 8188
rect 4312 8132 4316 8188
rect 4252 8128 4316 8132
rect 4332 8188 4396 8192
rect 4332 8132 4336 8188
rect 4336 8132 4392 8188
rect 4392 8132 4396 8188
rect 4332 8128 4396 8132
rect 4412 8188 4476 8192
rect 4412 8132 4416 8188
rect 4416 8132 4472 8188
rect 4472 8132 4476 8188
rect 4412 8128 4476 8132
rect 4492 8188 4556 8192
rect 4492 8132 4496 8188
rect 4496 8132 4552 8188
rect 4552 8132 4556 8188
rect 4492 8128 4556 8132
rect 1894 7644 1958 7648
rect 1894 7588 1898 7644
rect 1898 7588 1954 7644
rect 1954 7588 1958 7644
rect 1894 7584 1958 7588
rect 1974 7644 2038 7648
rect 1974 7588 1978 7644
rect 1978 7588 2034 7644
rect 2034 7588 2038 7644
rect 1974 7584 2038 7588
rect 2054 7644 2118 7648
rect 2054 7588 2058 7644
rect 2058 7588 2114 7644
rect 2114 7588 2118 7644
rect 2054 7584 2118 7588
rect 2134 7644 2198 7648
rect 2134 7588 2138 7644
rect 2138 7588 2194 7644
rect 2194 7588 2198 7644
rect 2134 7584 2198 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 3077 7644 3141 7648
rect 3077 7588 3081 7644
rect 3081 7588 3137 7644
rect 3137 7588 3141 7644
rect 3077 7584 3141 7588
rect 3780 7644 3844 7648
rect 3780 7588 3784 7644
rect 3784 7588 3840 7644
rect 3840 7588 3844 7644
rect 3780 7584 3844 7588
rect 3860 7644 3924 7648
rect 3860 7588 3864 7644
rect 3864 7588 3920 7644
rect 3920 7588 3924 7644
rect 3860 7584 3924 7588
rect 3940 7644 4004 7648
rect 3940 7588 3944 7644
rect 3944 7588 4000 7644
rect 4000 7588 4004 7644
rect 3940 7584 4004 7588
rect 4020 7644 4084 7648
rect 4020 7588 4024 7644
rect 4024 7588 4080 7644
rect 4080 7588 4084 7644
rect 4020 7584 4084 7588
rect 4723 7644 4787 7648
rect 4723 7588 4727 7644
rect 4727 7588 4783 7644
rect 4783 7588 4787 7644
rect 4723 7584 4787 7588
rect 4803 7644 4867 7648
rect 4803 7588 4807 7644
rect 4807 7588 4863 7644
rect 4863 7588 4867 7644
rect 4803 7584 4867 7588
rect 4883 7644 4947 7648
rect 4883 7588 4887 7644
rect 4887 7588 4943 7644
rect 4943 7588 4947 7644
rect 4883 7584 4947 7588
rect 4963 7644 5027 7648
rect 4963 7588 4967 7644
rect 4967 7588 5023 7644
rect 5023 7588 5027 7644
rect 4963 7584 5027 7588
rect 1423 7100 1487 7104
rect 1423 7044 1427 7100
rect 1427 7044 1483 7100
rect 1483 7044 1487 7100
rect 1423 7040 1487 7044
rect 1503 7100 1567 7104
rect 1503 7044 1507 7100
rect 1507 7044 1563 7100
rect 1563 7044 1567 7100
rect 1503 7040 1567 7044
rect 1583 7100 1647 7104
rect 1583 7044 1587 7100
rect 1587 7044 1643 7100
rect 1643 7044 1647 7100
rect 1583 7040 1647 7044
rect 1663 7100 1727 7104
rect 1663 7044 1667 7100
rect 1667 7044 1723 7100
rect 1723 7044 1727 7100
rect 1663 7040 1727 7044
rect 2366 7100 2430 7104
rect 2366 7044 2370 7100
rect 2370 7044 2426 7100
rect 2426 7044 2430 7100
rect 2366 7040 2430 7044
rect 2446 7100 2510 7104
rect 2446 7044 2450 7100
rect 2450 7044 2506 7100
rect 2506 7044 2510 7100
rect 2446 7040 2510 7044
rect 2526 7100 2590 7104
rect 2526 7044 2530 7100
rect 2530 7044 2586 7100
rect 2586 7044 2590 7100
rect 2526 7040 2590 7044
rect 2606 7100 2670 7104
rect 2606 7044 2610 7100
rect 2610 7044 2666 7100
rect 2666 7044 2670 7100
rect 2606 7040 2670 7044
rect 3309 7100 3373 7104
rect 3309 7044 3313 7100
rect 3313 7044 3369 7100
rect 3369 7044 3373 7100
rect 3309 7040 3373 7044
rect 3389 7100 3453 7104
rect 3389 7044 3393 7100
rect 3393 7044 3449 7100
rect 3449 7044 3453 7100
rect 3389 7040 3453 7044
rect 3469 7100 3533 7104
rect 3469 7044 3473 7100
rect 3473 7044 3529 7100
rect 3529 7044 3533 7100
rect 3469 7040 3533 7044
rect 3549 7100 3613 7104
rect 3549 7044 3553 7100
rect 3553 7044 3609 7100
rect 3609 7044 3613 7100
rect 3549 7040 3613 7044
rect 4252 7100 4316 7104
rect 4252 7044 4256 7100
rect 4256 7044 4312 7100
rect 4312 7044 4316 7100
rect 4252 7040 4316 7044
rect 4332 7100 4396 7104
rect 4332 7044 4336 7100
rect 4336 7044 4392 7100
rect 4392 7044 4396 7100
rect 4332 7040 4396 7044
rect 4412 7100 4476 7104
rect 4412 7044 4416 7100
rect 4416 7044 4472 7100
rect 4472 7044 4476 7100
rect 4412 7040 4476 7044
rect 4492 7100 4556 7104
rect 4492 7044 4496 7100
rect 4496 7044 4552 7100
rect 4552 7044 4556 7100
rect 4492 7040 4556 7044
rect 1894 6556 1958 6560
rect 1894 6500 1898 6556
rect 1898 6500 1954 6556
rect 1954 6500 1958 6556
rect 1894 6496 1958 6500
rect 1974 6556 2038 6560
rect 1974 6500 1978 6556
rect 1978 6500 2034 6556
rect 2034 6500 2038 6556
rect 1974 6496 2038 6500
rect 2054 6556 2118 6560
rect 2054 6500 2058 6556
rect 2058 6500 2114 6556
rect 2114 6500 2118 6556
rect 2054 6496 2118 6500
rect 2134 6556 2198 6560
rect 2134 6500 2138 6556
rect 2138 6500 2194 6556
rect 2194 6500 2198 6556
rect 2134 6496 2198 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 3077 6556 3141 6560
rect 3077 6500 3081 6556
rect 3081 6500 3137 6556
rect 3137 6500 3141 6556
rect 3077 6496 3141 6500
rect 3780 6556 3844 6560
rect 3780 6500 3784 6556
rect 3784 6500 3840 6556
rect 3840 6500 3844 6556
rect 3780 6496 3844 6500
rect 3860 6556 3924 6560
rect 3860 6500 3864 6556
rect 3864 6500 3920 6556
rect 3920 6500 3924 6556
rect 3860 6496 3924 6500
rect 3940 6556 4004 6560
rect 3940 6500 3944 6556
rect 3944 6500 4000 6556
rect 4000 6500 4004 6556
rect 3940 6496 4004 6500
rect 4020 6556 4084 6560
rect 4020 6500 4024 6556
rect 4024 6500 4080 6556
rect 4080 6500 4084 6556
rect 4020 6496 4084 6500
rect 4723 6556 4787 6560
rect 4723 6500 4727 6556
rect 4727 6500 4783 6556
rect 4783 6500 4787 6556
rect 4723 6496 4787 6500
rect 4803 6556 4867 6560
rect 4803 6500 4807 6556
rect 4807 6500 4863 6556
rect 4863 6500 4867 6556
rect 4803 6496 4867 6500
rect 4883 6556 4947 6560
rect 4883 6500 4887 6556
rect 4887 6500 4943 6556
rect 4943 6500 4947 6556
rect 4883 6496 4947 6500
rect 4963 6556 5027 6560
rect 4963 6500 4967 6556
rect 4967 6500 5023 6556
rect 5023 6500 5027 6556
rect 4963 6496 5027 6500
rect 1423 6012 1487 6016
rect 1423 5956 1427 6012
rect 1427 5956 1483 6012
rect 1483 5956 1487 6012
rect 1423 5952 1487 5956
rect 1503 6012 1567 6016
rect 1503 5956 1507 6012
rect 1507 5956 1563 6012
rect 1563 5956 1567 6012
rect 1503 5952 1567 5956
rect 1583 6012 1647 6016
rect 1583 5956 1587 6012
rect 1587 5956 1643 6012
rect 1643 5956 1647 6012
rect 1583 5952 1647 5956
rect 1663 6012 1727 6016
rect 1663 5956 1667 6012
rect 1667 5956 1723 6012
rect 1723 5956 1727 6012
rect 1663 5952 1727 5956
rect 2366 6012 2430 6016
rect 2366 5956 2370 6012
rect 2370 5956 2426 6012
rect 2426 5956 2430 6012
rect 2366 5952 2430 5956
rect 2446 6012 2510 6016
rect 2446 5956 2450 6012
rect 2450 5956 2506 6012
rect 2506 5956 2510 6012
rect 2446 5952 2510 5956
rect 2526 6012 2590 6016
rect 2526 5956 2530 6012
rect 2530 5956 2586 6012
rect 2586 5956 2590 6012
rect 2526 5952 2590 5956
rect 2606 6012 2670 6016
rect 2606 5956 2610 6012
rect 2610 5956 2666 6012
rect 2666 5956 2670 6012
rect 2606 5952 2670 5956
rect 3309 6012 3373 6016
rect 3309 5956 3313 6012
rect 3313 5956 3369 6012
rect 3369 5956 3373 6012
rect 3309 5952 3373 5956
rect 3389 6012 3453 6016
rect 3389 5956 3393 6012
rect 3393 5956 3449 6012
rect 3449 5956 3453 6012
rect 3389 5952 3453 5956
rect 3469 6012 3533 6016
rect 3469 5956 3473 6012
rect 3473 5956 3529 6012
rect 3529 5956 3533 6012
rect 3469 5952 3533 5956
rect 3549 6012 3613 6016
rect 3549 5956 3553 6012
rect 3553 5956 3609 6012
rect 3609 5956 3613 6012
rect 3549 5952 3613 5956
rect 4252 6012 4316 6016
rect 4252 5956 4256 6012
rect 4256 5956 4312 6012
rect 4312 5956 4316 6012
rect 4252 5952 4316 5956
rect 4332 6012 4396 6016
rect 4332 5956 4336 6012
rect 4336 5956 4392 6012
rect 4392 5956 4396 6012
rect 4332 5952 4396 5956
rect 4412 6012 4476 6016
rect 4412 5956 4416 6012
rect 4416 5956 4472 6012
rect 4472 5956 4476 6012
rect 4412 5952 4476 5956
rect 4492 6012 4556 6016
rect 4492 5956 4496 6012
rect 4496 5956 4552 6012
rect 4552 5956 4556 6012
rect 4492 5952 4556 5956
rect 1894 5468 1958 5472
rect 1894 5412 1898 5468
rect 1898 5412 1954 5468
rect 1954 5412 1958 5468
rect 1894 5408 1958 5412
rect 1974 5468 2038 5472
rect 1974 5412 1978 5468
rect 1978 5412 2034 5468
rect 2034 5412 2038 5468
rect 1974 5408 2038 5412
rect 2054 5468 2118 5472
rect 2054 5412 2058 5468
rect 2058 5412 2114 5468
rect 2114 5412 2118 5468
rect 2054 5408 2118 5412
rect 2134 5468 2198 5472
rect 2134 5412 2138 5468
rect 2138 5412 2194 5468
rect 2194 5412 2198 5468
rect 2134 5408 2198 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 3077 5468 3141 5472
rect 3077 5412 3081 5468
rect 3081 5412 3137 5468
rect 3137 5412 3141 5468
rect 3077 5408 3141 5412
rect 3780 5468 3844 5472
rect 3780 5412 3784 5468
rect 3784 5412 3840 5468
rect 3840 5412 3844 5468
rect 3780 5408 3844 5412
rect 3860 5468 3924 5472
rect 3860 5412 3864 5468
rect 3864 5412 3920 5468
rect 3920 5412 3924 5468
rect 3860 5408 3924 5412
rect 3940 5468 4004 5472
rect 3940 5412 3944 5468
rect 3944 5412 4000 5468
rect 4000 5412 4004 5468
rect 3940 5408 4004 5412
rect 4020 5468 4084 5472
rect 4020 5412 4024 5468
rect 4024 5412 4080 5468
rect 4080 5412 4084 5468
rect 4020 5408 4084 5412
rect 4723 5468 4787 5472
rect 4723 5412 4727 5468
rect 4727 5412 4783 5468
rect 4783 5412 4787 5468
rect 4723 5408 4787 5412
rect 4803 5468 4867 5472
rect 4803 5412 4807 5468
rect 4807 5412 4863 5468
rect 4863 5412 4867 5468
rect 4803 5408 4867 5412
rect 4883 5468 4947 5472
rect 4883 5412 4887 5468
rect 4887 5412 4943 5468
rect 4943 5412 4947 5468
rect 4883 5408 4947 5412
rect 4963 5468 5027 5472
rect 4963 5412 4967 5468
rect 4967 5412 5023 5468
rect 5023 5412 5027 5468
rect 4963 5408 5027 5412
rect 1423 4924 1487 4928
rect 1423 4868 1427 4924
rect 1427 4868 1483 4924
rect 1483 4868 1487 4924
rect 1423 4864 1487 4868
rect 1503 4924 1567 4928
rect 1503 4868 1507 4924
rect 1507 4868 1563 4924
rect 1563 4868 1567 4924
rect 1503 4864 1567 4868
rect 1583 4924 1647 4928
rect 1583 4868 1587 4924
rect 1587 4868 1643 4924
rect 1643 4868 1647 4924
rect 1583 4864 1647 4868
rect 1663 4924 1727 4928
rect 1663 4868 1667 4924
rect 1667 4868 1723 4924
rect 1723 4868 1727 4924
rect 1663 4864 1727 4868
rect 2366 4924 2430 4928
rect 2366 4868 2370 4924
rect 2370 4868 2426 4924
rect 2426 4868 2430 4924
rect 2366 4864 2430 4868
rect 2446 4924 2510 4928
rect 2446 4868 2450 4924
rect 2450 4868 2506 4924
rect 2506 4868 2510 4924
rect 2446 4864 2510 4868
rect 2526 4924 2590 4928
rect 2526 4868 2530 4924
rect 2530 4868 2586 4924
rect 2586 4868 2590 4924
rect 2526 4864 2590 4868
rect 2606 4924 2670 4928
rect 2606 4868 2610 4924
rect 2610 4868 2666 4924
rect 2666 4868 2670 4924
rect 2606 4864 2670 4868
rect 3309 4924 3373 4928
rect 3309 4868 3313 4924
rect 3313 4868 3369 4924
rect 3369 4868 3373 4924
rect 3309 4864 3373 4868
rect 3389 4924 3453 4928
rect 3389 4868 3393 4924
rect 3393 4868 3449 4924
rect 3449 4868 3453 4924
rect 3389 4864 3453 4868
rect 3469 4924 3533 4928
rect 3469 4868 3473 4924
rect 3473 4868 3529 4924
rect 3529 4868 3533 4924
rect 3469 4864 3533 4868
rect 3549 4924 3613 4928
rect 3549 4868 3553 4924
rect 3553 4868 3609 4924
rect 3609 4868 3613 4924
rect 3549 4864 3613 4868
rect 4252 4924 4316 4928
rect 4252 4868 4256 4924
rect 4256 4868 4312 4924
rect 4312 4868 4316 4924
rect 4252 4864 4316 4868
rect 4332 4924 4396 4928
rect 4332 4868 4336 4924
rect 4336 4868 4392 4924
rect 4392 4868 4396 4924
rect 4332 4864 4396 4868
rect 4412 4924 4476 4928
rect 4412 4868 4416 4924
rect 4416 4868 4472 4924
rect 4472 4868 4476 4924
rect 4412 4864 4476 4868
rect 4492 4924 4556 4928
rect 4492 4868 4496 4924
rect 4496 4868 4552 4924
rect 4552 4868 4556 4924
rect 4492 4864 4556 4868
rect 1894 4380 1958 4384
rect 1894 4324 1898 4380
rect 1898 4324 1954 4380
rect 1954 4324 1958 4380
rect 1894 4320 1958 4324
rect 1974 4380 2038 4384
rect 1974 4324 1978 4380
rect 1978 4324 2034 4380
rect 2034 4324 2038 4380
rect 1974 4320 2038 4324
rect 2054 4380 2118 4384
rect 2054 4324 2058 4380
rect 2058 4324 2114 4380
rect 2114 4324 2118 4380
rect 2054 4320 2118 4324
rect 2134 4380 2198 4384
rect 2134 4324 2138 4380
rect 2138 4324 2194 4380
rect 2194 4324 2198 4380
rect 2134 4320 2198 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 3077 4380 3141 4384
rect 3077 4324 3081 4380
rect 3081 4324 3137 4380
rect 3137 4324 3141 4380
rect 3077 4320 3141 4324
rect 3780 4380 3844 4384
rect 3780 4324 3784 4380
rect 3784 4324 3840 4380
rect 3840 4324 3844 4380
rect 3780 4320 3844 4324
rect 3860 4380 3924 4384
rect 3860 4324 3864 4380
rect 3864 4324 3920 4380
rect 3920 4324 3924 4380
rect 3860 4320 3924 4324
rect 3940 4380 4004 4384
rect 3940 4324 3944 4380
rect 3944 4324 4000 4380
rect 4000 4324 4004 4380
rect 3940 4320 4004 4324
rect 4020 4380 4084 4384
rect 4020 4324 4024 4380
rect 4024 4324 4080 4380
rect 4080 4324 4084 4380
rect 4020 4320 4084 4324
rect 4723 4380 4787 4384
rect 4723 4324 4727 4380
rect 4727 4324 4783 4380
rect 4783 4324 4787 4380
rect 4723 4320 4787 4324
rect 4803 4380 4867 4384
rect 4803 4324 4807 4380
rect 4807 4324 4863 4380
rect 4863 4324 4867 4380
rect 4803 4320 4867 4324
rect 4883 4380 4947 4384
rect 4883 4324 4887 4380
rect 4887 4324 4943 4380
rect 4943 4324 4947 4380
rect 4883 4320 4947 4324
rect 4963 4380 5027 4384
rect 4963 4324 4967 4380
rect 4967 4324 5023 4380
rect 5023 4324 5027 4380
rect 4963 4320 5027 4324
rect 1423 3836 1487 3840
rect 1423 3780 1427 3836
rect 1427 3780 1483 3836
rect 1483 3780 1487 3836
rect 1423 3776 1487 3780
rect 1503 3836 1567 3840
rect 1503 3780 1507 3836
rect 1507 3780 1563 3836
rect 1563 3780 1567 3836
rect 1503 3776 1567 3780
rect 1583 3836 1647 3840
rect 1583 3780 1587 3836
rect 1587 3780 1643 3836
rect 1643 3780 1647 3836
rect 1583 3776 1647 3780
rect 1663 3836 1727 3840
rect 1663 3780 1667 3836
rect 1667 3780 1723 3836
rect 1723 3780 1727 3836
rect 1663 3776 1727 3780
rect 2366 3836 2430 3840
rect 2366 3780 2370 3836
rect 2370 3780 2426 3836
rect 2426 3780 2430 3836
rect 2366 3776 2430 3780
rect 2446 3836 2510 3840
rect 2446 3780 2450 3836
rect 2450 3780 2506 3836
rect 2506 3780 2510 3836
rect 2446 3776 2510 3780
rect 2526 3836 2590 3840
rect 2526 3780 2530 3836
rect 2530 3780 2586 3836
rect 2586 3780 2590 3836
rect 2526 3776 2590 3780
rect 2606 3836 2670 3840
rect 2606 3780 2610 3836
rect 2610 3780 2666 3836
rect 2666 3780 2670 3836
rect 2606 3776 2670 3780
rect 3309 3836 3373 3840
rect 3309 3780 3313 3836
rect 3313 3780 3369 3836
rect 3369 3780 3373 3836
rect 3309 3776 3373 3780
rect 3389 3836 3453 3840
rect 3389 3780 3393 3836
rect 3393 3780 3449 3836
rect 3449 3780 3453 3836
rect 3389 3776 3453 3780
rect 3469 3836 3533 3840
rect 3469 3780 3473 3836
rect 3473 3780 3529 3836
rect 3529 3780 3533 3836
rect 3469 3776 3533 3780
rect 3549 3836 3613 3840
rect 3549 3780 3553 3836
rect 3553 3780 3609 3836
rect 3609 3780 3613 3836
rect 3549 3776 3613 3780
rect 4252 3836 4316 3840
rect 4252 3780 4256 3836
rect 4256 3780 4312 3836
rect 4312 3780 4316 3836
rect 4252 3776 4316 3780
rect 4332 3836 4396 3840
rect 4332 3780 4336 3836
rect 4336 3780 4392 3836
rect 4392 3780 4396 3836
rect 4332 3776 4396 3780
rect 4412 3836 4476 3840
rect 4412 3780 4416 3836
rect 4416 3780 4472 3836
rect 4472 3780 4476 3836
rect 4412 3776 4476 3780
rect 4492 3836 4556 3840
rect 4492 3780 4496 3836
rect 4496 3780 4552 3836
rect 4552 3780 4556 3836
rect 4492 3776 4556 3780
rect 1894 3292 1958 3296
rect 1894 3236 1898 3292
rect 1898 3236 1954 3292
rect 1954 3236 1958 3292
rect 1894 3232 1958 3236
rect 1974 3292 2038 3296
rect 1974 3236 1978 3292
rect 1978 3236 2034 3292
rect 2034 3236 2038 3292
rect 1974 3232 2038 3236
rect 2054 3292 2118 3296
rect 2054 3236 2058 3292
rect 2058 3236 2114 3292
rect 2114 3236 2118 3292
rect 2054 3232 2118 3236
rect 2134 3292 2198 3296
rect 2134 3236 2138 3292
rect 2138 3236 2194 3292
rect 2194 3236 2198 3292
rect 2134 3232 2198 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 3077 3292 3141 3296
rect 3077 3236 3081 3292
rect 3081 3236 3137 3292
rect 3137 3236 3141 3292
rect 3077 3232 3141 3236
rect 3780 3292 3844 3296
rect 3780 3236 3784 3292
rect 3784 3236 3840 3292
rect 3840 3236 3844 3292
rect 3780 3232 3844 3236
rect 3860 3292 3924 3296
rect 3860 3236 3864 3292
rect 3864 3236 3920 3292
rect 3920 3236 3924 3292
rect 3860 3232 3924 3236
rect 3940 3292 4004 3296
rect 3940 3236 3944 3292
rect 3944 3236 4000 3292
rect 4000 3236 4004 3292
rect 3940 3232 4004 3236
rect 4020 3292 4084 3296
rect 4020 3236 4024 3292
rect 4024 3236 4080 3292
rect 4080 3236 4084 3292
rect 4020 3232 4084 3236
rect 4723 3292 4787 3296
rect 4723 3236 4727 3292
rect 4727 3236 4783 3292
rect 4783 3236 4787 3292
rect 4723 3232 4787 3236
rect 4803 3292 4867 3296
rect 4803 3236 4807 3292
rect 4807 3236 4863 3292
rect 4863 3236 4867 3292
rect 4803 3232 4867 3236
rect 4883 3292 4947 3296
rect 4883 3236 4887 3292
rect 4887 3236 4943 3292
rect 4943 3236 4947 3292
rect 4883 3232 4947 3236
rect 4963 3292 5027 3296
rect 4963 3236 4967 3292
rect 4967 3236 5023 3292
rect 5023 3236 5027 3292
rect 4963 3232 5027 3236
rect 1423 2748 1487 2752
rect 1423 2692 1427 2748
rect 1427 2692 1483 2748
rect 1483 2692 1487 2748
rect 1423 2688 1487 2692
rect 1503 2748 1567 2752
rect 1503 2692 1507 2748
rect 1507 2692 1563 2748
rect 1563 2692 1567 2748
rect 1503 2688 1567 2692
rect 1583 2748 1647 2752
rect 1583 2692 1587 2748
rect 1587 2692 1643 2748
rect 1643 2692 1647 2748
rect 1583 2688 1647 2692
rect 1663 2748 1727 2752
rect 1663 2692 1667 2748
rect 1667 2692 1723 2748
rect 1723 2692 1727 2748
rect 1663 2688 1727 2692
rect 2366 2748 2430 2752
rect 2366 2692 2370 2748
rect 2370 2692 2426 2748
rect 2426 2692 2430 2748
rect 2366 2688 2430 2692
rect 2446 2748 2510 2752
rect 2446 2692 2450 2748
rect 2450 2692 2506 2748
rect 2506 2692 2510 2748
rect 2446 2688 2510 2692
rect 2526 2748 2590 2752
rect 2526 2692 2530 2748
rect 2530 2692 2586 2748
rect 2586 2692 2590 2748
rect 2526 2688 2590 2692
rect 2606 2748 2670 2752
rect 2606 2692 2610 2748
rect 2610 2692 2666 2748
rect 2666 2692 2670 2748
rect 2606 2688 2670 2692
rect 3309 2748 3373 2752
rect 3309 2692 3313 2748
rect 3313 2692 3369 2748
rect 3369 2692 3373 2748
rect 3309 2688 3373 2692
rect 3389 2748 3453 2752
rect 3389 2692 3393 2748
rect 3393 2692 3449 2748
rect 3449 2692 3453 2748
rect 3389 2688 3453 2692
rect 3469 2748 3533 2752
rect 3469 2692 3473 2748
rect 3473 2692 3529 2748
rect 3529 2692 3533 2748
rect 3469 2688 3533 2692
rect 3549 2748 3613 2752
rect 3549 2692 3553 2748
rect 3553 2692 3609 2748
rect 3609 2692 3613 2748
rect 3549 2688 3613 2692
rect 4252 2748 4316 2752
rect 4252 2692 4256 2748
rect 4256 2692 4312 2748
rect 4312 2692 4316 2748
rect 4252 2688 4316 2692
rect 4332 2748 4396 2752
rect 4332 2692 4336 2748
rect 4336 2692 4392 2748
rect 4392 2692 4396 2748
rect 4332 2688 4396 2692
rect 4412 2748 4476 2752
rect 4412 2692 4416 2748
rect 4416 2692 4472 2748
rect 4472 2692 4476 2748
rect 4412 2688 4476 2692
rect 4492 2748 4556 2752
rect 4492 2692 4496 2748
rect 4496 2692 4552 2748
rect 4552 2692 4556 2748
rect 4492 2688 4556 2692
rect 1894 2204 1958 2208
rect 1894 2148 1898 2204
rect 1898 2148 1954 2204
rect 1954 2148 1958 2204
rect 1894 2144 1958 2148
rect 1974 2204 2038 2208
rect 1974 2148 1978 2204
rect 1978 2148 2034 2204
rect 2034 2148 2038 2204
rect 1974 2144 2038 2148
rect 2054 2204 2118 2208
rect 2054 2148 2058 2204
rect 2058 2148 2114 2204
rect 2114 2148 2118 2204
rect 2054 2144 2118 2148
rect 2134 2204 2198 2208
rect 2134 2148 2138 2204
rect 2138 2148 2194 2204
rect 2194 2148 2198 2204
rect 2134 2144 2198 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 3077 2204 3141 2208
rect 3077 2148 3081 2204
rect 3081 2148 3137 2204
rect 3137 2148 3141 2204
rect 3077 2144 3141 2148
rect 3780 2204 3844 2208
rect 3780 2148 3784 2204
rect 3784 2148 3840 2204
rect 3840 2148 3844 2204
rect 3780 2144 3844 2148
rect 3860 2204 3924 2208
rect 3860 2148 3864 2204
rect 3864 2148 3920 2204
rect 3920 2148 3924 2204
rect 3860 2144 3924 2148
rect 3940 2204 4004 2208
rect 3940 2148 3944 2204
rect 3944 2148 4000 2204
rect 4000 2148 4004 2204
rect 3940 2144 4004 2148
rect 4020 2204 4084 2208
rect 4020 2148 4024 2204
rect 4024 2148 4080 2204
rect 4080 2148 4084 2204
rect 4020 2144 4084 2148
rect 4723 2204 4787 2208
rect 4723 2148 4727 2204
rect 4727 2148 4783 2204
rect 4783 2148 4787 2204
rect 4723 2144 4787 2148
rect 4803 2204 4867 2208
rect 4803 2148 4807 2204
rect 4807 2148 4863 2204
rect 4863 2148 4867 2204
rect 4803 2144 4867 2148
rect 4883 2204 4947 2208
rect 4883 2148 4887 2204
rect 4887 2148 4943 2204
rect 4943 2148 4947 2204
rect 4883 2144 4947 2148
rect 4963 2204 5027 2208
rect 4963 2148 4967 2204
rect 4967 2148 5023 2204
rect 5023 2148 5027 2204
rect 4963 2144 5027 2148
<< metal4 >>
rect 1415 8192 1735 8752
rect 1415 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1735 8192
rect 1415 7104 1735 8128
rect 1415 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1735 7104
rect 1415 6016 1735 7040
rect 1415 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1735 6016
rect 1415 4928 1735 5952
rect 1415 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1735 4928
rect 1415 3840 1735 4864
rect 1415 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1735 3840
rect 1415 2752 1735 3776
rect 1415 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1735 2752
rect 1415 2128 1735 2688
rect 1886 8736 2206 8752
rect 1886 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2206 8736
rect 1886 7648 2206 8672
rect 1886 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2206 7648
rect 1886 6560 2206 7584
rect 1886 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2206 6560
rect 1886 5472 2206 6496
rect 1886 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2206 5472
rect 1886 4384 2206 5408
rect 1886 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2206 4384
rect 1886 3296 2206 4320
rect 1886 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2206 3296
rect 1886 2208 2206 3232
rect 1886 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2206 2208
rect 1886 2128 2206 2144
rect 2358 8192 2678 8752
rect 2358 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2678 8192
rect 2358 7104 2678 8128
rect 2358 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2678 7104
rect 2358 6016 2678 7040
rect 2358 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2678 6016
rect 2358 4928 2678 5952
rect 2358 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2678 4928
rect 2358 3840 2678 4864
rect 2358 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2678 3840
rect 2358 2752 2678 3776
rect 2358 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2678 2752
rect 2358 2128 2678 2688
rect 2829 8736 3149 8752
rect 2829 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3149 8736
rect 2829 7648 3149 8672
rect 2829 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3149 7648
rect 2829 6560 3149 7584
rect 2829 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3149 6560
rect 2829 5472 3149 6496
rect 2829 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3149 5472
rect 2829 4384 3149 5408
rect 2829 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3149 4384
rect 2829 3296 3149 4320
rect 2829 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3149 3296
rect 2829 2208 3149 3232
rect 2829 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3149 2208
rect 2829 2128 3149 2144
rect 3301 8192 3621 8752
rect 3301 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3621 8192
rect 3301 7104 3621 8128
rect 3301 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3621 7104
rect 3301 6016 3621 7040
rect 3301 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3621 6016
rect 3301 4928 3621 5952
rect 3301 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3621 4928
rect 3301 3840 3621 4864
rect 3301 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3621 3840
rect 3301 2752 3621 3776
rect 3301 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3621 2752
rect 3301 2128 3621 2688
rect 3772 8736 4092 8752
rect 3772 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4092 8736
rect 3772 7648 4092 8672
rect 3772 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4092 7648
rect 3772 6560 4092 7584
rect 3772 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4092 6560
rect 3772 5472 4092 6496
rect 3772 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4092 5472
rect 3772 4384 4092 5408
rect 3772 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4092 4384
rect 3772 3296 4092 4320
rect 3772 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4092 3296
rect 3772 2208 4092 3232
rect 3772 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4092 2208
rect 3772 2128 4092 2144
rect 4244 8192 4564 8752
rect 4244 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4564 8192
rect 4244 7104 4564 8128
rect 4244 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4564 7104
rect 4244 6016 4564 7040
rect 4244 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4564 6016
rect 4244 4928 4564 5952
rect 4244 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4564 4928
rect 4244 3840 4564 4864
rect 4244 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4564 3840
rect 4244 2752 4564 3776
rect 4244 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4564 2752
rect 4244 2128 4564 2688
rect 4715 8736 5035 8752
rect 4715 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5035 8736
rect 4715 7648 5035 8672
rect 4715 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5035 7648
rect 4715 6560 5035 7584
rect 4715 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5035 6560
rect 4715 5472 5035 6496
rect 4715 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5035 5472
rect 4715 4384 5035 5408
rect 4715 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5035 4384
rect 4715 3296 5035 4320
rect 4715 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5035 3296
rect 4715 2208 5035 3232
rect 4715 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5035 2208
rect 4715 2128 5035 2144
use sky130_fd_sc_hd__dfxtp_1  _0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 1688980957
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1688980957
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_35
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_23
timestamp 1688980957
transform 1 0 3220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  grid_io_top_out_5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 5200 6808 6000 6928 0 FreeSans 480 0 0 0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal tristate
flabel metal3 s 5200 9528 6000 9648 0 FreeSans 480 0 0 0 bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 1 nsew signal input
flabel metal3 s 5200 1368 6000 1488 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 5200 4088 6000 4208 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal2 s 2962 10200 3018 11000 0 FreeSans 224 90 0 0 gfpga_pad_GPIO_PAD
port 4 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 prog_clk
port 5 nsew signal input
flabel metal4 s 1415 2128 1735 8752 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 2358 2128 2678 8752 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 3301 2128 3621 8752 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 4244 2128 4564 8752 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 1886 2128 2206 8752 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 2829 2128 3149 8752 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 3772 2128 4092 8752 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 4715 2128 5035 8752 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
rlabel metal1 2990 8160 2990 8160 0 vdd
rlabel via1 3069 8704 3069 8704 0 vss
rlabel metal1 4830 8466 4830 8466 0 bottom_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4830 2414 4830 2414 0 ccff_head
rlabel metal2 4370 4301 4370 4301 0 ccff_tail
rlabel metal1 3220 8602 3220 8602 0 gfpga_pad_GPIO_PAD
rlabel metal1 3588 7378 3588 7378 0 net1
rlabel metal1 4278 2618 4278 2618 0 net2
rlabel metal2 4554 4420 4554 4420 0 net3
rlabel metal1 3312 7514 3312 7514 0 net4
rlabel metal1 4738 7174 4738 7174 0 net5
rlabel metal3 935 8228 935 8228 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 6000 11000
<< end >>
