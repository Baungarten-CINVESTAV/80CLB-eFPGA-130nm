magic
tech sky130A
magscale 1 2
timestamp 1708121278
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 934 1640 29048 27872
<< metal2 >>
rect 3790 29200 3846 30000
rect 11242 29200 11298 30000
rect 18694 29200 18750 30000
rect 26146 29200 26202 30000
rect 3790 0 3846 800
rect 11242 0 11298 800
rect 18694 0 18750 800
rect 26146 0 26202 800
<< obsm2 >>
rect 938 29144 3734 29200
rect 3902 29144 11186 29200
rect 11354 29144 18638 29200
rect 18806 29144 26090 29200
rect 26258 29144 29042 29200
rect 938 856 29042 29144
rect 938 734 3734 856
rect 3902 734 11186 856
rect 11354 734 18638 856
rect 18806 734 26090 856
rect 26258 734 29042 856
<< metal3 >>
rect 0 27208 800 27328
rect 29200 26936 30000 27056
rect 0 23672 800 23792
rect 29200 22040 30000 22160
rect 0 20136 800 20256
rect 29200 17144 30000 17264
rect 0 16600 800 16720
rect 0 13064 800 13184
rect 29200 12248 30000 12368
rect 0 9528 800 9648
rect 29200 7352 30000 7472
rect 0 5992 800 6112
rect 29200 2456 30000 2576
<< obsm3 >>
rect 800 27408 29200 27777
rect 880 27136 29200 27408
rect 880 27128 29120 27136
rect 800 26856 29120 27128
rect 800 23872 29200 26856
rect 880 23592 29200 23872
rect 800 22240 29200 23592
rect 800 21960 29120 22240
rect 800 20336 29200 21960
rect 880 20056 29200 20336
rect 800 17344 29200 20056
rect 800 17064 29120 17344
rect 800 16800 29200 17064
rect 880 16520 29200 16800
rect 800 13264 29200 16520
rect 880 12984 29200 13264
rect 800 12448 29200 12984
rect 800 12168 29120 12448
rect 800 9728 29200 12168
rect 880 9448 29200 9728
rect 800 7552 29200 9448
rect 800 7272 29120 7552
rect 800 6192 29200 7272
rect 880 5912 29200 6192
rect 800 2656 29200 5912
rect 800 2376 29120 2656
rect 800 1940 29200 2376
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< obsm4 >>
rect 4843 2048 7810 18053
rect 8290 2048 11283 18053
rect 11763 2048 14756 18053
rect 15236 2048 18229 18053
rect 18709 2048 21702 18053
rect 22182 2048 25175 18053
rect 25655 2048 26069 18053
rect 4843 1939 26069 2048
<< labels >>
rlabel metal2 s 3790 0 3846 800 6 bottom_width_0_height_0_subtile_0__pin_I_2_
port 1 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 bottom_width_0_height_0_subtile_0__pin_I_6_
port 2 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 bottom_width_0_height_0_subtile_0__pin_O_0_
port 3 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 bottom_width_0_height_0_subtile_0__pin_clk_0_
port 4 nsew signal input
rlabel metal3 s 29200 22040 30000 22160 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 29200 26936 30000 27056 6 ccff_tail
port 6 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 clk
port 7 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 left_width_0_height_0_subtile_0__pin_I_3_
port 8 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 left_width_0_height_0_subtile_0__pin_I_7_
port 9 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 left_width_0_height_0_subtile_0__pin_O_1_
port 10 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 prog_clk
port 11 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 reset
port 12 nsew signal input
rlabel metal3 s 29200 2456 30000 2576 6 right_width_0_height_0_subtile_0__pin_I_1_
port 13 nsew signal input
rlabel metal3 s 29200 7352 30000 7472 6 right_width_0_height_0_subtile_0__pin_I_5_
port 14 nsew signal input
rlabel metal3 s 29200 12248 30000 12368 6 right_width_0_height_0_subtile_0__pin_I_9_
port 15 nsew signal input
rlabel metal3 s 29200 17144 30000 17264 6 right_width_0_height_0_subtile_0__pin_O_3_
port 16 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 set
port 17 nsew signal input
rlabel metal2 s 3790 29200 3846 30000 6 top_width_0_height_0_subtile_0__pin_I_0_
port 18 nsew signal input
rlabel metal2 s 11242 29200 11298 30000 6 top_width_0_height_0_subtile_0__pin_I_4_
port 19 nsew signal input
rlabel metal2 s 18694 29200 18750 30000 6 top_width_0_height_0_subtile_0__pin_I_8_
port 20 nsew signal input
rlabel metal2 s 26146 29200 26202 30000 6 top_width_0_height_0_subtile_0__pin_O_2_
port 21 nsew signal output
rlabel metal4 s 4417 2128 4737 27792 6 vdd
port 22 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vdd
port 22 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vdd
port 22 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vdd
port 22 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vss
port 23 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vss
port 23 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vss
port 23 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vss
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3327318
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/grid_clb/runs/24_02_16_16_06/results/signoff/grid_clb.magic.gds
string GDS_START 183766
<< end >>

