* NGSPICE file created from cby_8__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

.subckt cby_8__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] left_grid_right_width_0_height_0_subtile_0__pin_I_1_
+ left_grid_right_width_0_height_0_subtile_0__pin_I_5_ left_grid_right_width_0_height_0_subtile_0__pin_I_9_
+ prog_clk right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_ vdd vss
XFILLER_0_13_95 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_062_ _012_ vss vss vdd vdd _040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_74 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_114_ mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net41 sky130_fd_sc_hd__inv_2
Xoutput20 net20 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 vss vss vdd vdd right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
Xoutput31 net31 vss vss vdd vdd chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_13_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_061_ mem_right_ipin_1.DFF_1_.Q vss vss vdd vdd _012_ sky130_fd_sc_hd__clkbuf_1
X_113_ net13 vss vss vdd vdd mux_right_ipin_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_0_19 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput21 net21 vss vss vdd vdd chany_bottom_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 vss vss vdd vdd chany_top_out[2] sky130_fd_sc_hd__buf_2
X_060_ _011_ vss vss vdd vdd _041_ sky130_fd_sc_hd__clkbuf_1
X_112_ net4 vss vss vdd vdd mux_right_ipin_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_9_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput33 net33 vss vss vdd vdd chany_top_out[3] sky130_fd_sc_hd__buf_2
Xoutput22 net22 vss vss vdd vdd chany_bottom_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_111_ mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net40 sky130_fd_sc_hd__inv_2
XFILLER_0_10_88 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xoutput34 net34 vss vss vdd vdd chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vss vss vdd vdd chany_bottom_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_66 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_67 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_4_42 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_110_ net16 vss vss vdd vdd mux_right_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_0_1_98 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput35 net35 vss vss vdd vdd chany_top_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput24 net24 vss vss vdd vdd chany_bottom_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_35 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_32 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_169_ mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out _035_ vss vss vdd vdd mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_13_79 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_46 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_98 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput36 net36 vss vss vdd vdd chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput25 net25 vss vss vdd vdd chany_bottom_out[4] sky130_fd_sc_hd__clkbuf_4
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_099_ mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net42 sky130_fd_sc_hd__inv_2
X_168_ mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out _034_ vss vss vdd vdd mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
Xoutput37 net37 vss vss vdd vdd chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vss vss vdd vdd chany_bottom_out[5] sky130_fd_sc_hd__clkbuf_4
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_56 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_11_91 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_098_ _008_ vss vss vdd vdd _016_ sky130_fd_sc_hd__clkbuf_1
X_167_ mux_left_ipin_0.INVTX1_1_.out _033_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput38 net38 vss vss vdd vdd chany_top_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 vss vss vdd vdd chany_bottom_out[6] sky130_fd_sc_hd__clkbuf_4
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_097_ mem_left_ipin_0.DFF_1_.Q vss vss vdd vdd _008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_25 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_36 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_166_ mux_right_ipin_0.INVTX1_3_.out _032_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xoutput39 net39 vss vss vdd vdd left_grid_right_width_0_height_0_subtile_0__pin_I_1_
+ sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 vss vss vdd vdd chany_bottom_out[7] sky130_fd_sc_hd__clkbuf_4
X_149_ net2 vss vss vdd vdd net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_38 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_46 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_14 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_60 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_165_ mux_right_ipin_0.INVTX1_5_.out _031_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_096_ _007_ vss vss vdd vdd _017_ sky130_fd_sc_hd__clkbuf_1
X_148_ net3 vss vss vdd vdd net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_48 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xoutput29 net29 vss vss vdd vdd chany_bottom_out[8] sky130_fd_sc_hd__clkbuf_4
X_079_ mem_right_ipin_0.DFF_1_.Q vss vss vdd vdd _002_ sky130_fd_sc_hd__clkbuf_1
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_181_ mux_right_ipin_2.INVTX1_0_.out _047_ vss vss vdd vdd mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_095_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _007_ sky130_fd_sc_hd__clkbuf_1
X_164_ mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out _030_ vss vss vdd vdd mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_078_ _001_ vss vss vdd vdd _031_ sky130_fd_sc_hd__clkbuf_1
X_147_ net4 vss vss vdd vdd net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_26 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_180_ mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out _046_ vss vss vdd vdd mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_4_49 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_094_ _006_ vss vss vdd vdd _020_ sky130_fd_sc_hd__clkbuf_1
X_163_ net44 _029_ vss vss vdd vdd mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_5_92 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_077_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_71 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_146_ net5 vss vss vdd vdd net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_093_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _006_ sky130_fd_sc_hd__clkbuf_1
X_162_ mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out _028_ vss vss vdd vdd mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_3_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput1 ccff_head vss vss vdd vdd net1 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
X_076_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _037_ sky130_fd_sc_hd__inv_2
X_145_ net6 vss vss vdd vdd net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_059_ mem_right_ipin_1.DFF_0_.Q vss vss vdd vdd _011_ sky130_fd_sc_hd__clkbuf_1
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_092_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _024_ sky130_fd_sc_hd__inv_2
X_161_ mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out _027_ vss vss vdd vdd mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput2 chany_bottom_in[0] vss vss vdd vdd net2 sky130_fd_sc_hd__buf_1
X_127_ clknet_1_0__leaf_prog_clk net49 vss vss vdd vdd mem_right_ipin_2.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_075_ mem_right_ipin_0.DFF_1_.Q vss vss vdd vdd _035_ sky130_fd_sc_hd__inv_2
X_144_ net7 vss vss vdd vdd net35 sky130_fd_sc_hd__clkbuf_1
X_058_ mem_right_ipin_1.DFF_0_.Q vss vss vdd vdd _043_ sky130_fd_sc_hd__inv_2
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_87 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_160_ mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out _026_ vss vss vdd vdd mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_091_ mem_left_ipin_0.DFF_1_.Q vss vss vdd vdd _026_ sky130_fd_sc_hd__inv_2
X_074_ _000_ vss vss vdd vdd _028_ sky130_fd_sc_hd__clkbuf_1
Xinput3 chany_bottom_in[1] vss vss vdd vdd net3 sky130_fd_sc_hd__buf_1
X_143_ net8 vss vss vdd vdd net36 sky130_fd_sc_hd__clkbuf_1
X_057_ mem_right_ipin_1.DFF_1_.Q vss vss vdd vdd _042_ sky130_fd_sc_hd__inv_2
X_126_ clknet_1_0__leaf_prog_clk net47 vss vss vdd vdd net20 sky130_fd_sc_hd__dfxtp_1
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_109_ net3 vss vss vdd vdd mux_right_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_090_ _005_ vss vss vdd vdd _018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput4 chany_bottom_in[2] vss vss vdd vdd net4 sky130_fd_sc_hd__buf_1
X_056_ _010_ vss vss vdd vdd _044_ sky130_fd_sc_hd__clkbuf_1
X_125_ clknet_1_0__leaf_prog_clk net51 vss vss vdd vdd mem_right_ipin_1.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_142_ net9 vss vss vdd vdd net37 sky130_fd_sc_hd__clkbuf_1
X_073_ mem_right_ipin_0.DFF_2_.Q vss vss vdd vdd _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_97 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_163__44 vss vss vdd vdd net44 _163__44/LO sky130_fd_sc_hd__conb_1
X_108_ net12 vss vss vdd vdd mux_right_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XTAP_50 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ net10 vss vss vdd vdd net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_86 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_072_ _015_ vss vss vdd vdd _032_ sky130_fd_sc_hd__clkbuf_1
Xinput5 chany_bottom_in[3] vss vss vdd vdd net5 sky130_fd_sc_hd__buf_1
X_055_ net20 vss vss vdd vdd _010_ sky130_fd_sc_hd__clkbuf_1
X_124_ clknet_1_0__leaf_prog_clk net48 vss vss vdd vdd mem_right_ipin_1.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_107_ net7 vss vss vdd vdd mux_right_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XTAP_51 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ net11 vss vss vdd vdd net21 sky130_fd_sc_hd__clkbuf_1
X_071_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _015_ sky130_fd_sc_hd__clkbuf_1
Xinput6 chany_bottom_in[4] vss vss vdd vdd net6 sky130_fd_sc_hd__buf_1
X_106_ mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net39 sky130_fd_sc_hd__inv_2
X_054_ _009_ vss vss vdd vdd _045_ sky130_fd_sc_hd__clkbuf_1
X_123_ clknet_1_1__leaf_prog_clk net50 vss vss vdd vdd mem_right_ipin_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_41 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _038_ sky130_fd_sc_hd__inv_2
Xinput7 chany_bottom_in[5] vss vss vdd vdd net7 sky130_fd_sc_hd__buf_1
XTAP_30 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_053_ mem_right_ipin_2.DFF_0_.Q vss vss vdd vdd _009_ sky130_fd_sc_hd__clkbuf_1
X_122_ clknet_1_0__leaf_prog_clk net52 vss vss vdd vdd mem_right_ipin_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
Xinput10 chany_bottom_in[8] vss vss vdd vdd net10 sky130_fd_sc_hd__buf_1
X_105_ net19 vss vss vdd vdd mux_left_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XTAP_42 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_31 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 chany_bottom_in[6] vss vss vdd vdd net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_35 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput11 chany_top_in[0] vss vss vdd vdd net11 sky130_fd_sc_hd__buf_1
X_052_ mem_right_ipin_2.DFF_0_.Q vss vss vdd vdd _047_ sky130_fd_sc_hd__inv_2
X_121_ clknet_1_0__leaf_prog_clk net54 vss vss vdd vdd mem_right_ipin_0.DFF_2_.Q sky130_fd_sc_hd__dfxtp_1
X_104_ net11 vss vss vdd vdd mux_left_ipin_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_43 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput9 chany_bottom_in[7] vss vss vdd vdd net9 sky130_fd_sc_hd__clkbuf_1
XTAP_32 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 chany_top_in[1] vss vss vdd vdd net12 sky130_fd_sc_hd__buf_1
X_120_ clknet_1_1__leaf_prog_clk net1 vss vss vdd vdd mem_left_ipin_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_47 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_68 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_103_ net2 vss vss vdd vdd mux_left_ipin_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
Xhold1 mem_right_ipin_2.DFF_0_.Q vss vss vdd vdd net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_69 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_44 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_59 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_33 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 chany_top_in[2] vss vss vdd vdd net13 sky130_fd_sc_hd__buf_1
XFILLER_0_12_93 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_179_ mux_right_ipin_2.INVTX1_1_.out _045_ vss vss vdd vdd mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_102_ net6 vss vss vdd vdd mux_left_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
Xhold2 mem_right_ipin_1.DFF_0_.Q vss vss vdd vdd net48 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_45 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 chany_top_in[3] vss vss vdd vdd net14 sky130_fd_sc_hd__buf_1
XFILLER_0_12_72 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_178_ net46 _044_ vss vss vdd vdd mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_101_ net15 vss vss vdd vdd mux_left_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_3_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xhold3 mem_right_ipin_1.DFF_1_.Q vss vss vdd vdd net49 sky130_fd_sc_hd__dlygate4sd3_1
X_150__43 vss vss vdd vdd net43 _150__43/LO sky130_fd_sc_hd__conb_1
XFILLER_0_0_71 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_46 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 chany_top_in[4] vss vss vdd vdd net15 sky130_fd_sc_hd__buf_1
X_178__46 vss vss vdd vdd net46 _178__46/LO sky130_fd_sc_hd__conb_1
X_100_ net10 vss vss vdd vdd mux_left_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_177_ mux_right_ipin_1.INVTX1_0_.out _043_ vss vss vdd vdd mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_93 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xhold4 mem_left_ipin_0.DFF_2_.Q vss vss vdd vdd net50 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_47 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_50 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_18 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput16 chany_top_in[5] vss vss vdd vdd net16 sky130_fd_sc_hd__buf_1
X_176_ mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out _042_ vss vss vdd vdd mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_159_ mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out _025_ vss vss vdd vdd mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_9_71 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold5 mem_right_ipin_0.DFF_2_.Q vss vss vdd vdd net51 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_48 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_37 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput17 chany_top_in[6] vss vss vdd vdd net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_175_ mux_right_ipin_1.INVTX1_1_.out _041_ vss vss vdd vdd mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_51 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_158_ mux_left_ipin_0.INVTX1_4_.out _024_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_089_ mem_left_ipin_0.DFF_2_.Q vss vss vdd vdd _005_ sky130_fd_sc_hd__clkbuf_1
Xhold6 mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd net52 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_49 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_63 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput18 chany_top_in[7] vss vss vdd vdd net18 sky130_fd_sc_hd__clkbuf_1
X_174_ net45 _040_ vss vss vdd vdd mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_157_ mux_left_ipin_0.INVTX1_2_.out _023_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_088_ _004_ vss vss vdd vdd _019_ sky130_fd_sc_hd__clkbuf_1
Xhold7 mem_left_ipin_0.DFF_1_.Q vss vss vdd vdd net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_96 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_39 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_28 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 chany_top_in[8] vss vss vdd vdd net19 sky130_fd_sc_hd__buf_1
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_173_ mux_left_ipin_0.INVTX1_0_.out _039_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold8 mem_right_ipin_0.DFF_1_.Q vss vss vdd vdd net54 sky130_fd_sc_hd__dlygate4sd3_1
X_087_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _004_ sky130_fd_sc_hd__clkbuf_1
X_156_ mux_left_ipin_0.INVTX1_0_.out _022_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_9_63 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_139_ net12 vss vss vdd vdd net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_32 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_43 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_0_76 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_29 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out _021_ vss vss vdd vdd mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_086_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _023_ sky130_fd_sc_hd__inv_2
X_172_ mux_right_ipin_0.INVTX1_2_.out _038_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold9 mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_97 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_069_ _014_ vss vss vdd vdd _030_ sky130_fd_sc_hd__clkbuf_1
X_138_ net13 vss vss vdd vdd net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_21 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_171_ mux_right_ipin_0.INVTX1_4_.out _037_ vss vss vdd vdd mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_154_ mux_left_ipin_0.INVTX1_5_.out _020_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_085_ _003_ vss vss vdd vdd _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_068_ mem_right_ipin_0.DFF_1_.Q vss vss vdd vdd _014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_12 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_137_ net14 vss vss vdd vdd net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_89 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_88 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_174__45 vss vss vdd vdd net45 _174__45/LO sky130_fd_sc_hd__conb_1
X_170_ mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out _036_ vss vss vdd vdd mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_45 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_084_ mem_left_ipin_0.DFF_1_.Q vss vss vdd vdd _003_ sky130_fd_sc_hd__clkbuf_1
X_153_ mux_left_ipin_0.INVTX1_3_.out _019_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_136_ net15 vss vss vdd vdd net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_067_ _013_ vss vss vdd vdd _033_ sky130_fd_sc_hd__clkbuf_1
X_119_ clknet_1_1__leaf_prog_clk net55 vss vss vdd vdd mem_left_ipin_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_152_ mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out _018_ vss vss vdd vdd mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_083_ mem_left_ipin_0.DFF_0_.Q vss vss vdd vdd _022_ sky130_fd_sc_hd__inv_2
X_135_ net16 vss vss vdd vdd net26 sky130_fd_sc_hd__clkbuf_1
X_118_ clknet_1_1__leaf_prog_clk net53 vss vss vdd vdd mem_left_ipin_0.DFF_2_.Q sky130_fd_sc_hd__dfxtp_1
X_066_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _013_ sky130_fd_sc_hd__clkbuf_1
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_49 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_134_ net17 vss vss vdd vdd net27 sky130_fd_sc_hd__clkbuf_1
X_082_ mem_left_ipin_0.DFF_1_.Q vss vss vdd vdd _025_ sky130_fd_sc_hd__inv_2
X_151_ mux_left_ipin_0.INVTX1_1_.out _017_ vss vss vdd vdd mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_065_ mem_right_ipin_0.DFF_0_.Q vss vss vdd vdd _039_ sky130_fd_sc_hd__inv_2
X_117_ net20 vss vss vdd vdd _046_ sky130_fd_sc_hd__inv_2
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_150_ net43 _016_ vss vss vdd vdd mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_081_ mem_left_ipin_0.DFF_2_.Q vss vss vdd vdd _027_ sky130_fd_sc_hd__inv_2
X_133_ net18 vss vss vdd vdd net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_94 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_80 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_0_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_064_ mem_right_ipin_0.DFF_1_.Q vss vss vdd vdd _036_ sky130_fd_sc_hd__inv_2
X_116_ net14 vss vss vdd vdd mux_right_ipin_2.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_4_9 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput40 net40 vss vss vdd vdd left_grid_right_width_0_height_0_subtile_0__pin_I_5_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_3_38 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_132_ net19 vss vss vdd vdd net29 sky130_fd_sc_hd__clkbuf_1
X_080_ _002_ vss vss vdd vdd _029_ sky130_fd_sc_hd__clkbuf_1
X_063_ mem_right_ipin_0.DFF_2_.Q vss vss vdd vdd _034_ sky130_fd_sc_hd__inv_2
X_115_ net5 vss vss vdd vdd mux_right_ipin_2.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_1_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput41 net41 vss vss vdd vdd left_grid_right_width_0_height_0_subtile_0__pin_I_9_
+ sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 vss vss vdd vdd chany_top_out[0] sky130_fd_sc_hd__buf_2
.ends

