magic
tech sky130A
magscale 1 2
timestamp 1708041461
<< obsli1 >>
rect 1104 2159 14812 17425
<< obsm1 >>
rect 382 1232 15074 17456
<< metal2 >>
rect 570 0 626 800
rect 1306 0 1362 800
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
<< obsm2 >>
rect 388 856 15070 18601
rect 388 711 514 856
rect 682 711 1250 856
rect 1418 711 1986 856
rect 2154 711 2722 856
rect 2890 711 3458 856
rect 3626 711 4194 856
rect 4362 711 4930 856
rect 5098 711 5666 856
rect 5834 711 6402 856
rect 6570 711 7138 856
rect 7306 711 7874 856
rect 8042 711 8610 856
rect 8778 711 9346 856
rect 9514 711 10082 856
rect 10250 711 10818 856
rect 10986 711 11554 856
rect 11722 711 12290 856
rect 12458 711 13026 856
rect 13194 711 13762 856
rect 13930 711 14498 856
rect 14666 711 15070 856
<< metal3 >>
rect 0 18504 800 18624
rect 15200 18504 16000 18624
rect 0 17688 800 17808
rect 15200 17688 16000 17808
rect 0 16872 800 16992
rect 15200 16872 16000 16992
rect 0 16056 800 16176
rect 15200 16056 16000 16176
rect 0 15240 800 15360
rect 15200 15240 16000 15360
rect 0 14424 800 14544
rect 15200 14424 16000 14544
rect 0 13608 800 13728
rect 15200 13608 16000 13728
rect 0 12792 800 12912
rect 15200 12792 16000 12912
rect 0 11976 800 12096
rect 15200 11976 16000 12096
rect 0 11160 800 11280
rect 15200 11160 16000 11280
rect 0 10344 800 10464
rect 15200 10344 16000 10464
rect 0 9528 800 9648
rect 15200 9528 16000 9648
rect 0 8712 800 8832
rect 15200 8712 16000 8832
rect 0 7896 800 8016
rect 15200 7896 16000 8016
rect 0 7080 800 7200
rect 15200 7080 16000 7200
rect 0 6264 800 6384
rect 15200 6264 16000 6384
rect 0 5448 800 5568
rect 15200 5448 16000 5568
rect 0 4632 800 4752
rect 15200 4632 16000 4752
rect 0 3816 800 3936
rect 15200 3816 16000 3936
rect 0 3000 800 3120
rect 15200 3000 16000 3120
rect 0 2184 800 2304
rect 15200 2184 16000 2304
rect 15200 1368 16000 1488
<< obsm3 >>
rect 880 18424 15120 18597
rect 565 17888 15210 18424
rect 880 17608 15120 17888
rect 565 17072 15210 17608
rect 880 16792 15120 17072
rect 565 16256 15210 16792
rect 880 15976 15120 16256
rect 565 15440 15210 15976
rect 880 15160 15120 15440
rect 565 14624 15210 15160
rect 880 14344 15120 14624
rect 565 13808 15210 14344
rect 880 13528 15120 13808
rect 565 12992 15210 13528
rect 880 12712 15120 12992
rect 565 12176 15210 12712
rect 880 11896 15120 12176
rect 565 11360 15210 11896
rect 880 11080 15120 11360
rect 565 10544 15210 11080
rect 880 10264 15120 10544
rect 565 9728 15210 10264
rect 880 9448 15120 9728
rect 565 8912 15210 9448
rect 880 8632 15120 8912
rect 565 8096 15210 8632
rect 880 7816 15120 8096
rect 565 7280 15210 7816
rect 880 7000 15120 7280
rect 565 6464 15210 7000
rect 880 6184 15120 6464
rect 565 5648 15210 6184
rect 880 5368 15120 5648
rect 565 4832 15210 5368
rect 880 4552 15120 4832
rect 565 4016 15210 4552
rect 880 3736 15120 4016
rect 565 3200 15210 3736
rect 880 2920 15120 3200
rect 565 2384 15210 2920
rect 880 2104 15120 2384
rect 565 1568 15210 2104
rect 565 1288 15120 1568
rect 565 715 15210 1288
<< metal4 >>
rect 2657 2128 2977 17456
rect 4370 2128 4690 17456
rect 6084 2128 6404 17456
rect 7797 2128 8117 17456
rect 9511 2128 9831 17456
rect 11224 2128 11544 17456
rect 12938 2128 13258 17456
rect 14651 2128 14971 17456
<< obsm4 >>
rect 795 2048 2577 14517
rect 3057 2048 4290 14517
rect 4770 2048 6004 14517
rect 6484 2048 7717 14517
rect 8197 2048 9431 14517
rect 9911 2048 11144 14517
rect 11624 2048 12821 14517
rect 795 715 12821 2048
<< labels >>
rlabel metal2 s 7930 0 7986 800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 1 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 2 nsew signal input
rlabel metal3 s 15200 17688 16000 17808 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 15200 18504 16000 18624 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 chanx_left_in[0]
port 5 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[1]
port 6 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 chanx_left_in[2]
port 7 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 chanx_left_in[3]
port 8 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[4]
port 9 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[5]
port 10 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 chanx_left_in[6]
port 11 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[7]
port 12 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 chanx_left_in[8]
port 13 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_out[0]
port 14 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 chanx_left_out[1]
port 15 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[2]
port 16 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[3]
port 17 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 chanx_left_out[4]
port 18 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 19 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[6]
port 20 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 chanx_left_out[7]
port 21 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 chanx_left_out[8]
port 22 nsew signal output
rlabel metal3 s 15200 1368 16000 1488 6 chanx_right_in[0]
port 23 nsew signal input
rlabel metal3 s 15200 2184 16000 2304 6 chanx_right_in[1]
port 24 nsew signal input
rlabel metal3 s 15200 3000 16000 3120 6 chanx_right_in[2]
port 25 nsew signal input
rlabel metal3 s 15200 3816 16000 3936 6 chanx_right_in[3]
port 26 nsew signal input
rlabel metal3 s 15200 4632 16000 4752 6 chanx_right_in[4]
port 27 nsew signal input
rlabel metal3 s 15200 5448 16000 5568 6 chanx_right_in[5]
port 28 nsew signal input
rlabel metal3 s 15200 6264 16000 6384 6 chanx_right_in[6]
port 29 nsew signal input
rlabel metal3 s 15200 7080 16000 7200 6 chanx_right_in[7]
port 30 nsew signal input
rlabel metal3 s 15200 7896 16000 8016 6 chanx_right_in[8]
port 31 nsew signal input
rlabel metal3 s 15200 8712 16000 8832 6 chanx_right_out[0]
port 32 nsew signal output
rlabel metal3 s 15200 9528 16000 9648 6 chanx_right_out[1]
port 33 nsew signal output
rlabel metal3 s 15200 10344 16000 10464 6 chanx_right_out[2]
port 34 nsew signal output
rlabel metal3 s 15200 11160 16000 11280 6 chanx_right_out[3]
port 35 nsew signal output
rlabel metal3 s 15200 11976 16000 12096 6 chanx_right_out[4]
port 36 nsew signal output
rlabel metal3 s 15200 12792 16000 12912 6 chanx_right_out[5]
port 37 nsew signal output
rlabel metal3 s 15200 13608 16000 13728 6 chanx_right_out[6]
port 38 nsew signal output
rlabel metal3 s 15200 14424 16000 14544 6 chanx_right_out[7]
port 39 nsew signal output
rlabel metal3 s 15200 15240 16000 15360 6 chanx_right_out[8]
port 40 nsew signal output
rlabel metal2 s 570 0 626 800 6 chany_bottom_in[0]
port 41 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 chany_bottom_in[1]
port 42 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 chany_bottom_in[2]
port 43 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_in[3]
port 44 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_in[4]
port 45 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[5]
port 46 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[6]
port 47 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[7]
port 48 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[8]
port 49 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_out[0]
port 50 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_out[1]
port 51 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_out[2]
port 52 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_out[3]
port 53 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_out[4]
port 54 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_out[5]
port 55 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[6]
port 56 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[7]
port 57 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[8]
port 58 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 59 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 60 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 prog_clk
port 61 nsew signal input
rlabel metal3 s 15200 16056 16000 16176 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 62 nsew signal input
rlabel metal3 s 15200 16872 16000 16992 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 63 nsew signal input
rlabel metal4 s 2657 2128 2977 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 17456 6 vss
port 65 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1121050
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_1__10_/runs/24_02_15_17_56/results/signoff/sb_1__10_.magic.gds
string GDS_START 113884
<< end >>

