* NGSPICE file created from grid_clb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_1 abstract view
.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt grid_clb bottom_width_0_height_0_subtile_0__pin_I_2_ bottom_width_0_height_0_subtile_0__pin_I_6_
+ bottom_width_0_height_0_subtile_0__pin_O_0_ bottom_width_0_height_0_subtile_0__pin_clk_0_
+ ccff_head ccff_tail clk left_width_0_height_0_subtile_0__pin_I_3_ left_width_0_height_0_subtile_0__pin_I_7_
+ left_width_0_height_0_subtile_0__pin_O_1_ prog_clk reset right_width_0_height_0_subtile_0__pin_I_1_
+ right_width_0_height_0_subtile_0__pin_I_5_ right_width_0_height_0_subtile_0__pin_I_9_
+ right_width_0_height_0_subtile_0__pin_O_3_ set top_width_0_height_0_subtile_0__pin_I_0_
+ top_width_0_height_0_subtile_0__pin_I_4_ top_width_0_height_0_subtile_0__pin_I_8_
+ top_width_0_height_0_subtile_0__pin_O_2_ vdd vss
X_2106_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out _0352_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2037_ clknet_4_0_0_prog_clk net90 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_177 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1270_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0082_
+ sky130_fd_sc_hd__clkbuf_1
X_1606_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0377_
+ sky130_fd_sc_hd__inv_2
X_0985_ _0293_ vss vss vdd vdd _0702_ sky130_fd_sc_hd__clkbuf_1
X_2655_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ _0901_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_1537_ _0177_ vss vss vdd vdd _0361_ sky130_fd_sc_hd__clkbuf_1
X_2586_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ _0832_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_1399_ _0127_ vss vss vdd vdd _0507_ sky130_fd_sc_hd__clkbuf_1
X_1468_ _0151_ vss vss vdd vdd _0534_ sky130_fd_sc_hd__clkbuf_1
X_2440_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out _0686_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1322_ _0099_ vss vss vdd vdd _0847_ sky130_fd_sc_hd__inv_2
X_1253_ _0075_ vss vss vdd vdd _0871_ sky130_fd_sc_hd__clkbuf_1
X_2371_ net57 _0617_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1184_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd _0052_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_169 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0968_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0687_
+ sky130_fd_sc_hd__inv_2
X_2569_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ _0815_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_2638_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ _0884_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_37_169 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_45_49 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1871_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ sky130_fd_sc_hd__inv_2
X_1940_ clknet_4_15_0_prog_clk net175 vss vss vdd vdd net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2423_ net27 _0669_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1305_ _0093_ vss vss vdd vdd _0676_ sky130_fd_sc_hd__buf_1
X_2354_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out _0600_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1236_ _0070_ vss vss vdd vdd _0610_ sky130_fd_sc_hd__clkbuf_1
X_2285_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out _0531_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_35_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1167_ _0046_ vss vss vdd vdd _0588_ sky130_fd_sc_hd__clkbuf_1
X_1098_ _0012_ vss vss vdd vdd _0735_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1021_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0306_
+ sky130_fd_sc_hd__clkbuf_1
X_1854_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ sky130_fd_sc_hd__inv_2
X_1923_ clknet_4_10_0_prog_clk net107 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1785_ _0263_ vss vss vdd vdd _0664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_51 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2406_ net35 _0652_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2199_ net26 _0445_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1219_ _0063_ vss vss vdd vdd _0599_ sky130_fd_sc_hd__inv_2
X_2337_ net28 _0583_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2268_ net24 _0514_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold63 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd net97 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold41 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ vss vss vdd vdd net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd net152
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd net163
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_337 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0189_ sky130_fd_sc_hd__clkbuf_1
XTAP_315 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_186 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2122_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out _0368_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
X_2053_ clknet_4_2_0_prog_clk net75 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ sky130_fd_sc_hd__dfxtp_1
X_2511__62 vss vss vdd vdd net62 _2511__62/LO sky130_fd_sc_hd__conb_1
XFILLER_0_29_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1004_ _0288_ vss vss vdd vdd _0677_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_234 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1906_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ sky130_fd_sc_hd__inv_2
X_1837_ net9 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out
+ sky130_fd_sc_hd__inv_2
X_1768_ _0096_ vss vss vdd vdd _0653_ sky130_fd_sc_hd__inv_2
X_1699_ _0235_ vss vss vdd vdd _0442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_197 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_28 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1622_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0814_ sky130_fd_sc_hd__inv_2
X_1553_ _0183_ vss vss vdd vdd _0358_ sky130_fd_sc_hd__clkbuf_1
XTAP_134 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0516_
+ sky130_fd_sc_hd__inv_2
X_2105_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out _0351_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2036_ _0008_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ _0006_ _0007_ vss vss vdd vdd _2036_/Q logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ sky130_fd_sc_hd__dfbbn_1
X_0984_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q vss vss vdd vdd _0293_
+ sky130_fd_sc_hd__clkbuf_1
X_1536_ _0176_ vss vss vdd vdd _0177_ sky130_fd_sc_hd__clkbuf_1
X_2585_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ _0831_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_1605_ _0195_ vss vss vdd vdd _0372_ sky130_fd_sc_hd__inv_2
X_2654_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ _0900_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_14_215 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1398_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q vss vss vdd vdd _0127_
+ sky130_fd_sc_hd__clkbuf_1
X_1467_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q vss vss vdd vdd _0151_
+ sky130_fd_sc_hd__clkbuf_1
X_2019_ clknet_4_4_0_prog_clk net138 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_270 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_229 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_6_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1321_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0099_ sky130_fd_sc_hd__buf_6
X_1252_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0075_ sky130_fd_sc_hd__clkbuf_1
X_2370_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out _0616_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1183_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0573_
+ sky130_fd_sc_hd__inv_2
X_0967_ _0287_ vss vss vdd vdd _0701_ sky130_fd_sc_hd__clkbuf_1
X_1519_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0816_ sky130_fd_sc_hd__inv_2
X_2568_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ _0814_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_2637_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ _0883_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2499_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out _0745_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_37_148 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_36_192 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1870_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_10_20 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2353_ net22 _0599_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2422_ net21 _0668_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1304_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q vss vss vdd vdd _0093_
+ sky130_fd_sc_hd__clkbuf_1
X_1235_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd _0070_
+ sky130_fd_sc_hd__clkbuf_1
X_1166_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0046_
+ sky130_fd_sc_hd__clkbuf_1
X_2284_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out _0530_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_35_83 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_19_159 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1097_ _0020_ vss vss vdd vdd _0749_ sky130_fd_sc_hd__clkbuf_1
X_1999_ clknet_4_14_0_prog_clk net193 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_192 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_33_140 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1020_ _0305_ vss vss vdd vdd _0731_ sky130_fd_sc_hd__clkbuf_1
X_1922_ clknet_4_10_0_prog_clk net116 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1853_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ sky130_fd_sc_hd__inv_2
X_1784_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd _0263_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_74 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2336_ net32 _0582_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2405_ net38 _0651_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2198_ net20 _0444_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_27_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1149_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0039_ sky130_fd_sc_hd__clkbuf_1
X_1218_ _0064_ vss vss vdd vdd _0613_ sky130_fd_sc_hd__clkbuf_1
X_2267_ net30 _0513_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold42 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd net153
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd net164
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_38_221 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_338 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_154 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2121_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out _0367_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2052_ clknet_4_2_0_prog_clk net105 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1003_ _0299_ vss vss vdd vdd _0691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_9 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1905_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ sky130_fd_sc_hd__inv_2
X_1836_ net13 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out
+ sky130_fd_sc_hd__inv_2
X_1698_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd _0235_
+ sky130_fd_sc_hd__clkbuf_1
X_1767_ _0257_ vss vss vdd vdd _0667_ sky130_fd_sc_hd__clkbuf_1
X_2319_ net46 _0565_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1621_ _0207_ vss vss vdd vdd _0803_ sky130_fd_sc_hd__clkbuf_1
X_1552_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd _0183_
+ sky130_fd_sc_hd__clkbuf_1
X_2104_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out _0350_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_124 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _0146_ vss vss vdd vdd _0510_ sky130_fd_sc_hd__inv_2
X_2035_ clknet_4_1_0_prog_clk net157 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1819_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0768_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_162 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2175__50 vss vss vdd vdd net50 _2175__50/LO sky130_fd_sc_hd__conb_1
X_0983_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q vss vss vdd vdd _0690_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_205 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1535_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd _0176_
+ sky130_fd_sc_hd__buf_6
X_1604_ _0202_ vss vss vdd vdd _0386_ sky130_fd_sc_hd__clkbuf_1
X_2584_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ _0830_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
X_2653_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ _0899_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1397_ _0126_ vss vss vdd vdd _0508_ sky130_fd_sc_hd__buf_1
X_1466_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q vss vss vdd vdd _0522_
+ sky130_fd_sc_hd__inv_2
X_2018_ clknet_4_4_0_prog_clk net84 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_208 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1320_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0851_ sky130_fd_sc_hd__inv_2
X_1251_ _0063_ vss vss vdd vdd _0593_ sky130_fd_sc_hd__inv_2
X_1182_ _0044_ vss vss vdd vdd _0568_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2636_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ _0882_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_0966_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0287_
+ sky130_fd_sc_hd__clkbuf_1
X_1518_ _0169_ vss vss vdd vdd _0804_ sky130_fd_sc_hd__clkbuf_1
X_2567_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ _0813_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_2498_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out _0744_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1449_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0145_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_19 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1303_ _0033_ vss vss vdd vdd _0874_ sky130_fd_sc_hd__inv_2
X_2352_ net24 _0598_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2421_ net29 _0667_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2283_ net26 _0529_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1234_ _0069_ vss vss vdd vdd _0615_ sky130_fd_sc_hd__clkbuf_1
X_1165_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q vss vss vdd vdd _0577_
+ sky130_fd_sc_hd__inv_2
X_1096_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd _0020_
+ sky130_fd_sc_hd__clkbuf_1
X_1998_ clknet_4_15_0_prog_clk net153 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2619_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ _0865_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_0949_ _0277_ vss vss vdd vdd _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_171 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_1852_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ sky130_fd_sc_hd__inv_2
X_1921_ clknet_4_10_0_prog_clk net100 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1783_ _0262_ vss vss vdd vdd _0670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_42 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2404_ net43 _0650_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2335_ net36 _0581_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2266_ net34 _0512_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2197_ net28 _0443_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1148_ _0038_ vss vss vdd vdd _0864_ sky130_fd_sc_hd__clkbuf_1
X_1217_ _0063_ vss vss vdd vdd _0064_ sky130_fd_sc_hd__clkbuf_1
X_1079_ _0014_ vss vss vdd vdd _0756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_144 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xhold65 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd net165
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q vss vss vdd vdd net154
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q vss vss vdd vdd net77
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd net110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_233 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_328 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out _0366_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2051_ clknet_4_2_0_prog_clk net131 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1002_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd _0299_
+ sky130_fd_sc_hd__clkbuf_1
X_1835_ net5 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_32_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_29_233 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1904_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ sky130_fd_sc_hd__inv_2
X_1697_ _0234_ vss vss vdd vdd _0447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_122 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_188 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1766_ _0096_ vss vss vdd vdd _0257_ sky130_fd_sc_hd__clkbuf_1
X_2249_ net44 _0495_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2318_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out _0564_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_258 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_26_225 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1620_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0207_ sky130_fd_sc_hd__clkbuf_1
X_1551_ _0182_ vss vss vdd vdd _0363_ sky130_fd_sc_hd__clkbuf_1
XTAP_114 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1482_ _0156_ vss vss vdd vdd _0524_ sky130_fd_sc_hd__clkbuf_1
X_2103_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out _0349_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_125 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ clknet_4_1_0_prog_clk net110 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1818_ _0028_ vss vss vdd vdd _0762_ sky130_fd_sc_hd__inv_2
X_1749_ _0162_ vss vss vdd vdd _0538_ sky130_fd_sc_hd__inv_2
X_2652_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ _0898_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
X_0982_ _0288_ vss vss vdd vdd _0681_ sky130_fd_sc_hd__inv_2
X_1534_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0351_
+ sky130_fd_sc_hd__inv_2
X_1603_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd _0202_
+ sky130_fd_sc_hd__clkbuf_1
X_2583_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ _0829_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1465_ _0146_ vss vss vdd vdd _0513_ sky130_fd_sc_hd__inv_2
X_1396_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q vss vss vdd vdd _0126_
+ sky130_fd_sc_hd__clkbuf_1
X_2017_ _0005_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ _0003_ _0004_ vss vss vdd vdd _2017_/Q logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ sky130_fd_sc_hd__dfbbn_1
Xhold140 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd net207
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1181_ _0051_ vss vss vdd vdd _0582_ sky130_fd_sc_hd__clkbuf_1
X_1250_ _0074_ vss vss vdd vdd _0607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_40_63 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2635_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ _0881_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_0965_ _0286_ vss vss vdd vdd _0703_ sky130_fd_sc_hd__clkbuf_1
X_1517_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0169_ sky130_fd_sc_hd__clkbuf_1
X_2566_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ _0812_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_1448_ _0144_ vss vss vdd vdd _0535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_63 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_275 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2497_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out _0743_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1379_ _0110_ vss vss vdd vdd _0454_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_128 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_28_117 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2420_ net33 _0666_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1302_ _0092_ vss vss vdd vdd _0867_ sky130_fd_sc_hd__clkbuf_1
X_1233_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0069_
+ sky130_fd_sc_hd__clkbuf_1
X_2351_ net30 _0597_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2282_ net20 _0528_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_86 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_35_41 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1164_ _0044_ vss vss vdd vdd _0571_ sky130_fd_sc_hd__inv_2
X_1095_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0741_
+ sky130_fd_sc_hd__inv_2
X_1997_ clknet_4_14_0_prog_clk net94 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_0948_ _0277_ vss vss vdd vdd _0330_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_139 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_2549_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ _0795_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_42_175 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2618_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ _0864_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_18_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1851_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_24_120 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1920_ clknet_4_10_0_prog_clk net99 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_197 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1782_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0262_
+ sky130_fd_sc_hd__clkbuf_1
X_2403_ net46 _0649_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_73 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_46_40 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2196_ net32 _0442_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1216_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd _0063_
+ sky130_fd_sc_hd__buf_6
X_2334_ net40 _0580_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2265_ net38 _0511_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1147_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0038_ sky130_fd_sc_hd__clkbuf_1
X_1078_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0014_
+ sky130_fd_sc_hd__clkbuf_1
Xhold11 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ vss vss vdd vdd net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q vss vss vdd vdd net155
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd net166
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_329 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ clknet_4_2_0_prog_clk net118 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1001_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0684_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_16_43 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_76 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_16_98 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_44_259 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2578__65 vss vss vdd vdd net65 _2578__65/LO sky130_fd_sc_hd__conb_1
X_1834_ net1 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out
+ sky130_fd_sc_hd__inv_2
X_1903_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ sky130_fd_sc_hd__inv_2
X_1765_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0658_
+ sky130_fd_sc_hd__inv_2
X_1696_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0234_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_134 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_156 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2179_ net46 _0425_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2248_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out _0494_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_2317_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out _0563_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_26_248 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1550_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0182_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_126 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd _0156_
+ sky130_fd_sc_hd__clkbuf_1
X_2102_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out _0348_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_27_42 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_159 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ clknet_4_1_0_prog_clk net112 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_204 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_40_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1817_ _0273_ vss vss vdd vdd _0776_ sky130_fd_sc_hd__clkbuf_1
X_1748_ _0251_ vss vss vdd vdd _0552_ sky130_fd_sc_hd__clkbuf_1
X_1679_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd _0228_
+ sky130_fd_sc_hd__buf_6
XFILLER_0_7_74 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_0981_ _0292_ vss vss vdd vdd _0695_ sky130_fd_sc_hd__clkbuf_1
X_1602_ _0201_ vss vss vdd vdd _0391_ sky130_fd_sc_hd__clkbuf_1
X_2582_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ _0828_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_2651_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ _0897_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
X_1533_ _0175_ vss vss vdd vdd _0365_ sky130_fd_sc_hd__clkbuf_1
X_1395_ _0125_ vss vss vdd vdd _0827_ sky130_fd_sc_hd__clkbuf_1
X_1464_ _0150_ vss vss vdd vdd _0527_ sky130_fd_sc_hd__clkbuf_1
X_2016_ clknet_4_6_0_prog_clk net133 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold130 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd net197
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_284 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_21 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1180_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd _0051_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_181 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_237 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0964_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q vss vss vdd vdd _0286_
+ sky130_fd_sc_hd__clkbuf_1
X_2565_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ _0811_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
X_1516_ _0168_ vss vss vdd vdd _0797_ sky130_fd_sc_hd__clkbuf_1
X_2634_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ _0880_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_1378_ _0120_ vss vss vdd vdd _0468_ sky130_fd_sc_hd__clkbuf_1
X_1447_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q vss vss vdd vdd _0144_
+ sky130_fd_sc_hd__clkbuf_1
X_2496_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out _0742_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_151 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1301_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0092_ sky130_fd_sc_hd__clkbuf_1
X_2350_ net34 _0596_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1232_ _0068_ vss vss vdd vdd _0618_ sky130_fd_sc_hd__clkbuf_1
X_2281_ net28 _0527_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1163_ _0045_ vss vss vdd vdd _0585_ sky130_fd_sc_hd__clkbuf_1
X_1094_ _0012_ vss vss vdd vdd _0736_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_184 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_0947_ _0279_ vss vss vdd vdd _0904_ sky130_fd_sc_hd__clkbuf_1
X_1996_ clknet_4_11_0_prog_clk net184 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2548_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ _0794_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_2617_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ _0863_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_5_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_2479_ net27 _0725_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_18_184 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1850_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ sky130_fd_sc_hd__inv_2
X_1781_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q vss vss vdd vdd _0660_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_21_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2402_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out _0648_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_2333_ net44 _0579_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_96 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2195_ net36 _0441_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1146_ _0033_ vss vss vdd vdd _0879_ sky130_fd_sc_hd__inv_2
X_1215_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0603_
+ sky130_fd_sc_hd__inv_2
X_2264_ net42 _0510_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2427__59 vss vss vdd vdd net59 _2427__59/LO sky130_fd_sc_hd__conb_1
X_1077_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q vss vss vdd vdd _0745_
+ sky130_fd_sc_hd__inv_2
X_1979_ clknet_4_9_0_prog_clk net198 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
Xhold56 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd net156
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd net134 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_319 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _0288_ vss vss vdd vdd _0678_ sky130_fd_sc_hd__inv_2
X_1902_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ sky130_fd_sc_hd__inv_2
X_1764_ _0096_ vss vss vdd vdd _0654_ sky130_fd_sc_hd__inv_2
X_1833_ net8 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out
+ sky130_fd_sc_hd__inv_2
X_1695_ _0233_ vss vss vdd vdd _0450_ sky130_fd_sc_hd__clkbuf_1
X_2316_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out _0562_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2178_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out _0424_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_2247_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out _0493_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1129_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0032_ sky130_fd_sc_hd__clkbuf_1
XTAP_127 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _0155_ vss vss vdd vdd _0530_ sky130_fd_sc_hd__clkbuf_1
X_2101_ net23 _0347_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2032_ clknet_4_1_0_prog_clk net113 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1678_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0435_
+ sky130_fd_sc_hd__inv_2
X_1816_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd _0273_
+ sky130_fd_sc_hd__clkbuf_1
X_1747_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd _0251_
+ sky130_fd_sc_hd__clkbuf_1
X_0980_ _0288_ vss vss vdd vdd _0292_ sky130_fd_sc_hd__clkbuf_1
X_1532_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0175_
+ sky130_fd_sc_hd__clkbuf_1
X_1601_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0201_
+ sky130_fd_sc_hd__clkbuf_1
X_2581_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ _0827_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2650_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ _0896_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_1394_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0125_ sky130_fd_sc_hd__clkbuf_1
X_1463_ _0146_ vss vss vdd vdd _0150_ sky130_fd_sc_hd__clkbuf_1
X_2015_ clknet_4_7_0_prog_clk net70 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold120 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd net187
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd net198
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_193 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_40_43 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0963_ _0285_ vss vss vdd vdd _0704_ sky130_fd_sc_hd__clkbuf_1
X_2564_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ _0810_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
X_1515_ _0165_ vss vss vdd vdd _0168_ sky130_fd_sc_hd__clkbuf_1
X_2633_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ _0879_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
X_2495_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out _0741_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1377_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd _0120_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_32 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1446_ _0143_ vss vss vdd vdd _0536_ sky130_fd_sc_hd__buf_1
XFILLER_0_36_163 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_36_152 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_35_32 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1300_ _0080_ vss vss vdd vdd _0621_ sky130_fd_sc_hd__inv_2
X_1231_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q vss vss vdd vdd _0068_
+ sky130_fd_sc_hd__clkbuf_1
X_1162_ _0044_ vss vss vdd vdd _0045_ sky130_fd_sc_hd__clkbuf_1
X_2280_ net32 _0526_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_77 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_108 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1093_ _0019_ vss vss vdd vdd _0750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_152 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2616_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ _0862_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_0946_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0279_ sky130_fd_sc_hd__clkbuf_1
X_1995_ clknet_4_11_0_prog_clk net188 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2547_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ _0793_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_1429_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q vss vss vdd vdd _0492_
+ sky130_fd_sc_hd__inv_2
X_2478_ net21 _0724_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1780_ _0096_ vss vss vdd vdd _0651_ sky130_fd_sc_hd__inv_2
X_2401_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out _0647_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2332_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out _0578_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
X_2194_ net40 _0440_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1145_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0884_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1214_ _0062_ vss vss vdd vdd _0617_ sky130_fd_sc_hd__clkbuf_1
X_2263_ net46 _0509_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1076_ _0012_ vss vss vdd vdd _0739_ sky130_fd_sc_hd__inv_2
X_1978_ clknet_4_9_0_prog_clk net173 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_15_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0929_ _0009_ net11 vss vss vdd vdd _0010_ sky130_fd_sc_hd__nand2_1
Xhold13 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q vss vss vdd vdd net146
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd net91 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_309 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_1832_ net12 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out
+ sky130_fd_sc_hd__inv_2
X_1901_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ sky130_fd_sc_hd__inv_2
X_1694_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q vss vss vdd vdd _0233_
+ sky130_fd_sc_hd__clkbuf_1
X_1763_ _0256_ vss vss vdd vdd _0858_ sky130_fd_sc_hd__buf_1
X_2246_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out _0492_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2315_ net55 _0561_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2177_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out _0423_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1059_ _0307_ vss vss vdd vdd _0705_ sky130_fd_sc_hd__inv_2
X_1128_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ vss vss vdd vdd _0856_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_294 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2100_ net24 _0346_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_128 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_43 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2031_ clknet_4_4_0_prog_clk net82 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ sky130_fd_sc_hd__dfxtp_1
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1815_ _0272_ vss vss vdd vdd _0782_ sky130_fd_sc_hd__clkbuf_1
X_1677_ _0227_ vss vss vdd vdd _0449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_242 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1746_ _0250_ vss vss vdd vdd _0558_ sky130_fd_sc_hd__clkbuf_1
X_2229_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out _0475_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_261 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_31_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1531_ _0174_ vss vss vdd vdd _0367_ sky130_fd_sc_hd__clkbuf_1
X_1600_ _0200_ vss vss vdd vdd _0394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_169 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1462_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0518_
+ sky130_fd_sc_hd__inv_2
X_2580_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ _0826_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_22_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1393_ _0099_ vss vss vdd vdd _0842_ sky130_fd_sc_hd__inv_2
X_2014_ clknet_4_7_0_prog_clk net101 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ sky130_fd_sc_hd__dfxtp_1
Xhold110 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q vss vss vdd vdd net177
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _0162_ vss vss vdd vdd _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold121 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd net188
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_280 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2632_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ _0878_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
X_0962_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q vss vss vdd vdd _0285_
+ sky130_fd_sc_hd__clkbuf_1
X_2563_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ _0809_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_1514_ _0165_ vss vss vdd vdd _0812_ sky130_fd_sc_hd__inv_2
X_1445_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q vss vss vdd vdd _0143_
+ sky130_fd_sc_hd__clkbuf_1
X_2494_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out _0740_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1376_ _0119_ vss vss vdd vdd _0474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_44 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_45_131 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1230_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q vss vss vdd vdd _0606_
+ sky130_fd_sc_hd__inv_2
X_1161_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd _0044_
+ sky130_fd_sc_hd__buf_6
X_1092_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd _0019_
+ sky130_fd_sc_hd__clkbuf_1
X_1994_ clknet_4_14_0_prog_clk net167 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2615_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ _0861_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_0945_ _0278_ vss vss vdd vdd _0900_ sky130_fd_sc_hd__clkbuf_1
X_2546_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ _0792_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1428_ _0129_ vss vss vdd vdd _0483_ sky130_fd_sc_hd__inv_2
X_2477_ net28 _0723_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1359_ _0110_ vss vss vdd vdd _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_131 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_33_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2400_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out _0646_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_21 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_2262_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out _0508_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_2331_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out _0577_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1213_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0062_
+ sky130_fd_sc_hd__clkbuf_1
X_2193_ net44 _0439_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1144_ _0037_ vss vss vdd vdd _0872_ sky130_fd_sc_hd__clkbuf_1
X_1075_ _0013_ vss vss vdd vdd _0753_ sky130_fd_sc_hd__clkbuf_1
X_1977_ clknet_4_9_0_prog_clk net155 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2529_ net45 _0775_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_0928_ net7 vss vss vdd vdd _0009_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_15_156 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold25 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_281 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1831_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ sky130_fd_sc_hd__inv_2
X_1900_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__inv_2
X_1693_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q vss vss vdd vdd _0438_
+ sky130_fd_sc_hd__inv_2
X_1762_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ vss vss vdd vdd _0256_ sky130_fd_sc_hd__clkbuf_1
X_2245_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out _0491_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2176_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out _0422_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2314_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out _0560_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1127_ _0031_ vss vss vdd vdd _0780_ sky130_fd_sc_hd__clkbuf_1
X_1058_ _0318_ vss vss vdd vdd _0719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_207 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput15 net15 vss vss vdd vdd bottom_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_262 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_2030_ clknet_4_4_0_prog_clk net83 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ sky130_fd_sc_hd__dfxtp_1
XTAP_129 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_77 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_43_33 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1814_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0272_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_284 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_251 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1745_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0250_
+ sky130_fd_sc_hd__clkbuf_1
X_1676_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0227_
+ sky130_fd_sc_hd__clkbuf_1
X_2228_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out _0474_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_30_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2159_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out _0405_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1530_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q vss vss vdd vdd _0174_
+ sky130_fd_sc_hd__clkbuf_1
X_1392_ _0124_ vss vss vdd vdd _0834_ sky130_fd_sc_hd__clkbuf_1
X_1461_ _0146_ vss vss vdd vdd _0514_ sky130_fd_sc_hd__inv_2
X_2013_ clknet_4_7_0_prog_clk net128 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ sky130_fd_sc_hd__dfxtp_1
Xhold133 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd net200
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd net167
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0546_
+ sky130_fd_sc_hd__inv_2
Xhold122 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q vss vss vdd vdd net189
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q vss vss vdd vdd net178
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q vss vss vdd vdd _0408_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_39_151 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0961_ _0284_ vss vss vdd vdd _0897_ sky130_fd_sc_hd__buf_1
X_2562_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ _0808_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_2631_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ _0877_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_1375_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0119_
+ sky130_fd_sc_hd__clkbuf_1
X_1513_ _0167_ vss vss vdd vdd _0802_ sky130_fd_sc_hd__clkbuf_1
X_1444_ _0142_ vss vss vdd vdd _0826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_246 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2493_ net22 _0739_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_290 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1160_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0575_
+ sky130_fd_sc_hd__inv_2
X_1091_ _0018_ vss vss vdd vdd _0755_ sky130_fd_sc_hd__clkbuf_1
X_1993_ clknet_4_14_0_prog_clk net150 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_143 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_0944_ _0277_ vss vss vdd vdd _0278_ sky130_fd_sc_hd__clkbuf_1
X_2545_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ _0791_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_2614_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ _0860_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1358_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0462_
+ sky130_fd_sc_hd__inv_2
X_1427_ _0137_ vss vss vdd vdd _0497_ sky130_fd_sc_hd__clkbuf_1
X_2476_ net33 _0722_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1289_ _0088_ vss vss vdd vdd _0637_ sky130_fd_sc_hd__clkbuf_1
X_2287__54 vss vss vdd vdd net54 _2287__54/LO sky130_fd_sc_hd__conb_1
XFILLER_0_24_102 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_46_44 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_46_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2192_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out _0438_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2261_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out _0507_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1212_ _0061_ vss vss vdd vdd _0619_ sky130_fd_sc_hd__clkbuf_1
X_2330_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out _0576_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1143_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0037_ sky130_fd_sc_hd__clkbuf_1
X_1074_ _0012_ vss vss vdd vdd _0013_ sky130_fd_sc_hd__clkbuf_1
X_1976_ clknet_4_3_0_prog_clk net171 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_102 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_15_135 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2528_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out _0774_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
Xhold37 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd net93 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ net47 _0705_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold15 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd net115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_293 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1830_ _0176_ vss vss vdd vdd _0341_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_238 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1761_ _0255_ vss vss vdd vdd _0668_ sky130_fd_sc_hd__clkbuf_1
X_1692_ _0228_ vss vss vdd vdd _0429_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_4_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_2313_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out _0559_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1126_ _0028_ vss vss vdd vdd _0031_ sky130_fd_sc_hd__clkbuf_1
X_2175_ net50 _0421_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2244_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out _0490_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1057_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd _0318_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_43_263 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1959_ clknet_4_6_0_prog_clk net197 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
Xoutput16 net16 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_0_34_274 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_119 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_68 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1813_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q vss vss vdd vdd _0772_
+ sky130_fd_sc_hd__inv_2
X_1744_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q vss vss vdd vdd _0548_
+ sky130_fd_sc_hd__inv_2
X_1675_ _0226_ vss vss vdd vdd _0451_ sky130_fd_sc_hd__clkbuf_1
X_2227_ net26 _0473_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2158_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out _0404_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2089_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ _0335_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_1109_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_241 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_22_200 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1391_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0124_ sky130_fd_sc_hd__clkbuf_1
X_1460_ _0149_ vss vss vdd vdd _0528_ sky130_fd_sc_hd__clkbuf_1
X_2012_ clknet_4_7_0_prog_clk net126 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_205 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold123 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q vss vss vdd vdd net190
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _0212_ vss vss vdd vdd _0399_ sky130_fd_sc_hd__inv_2
Xhold101 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd net168
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd net179
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_244 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold134 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd net201
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _0162_ vss vss vdd vdd _0542_ sky130_fd_sc_hd__inv_2
X_1589_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0197_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0960_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0284_ sky130_fd_sc_hd__clkbuf_1
X_2561_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ _0807_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_40_68 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1512_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0167_ sky130_fd_sc_hd__clkbuf_1
X_2492_ net25 _0738_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2630_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ _0876_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_1374_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q vss vss vdd vdd _0464_
+ sky130_fd_sc_hd__inv_2
X_2544__64 vss vss vdd vdd net64 _2544__64/LO sky130_fd_sc_hd__conb_1
X_1443_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_80 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XTAP_291 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out vss vss vdd vdd
+ net40 sky130_fd_sc_hd__clkbuf_4
X_1090_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0018_
+ sky130_fd_sc_hd__clkbuf_1
X_0943_ _0277_ vss vss vdd vdd _0331_ sky130_fd_sc_hd__inv_2
X_1992_ clknet_4_8_0_prog_clk net161 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2544_ net64 _0790_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_2613_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ _0859_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_2475_ net37 _0721_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1357_ _0110_ vss vss vdd vdd _0458_ sky130_fd_sc_hd__inv_2
X_1426_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd _0137_
+ sky130_fd_sc_hd__clkbuf_1
X_1288_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd _0088_
+ sky130_fd_sc_hd__clkbuf_1
X_2191_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out _0437_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2260_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out _0506_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1142_ _0036_ vss vss vdd vdd _0865_ sky130_fd_sc_hd__clkbuf_1
X_1211_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q vss vss vdd vdd _0061_
+ sky130_fd_sc_hd__clkbuf_1
X_1073_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd _0012_
+ sky130_fd_sc_hd__buf_6
X_1975_ clknet_4_3_0_prog_clk net202 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_169 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_30_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold27 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ vss vss vdd vdd net94 sky130_fd_sc_hd__dlygate4sd3_1
X_2527_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out _0773_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1409_ _0131_ vss vss vdd vdd _0504_ sky130_fd_sc_hd__clkbuf_1
Xhold16 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd net105 sky130_fd_sc_hd__dlygate4sd3_1
X_2458_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out _0704_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_8
X_2389_ net44 _0635_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold49 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd net116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_272 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1691_ _0232_ vss vss vdd vdd _0443_ sky130_fd_sc_hd__clkbuf_1
X_1760_ _0096_ vss vss vdd vdd _0255_ sky130_fd_sc_hd__clkbuf_1
X_2312_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out _0558_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1125_ _0030_ vss vss vdd vdd _0784_ sky130_fd_sc_hd__clkbuf_1
X_2174_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out _0420_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2243_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out _0489_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1056_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0712_
+ sky130_fd_sc_hd__inv_2
Xoutput17 net17 vss vss vdd vdd left_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1958_ clknet_4_6_0_prog_clk net187 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1889_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ sky130_fd_sc_hd__inv_2
XTAP_109 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_13 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_47 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1674_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q vss vss vdd vdd _0226_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_212 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1812_ _0028_ vss vss vdd vdd _0763_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1743_ _0162_ vss vss vdd vdd _0539_ sky130_fd_sc_hd__inv_2
X_2226_ net20 _0472_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_40_289 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2157_ net23 _0403_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1108_ _0012_ vss vss vdd vdd _0733_ sky130_fd_sc_hd__inv_2
X_2088_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ _0334_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_3 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_17_91 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1039_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q vss vss vdd vdd _0312_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_278 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_31_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_180 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1390_ _0123_ vss vss vdd vdd _0828_ sky130_fd_sc_hd__clkbuf_1
X_2011_ clknet_4_7_0_prog_clk net130 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1588_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q vss vss vdd vdd _0381_
+ sky130_fd_sc_hd__inv_2
X_1657_ _0220_ vss vss vdd vdd _0413_ sky130_fd_sc_hd__clkbuf_1
X_1726_ _0244_ vss vss vdd vdd _0556_ sky130_fd_sc_hd__clkbuf_1
Xhold135 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd net202
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd net191
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q vss vss vdd vdd net180
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd net169
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2209_ net38 _0455_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2483__61 vss vss vdd vdd net61 _2483__61/LO sky130_fd_sc_hd__conb_1
XFILLER_0_39_175 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_2560_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ _0806_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1511_ _0166_ vss vss vdd vdd _0798_ sky130_fd_sc_hd__clkbuf_1
X_2491_ net31 _0737_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1442_ _0099_ vss vss vdd vdd _0841_ sky130_fd_sc_hd__inv_2
X_1373_ _0110_ vss vss vdd vdd _0455_ sky130_fd_sc_hd__inv_2
X_1709_ _0238_ vss vss vdd vdd _0440_ sky130_fd_sc_hd__clkbuf_1
XTAP_292 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out vss vss vdd vdd
+ net30 sky130_fd_sc_hd__clkbuf_4
Xfanout41 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out vss vss vdd vdd
+ net41 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_69 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_156 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0942_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0277_ sky130_fd_sc_hd__buf_6
X_2612_ net66 _0858_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1991_ clknet_4_12_0_prog_clk net195 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2543_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ _0789_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_2474_ net41 _0720_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1425_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0489_
+ sky130_fd_sc_hd__inv_2
X_1356_ _0113_ vss vss vdd vdd _0472_ sky130_fd_sc_hd__clkbuf_1
X_1287_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0629_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_32_170 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_46_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2190_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out _0436_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1141_ _0033_ vss vss vdd vdd _0036_ sky130_fd_sc_hd__clkbuf_1
X_1210_ _0060_ vss vss vdd vdd _0620_ sky130_fd_sc_hd__buf_1
X_1072_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0743_
+ sky130_fd_sc_hd__inv_2
X_1974_ clknet_4_2_0_prog_clk net179 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
Xhold17 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd net84 sky130_fd_sc_hd__dlygate4sd3_1
X_2526_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out _0772_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1408_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0131_
+ sky130_fd_sc_hd__clkbuf_1
Xhold28 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd net95 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out _0634_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_2457_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out _0703_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold39 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd net106 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_46_240 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_14_181 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_107 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1690_ _0228_ vss vss vdd vdd _0232_ sky130_fd_sc_hd__clkbuf_1
X_2242_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out _0488_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2311_ net26 _0557_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1124_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0030_
+ sky130_fd_sc_hd__clkbuf_1
X_2173_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out _0419_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1055_ _0307_ vss vss vdd vdd _0706_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1957_ clknet_4_6_0_prog_clk net140 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_189 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput18 net18 vss vss vdd vdd right_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__clkbuf_4
X_1888_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_11_151 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2509_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out _0755_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1811_ _0271_ vss vss vdd vdd _0777_ sky130_fd_sc_hd__clkbuf_1
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1673_ _0225_ vss vss vdd vdd _0452_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_235 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1742_ _0249_ vss vss vdd vdd _0553_ sky130_fd_sc_hd__clkbuf_1
X_2225_ net28 _0471_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2156_ net25 _0402_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1107_ _0023_ vss vss vdd vdd _0747_ sky130_fd_sc_hd__clkbuf_1
X_2087_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ _0333_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_1038_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q vss vss vdd vdd _0718_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_81 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_7 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_22_246 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2010_ clknet_4_7_0_prog_clk net132 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1725_ _0162_ vss vss vdd vdd _0244_ sky130_fd_sc_hd__clkbuf_1
X_1587_ _0195_ vss vss vdd vdd _0375_ sky130_fd_sc_hd__inv_2
Xhold136 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q vss vss vdd vdd net203
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q vss vss vdd vdd net170
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd net192
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd _0220_
+ sky130_fd_sc_hd__clkbuf_1
Xhold114 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q vss vss vdd vdd net181
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2139_ net37 _0385_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2208_ net42 _0454_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_39_165 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1510_ _0165_ vss vss vdd vdd _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_205 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_227 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2490_ net35 _0736_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1441_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0848_ sky130_fd_sc_hd__inv_2
X_1372_ _0118_ vss vss vdd vdd _0469_ sky130_fd_sc_hd__clkbuf_1
X_1708_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd _0238_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_293 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1639_ _0214_ vss vss vdd vdd _0420_ sky130_fd_sc_hd__clkbuf_1
Xfanout31 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out vss vss vdd vdd
+ net31 sky130_fd_sc_hd__buf_2
Xfanout42 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out vss vss vdd vdd
+ net42 sky130_fd_sc_hd__clkbuf_4
Xfanout20 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net20 sky130_fd_sc_hd__buf_4
XFILLER_0_10_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1990_ clknet_4_12_0_prog_clk net168 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_102 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0941_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0335_ sky130_fd_sc_hd__inv_2
X_2542_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out _0788_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2611_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ _0857_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1355_ _0110_ vss vss vdd vdd _0113_ sky130_fd_sc_hd__clkbuf_1
X_2473_ net45 _0719_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1424_ _0129_ vss vss vdd vdd _0484_ sky130_fd_sc_hd__inv_2
X_1286_ _0080_ vss vss vdd vdd _0624_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_18_179 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_149 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1140_ _0033_ vss vss vdd vdd _0880_ sky130_fd_sc_hd__inv_2
X_1071_ _0323_ vss vss vdd vdd _0757_ sky130_fd_sc_hd__clkbuf_1
X_1973_ clknet_4_2_0_prog_clk net147 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2525_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out _0771_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_23_193 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_39_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1338_ _0099_ vss vss vdd vdd _0844_ sky130_fd_sc_hd__inv_2
X_1407_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q vss vss vdd vdd _0493_
+ sky130_fd_sc_hd__inv_2
X_2387_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out _0633_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
Xhold29 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd net96 sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out _0702_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold18 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd net85 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q vss vss vdd vdd _0633_
+ sky130_fd_sc_hd__inv_2
X_2241_ net22 _0487_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2172_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out _0418_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2310_ net20 _0556_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1123_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q vss vss vdd vdd _0773_
+ sky130_fd_sc_hd__inv_2
X_1054_ _0317_ vss vss vdd vdd _0720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_222 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1956_ clknet_4_5_0_prog_clk net177 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1887_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_7_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_124 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_22_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput19 net19 vss vss vdd vdd top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__clkbuf_4
X_2508_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out _0754_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2439_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out _0685_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1810_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd _0271_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_127 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1741_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd _0249_
+ sky130_fd_sc_hd__clkbuf_1
X_1672_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q vss vss vdd vdd _0225_
+ sky130_fd_sc_hd__clkbuf_1
X_2224_ net32 _0470_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2155_ net30 _0401_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1106_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd _0023_
+ sky130_fd_sc_hd__clkbuf_1
X_2086_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ _0332_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_1037_ _0307_ vss vss vdd vdd _0709_ sky130_fd_sc_hd__inv_2
X_1939_ clknet_4_15_0_prog_clk net194 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_3_0_prog_clk sky130_fd_sc_hd__clkbuf_8
Xhold115 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd net182
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd net193
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q vss vss vdd vdd net171
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ _0243_ vss vss vdd vdd _0560_ sky130_fd_sc_hd__clkbuf_1
X_1586_ _0196_ vss vss vdd vdd _0389_ sky130_fd_sc_hd__clkbuf_1
X_1655_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0405_
+ sky130_fd_sc_hd__inv_2
Xhold137 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_152 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2207_ net46 _0453_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2138_ net40 _0384_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_12_280 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1371_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd _0118_
+ sky130_fd_sc_hd__clkbuf_1
X_1440_ _0141_ vss vss vdd vdd _0837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_239 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_222 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1707_ _0237_ vss vss vdd vdd _0446_ sky130_fd_sc_hd__clkbuf_1
X_1638_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0214_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1569_ _0165_ vss vss vdd vdd _0809_ sky130_fd_sc_hd__inv_2
XTAP_294 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net21 sky130_fd_sc_hd__buf_4
Xfanout32 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out vss vss vdd vdd
+ net32 sky130_fd_sc_hd__clkbuf_4
Xfanout43 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out vss vss vdd vdd
+ net43 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_136 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_0940_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0337_ sky130_fd_sc_hd__inv_2
X_2541_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out _0787_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2610_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ _0856_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2472_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out _0718_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_1354_ _0112_ vss vss vdd vdd _0476_ sky130_fd_sc_hd__clkbuf_1
X_1423_ _0136_ vss vss vdd vdd _0498_ sky130_fd_sc_hd__clkbuf_1
X_1285_ _0087_ vss vss vdd vdd _0638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_194 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_32_150 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1070_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0323_
+ sky130_fd_sc_hd__clkbuf_1
X_1972_ clknet_4_1_0_prog_clk net180 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2524_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out _0770_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2455_ net60 _0701_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1337_ _0105_ vss vss vdd vdd _0835_ sky130_fd_sc_hd__clkbuf_1
X_1406_ _0129_ vss vss vdd vdd _0487_ sky130_fd_sc_hd__inv_2
Xhold19 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd net86 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out _0632_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1268_ _0080_ vss vss vdd vdd _0627_ sky130_fd_sc_hd__inv_2
X_1199_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0886_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_253 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_20_175 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2171_ net26 _0417_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1122_ _0028_ vss vss vdd vdd _0767_ sky130_fd_sc_hd__inv_2
X_2240_ net25 _0486_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1053_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd _0317_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_256 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1955_ clknet_4_5_0_prog_clk net207 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1886_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_22_61 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2438_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out _0684_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2507_ net27 _0753_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2369_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out _0615_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1671_ _0165_ vss vss vdd vdd _0806_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_16 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1740_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0545_
+ sky130_fd_sc_hd__inv_2
X_2223_ net36 _0469_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2154_ net34 _0400_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2085_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ _0331_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_1105_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0740_
+ sky130_fd_sc_hd__inv_2
X_1036_ _0311_ vss vss vdd vdd _0723_ sky130_fd_sc_hd__clkbuf_1
X_1938_ clknet_4_15_0_prog_clk net176 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1869_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_16_278 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold127 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd net194
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd net183
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q vss vss vdd vdd net172
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ _0212_ vss vss vdd vdd _0400_ sky130_fd_sc_hd__inv_2
X_1723_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0243_
+ sky130_fd_sc_hd__clkbuf_1
X_1585_ _0195_ vss vss vdd vdd _0196_ sky130_fd_sc_hd__clkbuf_1
X_2206_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out _0452_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_21_281 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2137_ net45 _0383_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1019_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q vss vss vdd vdd _0305_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_242 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_275 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1370_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0461_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_5_234 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1706_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0237_
+ sky130_fd_sc_hd__clkbuf_1
X_1637_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q vss vss vdd vdd _0409_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_5_278 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1568_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0815_ sky130_fd_sc_hd__inv_2
XTAP_295 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _0162_ vss vss vdd vdd _0163_ sky130_fd_sc_hd__clkbuf_1
Xfanout33 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out vss vss vdd vdd
+ net33 sky130_fd_sc_hd__clkbuf_2
Xfanout22 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net22 sky130_fd_sc_hd__buf_6
Xfanout44 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out vss vss vdd vdd
+ net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2540_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out _0786_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1422_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd _0136_
+ sky130_fd_sc_hd__clkbuf_1
X_2471_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out _0717_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1353_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0112_
+ sky130_fd_sc_hd__clkbuf_1
X_1284_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd _0087_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_71 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_33_129 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0999_ _0298_ vss vss vdd vdd _0692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_195 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_17_192 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_52 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1971_ clknet_4_1_0_prog_clk net191 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2523_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out _0769_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1405_ _0130_ vss vss vdd vdd _0501_ sky130_fd_sc_hd__clkbuf_1
X_2385_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out _0631_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2454_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out _0700_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_23_184 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1336_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0105_ sky130_fd_sc_hd__clkbuf_1
Xinput1 bottom_width_0_height_0_subtile_0__pin_I_2_ vss vss vdd vdd net1 sky130_fd_sc_hd__clkbuf_1
X_1198_ _0056_ vss vss vdd vdd _0873_ sky130_fd_sc_hd__clkbuf_1
X_1267_ _0081_ vss vss vdd vdd _0641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_265 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_46_232 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
X_1121_ _0029_ vss vss vdd vdd _0781_ sky130_fd_sc_hd__clkbuf_1
X_2170_ net21 _0416_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1052_ _0316_ vss vss vdd vdd _0726_ sky130_fd_sc_hd__clkbuf_1
X_1954_ clknet_4_5_0_prog_clk net165 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_148 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_22_40 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1885_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_11_132 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_2506_ net21 _0752_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2368_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out _0614_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_187 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2437_ net22 _0683_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1319_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0853_ sky130_fd_sc_hd__inv_2
X_2299_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out _0545_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1670_ _0224_ vss vss vdd vdd _0799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_202 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2222_ net40 _0468_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2153_ net38 _0399_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2084_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ _0330_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_7 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1035_ _0307_ vss vss vdd vdd _0311_ sky130_fd_sc_hd__clkbuf_1
X_1104_ _0012_ vss vss vdd vdd _0734_ sky130_fd_sc_hd__inv_2
X_1937_ clknet_4_15_0_prog_clk net146 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1799_ _0267_ vss vss vdd vdd _0779_ sky130_fd_sc_hd__clkbuf_1
X_1868_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ sky130_fd_sc_hd__inv_2
X_2399__58 vss vss vdd vdd net58 _2399__58/LO sky130_fd_sc_hd__conb_1
XFILLER_0_22_238 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_1584_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd _0195_
+ sky130_fd_sc_hd__buf_6
X_1653_ _0219_ vss vss vdd vdd _0414_ sky130_fd_sc_hd__clkbuf_1
Xhold128 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd net195
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd net173
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q vss vss vdd vdd net206
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q vss vss vdd vdd net184
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1722_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q vss vss vdd vdd _0549_
+ sky130_fd_sc_hd__inv_2
X_2205_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out _0451_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_44_93 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2136_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out _0382_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_1018_ _0304_ vss vss vdd vdd _0732_ sky130_fd_sc_hd__buf_1
XFILLER_0_8_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_39_124 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_219 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1705_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q vss vss vdd vdd _0436_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1567_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0818_ sky130_fd_sc_hd__inv_2
X_1636_ _0212_ vss vss vdd vdd _0403_ sky130_fd_sc_hd__inv_2
XTAP_241 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ net48 _0365_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_296 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd _0162_
+ sky130_fd_sc_hd__buf_6
Xfanout23 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net23 sky130_fd_sc_hd__buf_2
Xfanout45 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out vss vss vdd vdd
+ net45 sky130_fd_sc_hd__clkbuf_2
Xfanout34 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out vss vss vdd vdd
+ net34 sky130_fd_sc_hd__clkbuf_4
X_1421_ _0135_ vss vss vdd vdd _0503_ sky130_fd_sc_hd__clkbuf_1
X_2470_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out _0716_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1352_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q vss vss vdd vdd _0465_
+ sky130_fd_sc_hd__inv_2
X_1283_ _0086_ vss vss vdd vdd _0643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_174 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_33_108 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0998_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd _0298_
+ sky130_fd_sc_hd__clkbuf_1
X_1619_ _0195_ vss vss vdd vdd _0369_ sky130_fd_sc_hd__inv_2
X_2599_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ _0845_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_24_108 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1970_ clknet_4_0_0_prog_clk net162 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2522_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out _0768_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1335_ _0104_ vss vss vdd vdd _0830_ sky130_fd_sc_hd__clkbuf_1
X_1404_ _0129_ vss vss vdd vdd _0130_ sky130_fd_sc_hd__clkbuf_1
X_2384_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out _0630_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2453_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out _0699_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput2 bottom_width_0_height_0_subtile_0__pin_I_6_ vss vss vdd vdd net2 sky130_fd_sc_hd__buf_1
X_1197_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0056_ sky130_fd_sc_hd__clkbuf_1
X_1266_ _0080_ vss vss vdd vdd _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_130 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_14_141 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_174 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_32_19 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_37_255 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_166 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1120_ _0028_ vss vss vdd vdd _0029_ sky130_fd_sc_hd__clkbuf_1
X_1051_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0316_
+ sky130_fd_sc_hd__clkbuf_1
X_1953_ clknet_4_7_0_prog_clk net76 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_222 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_28_200 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1884_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_43_236 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2505_ net29 _0751_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_144 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_11_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1318_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0854_ sky130_fd_sc_hd__inv_2
X_2367_ net26 _0613_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2436_ net24 _0682_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2298_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out _0544_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1249_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd _0074_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_73 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_225 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_25_269 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2221_ net44 _0467_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2152_ net42 _0398_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2083_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ _0329_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_85 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1034_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0714_
+ sky130_fd_sc_hd__inv_2
X_1103_ _0022_ vss vss vdd vdd _0748_ sky130_fd_sc_hd__clkbuf_1
X_1867_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ sky130_fd_sc_hd__inv_2
X_1936_ _0002_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ _0000_ _0001_ vss vss vdd vdd _1936_/Q logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ sky130_fd_sc_hd__dfbbn_1
XFILLER_0_16_236 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1798_ _0028_ vss vss vdd vdd _0267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_239 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2419_ net37 _0665_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_30_294 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1721_ _0242_ vss vss vdd vdd _0824_ sky130_fd_sc_hd__buf_1
X_1583_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0379_
+ sky130_fd_sc_hd__inv_2
Xhold107 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q vss vss vdd vdd net174
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd _0219_
+ sky130_fd_sc_hd__clkbuf_1
Xhold118 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd net185
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd net196
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2135_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out _0381_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2204_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out _0450_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1017_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q vss vss vdd vdd _0304_
+ sky130_fd_sc_hd__clkbuf_1
X_1919_ clknet_4_8_0_prog_clk net136 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_72 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_8_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_39_169 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_14_42 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1704_ _0228_ vss vss vdd vdd _0427_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_2_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1566_ _0188_ vss vss vdd vdd _0805_ sky130_fd_sc_hd__clkbuf_1
X_1635_ _0213_ vss vss vdd vdd _0417_ sky130_fd_sc_hd__clkbuf_1
XTAP_275 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0547_
+ sky130_fd_sc_hd__inv_2
X_2118_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out _0364_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_297 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ clknet_4_2_0_prog_clk net124 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ sky130_fd_sc_hd__dfxtp_1
Xfanout46 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out vss vss vdd vdd
+ net46 sky130_fd_sc_hd__clkbuf_4
Xfanout24 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net24 sky130_fd_sc_hd__buf_6
Xfanout35 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out vss vss vdd vdd
+ net35 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_161 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1351_ _0110_ vss vss vdd vdd _0459_ sky130_fd_sc_hd__inv_2
X_1420_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0135_
+ sky130_fd_sc_hd__clkbuf_1
X_1282_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0086_
+ sky130_fd_sc_hd__clkbuf_1
X_1618_ _0206_ vss vss vdd vdd _0383_ sky130_fd_sc_hd__clkbuf_1
X_0997_ _0297_ vss vss vdd vdd _0698_ sky130_fd_sc_hd__clkbuf_1
X_1549_ _0181_ vss vss vdd vdd _0366_ sky130_fd_sc_hd__clkbuf_1
X_2598_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ _0844_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_32_164 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_46_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2521_ net23 _0767_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_23_164 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1334_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0104_ sky130_fd_sc_hd__clkbuf_1
X_1403_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd _0129_
+ sky130_fd_sc_hd__buf_6
X_1265_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd _0080_
+ sky130_fd_sc_hd__buf_6
X_2383_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out _0629_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2452_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out _0698_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2371__57 vss vss vdd vdd net57 _2371__57/LO sky130_fd_sc_hd__conb_1
Xinput3 ccff_head vss vss vdd vdd net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ _0044_ vss vss vdd vdd _0565_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_153 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1050_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q vss vss vdd vdd _0716_
+ sky130_fd_sc_hd__inv_2
X_1952_ clknet_4_7_0_prog_clk net186 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1883_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ sky130_fd_sc_hd__inv_2
X_2435_ net31 _0681_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2504_ net32 _0750_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1317_ _0098_ vss vss vdd vdd _0823_ sky130_fd_sc_hd__clkbuf_1
X_2297_ net22 _0543_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1248_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0600_
+ sky130_fd_sc_hd__inv_2
X_2366_ net20 _0612_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1179_ _0050_ vss vss vdd vdd _0587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_15_0_prog_clk sky130_fd_sc_hd__clkbuf_8
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2220_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out _0466_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
X_2151_ net47 _0397_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1102_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q vss vss vdd vdd _0022_
+ sky130_fd_sc_hd__clkbuf_1
X_2082_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ _0328_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_33_52 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_17_75 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1033_ _0307_ vss vss vdd vdd _0710_ sky130_fd_sc_hd__inv_2
X_1797_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0770_
+ sky130_fd_sc_hd__inv_2
X_1935_ clknet_4_13_0_prog_clk net79 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1866_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ sky130_fd_sc_hd__inv_2
X_2418_ net41 _0664_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2349_ net38 _0595_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_38_19 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold108 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q vss vss vdd vdd net175
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1720_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ vss vss vdd vdd _0242_ sky130_fd_sc_hd__clkbuf_1
X_1651_ _0218_ vss vss vdd vdd _0419_ sky130_fd_sc_hd__clkbuf_1
X_1582_ _0194_ vss vss vdd vdd _0393_ sky130_fd_sc_hd__clkbuf_1
Xhold119 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q vss vss vdd vdd net186
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2203_ net51 _0449_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2134_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out _0380_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1016_ _0303_ vss vss vdd vdd _0895_ sky130_fd_sc_hd__clkbuf_1
X_1849_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ sky130_fd_sc_hd__inv_2
X_1918_ clknet_4_10_0_prog_clk net68 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
X_1703_ _0236_ vss vss vdd vdd _0441_ sky130_fd_sc_hd__clkbuf_1
X_1634_ _0212_ vss vss vdd vdd _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_259 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1565_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0188_ sky130_fd_sc_hd__clkbuf_1
XTAP_298 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _0161_ vss vss vdd vdd _0561_ sky130_fd_sc_hd__clkbuf_1
X_2117_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out _0363_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2048_ clknet_4_2_0_prog_clk net120 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_3 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xfanout47 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out vss vss vdd vdd
+ net47 sky130_fd_sc_hd__clkbuf_2
Xfanout36 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out vss vss vdd vdd
+ net36 sky130_fd_sc_hd__clkbuf_4
Xfanout25 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net25 sky130_fd_sc_hd__buf_2
XFILLER_0_3_6 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_35_140 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1350_ _0111_ vss vss vdd vdd _0473_ sky130_fd_sc_hd__clkbuf_1
X_1281_ _0085_ vss vss vdd vdd _0646_ sky130_fd_sc_hd__clkbuf_1
X_0996_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0297_
+ sky130_fd_sc_hd__clkbuf_1
X_1617_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd _0206_
+ sky130_fd_sc_hd__clkbuf_1
X_2597_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ _0843_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_1548_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q vss vss vdd vdd _0181_
+ sky130_fd_sc_hd__clkbuf_1
X_1479_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0155_
+ sky130_fd_sc_hd__clkbuf_1
X_2520_ net25 _0766_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1402_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0491_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_11_44 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2451_ net27 _0697_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_1333_ _0099_ vss vss vdd vdd _0845_ sky130_fd_sc_hd__inv_2
X_2382_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out _0628_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1264_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0631_
+ sky130_fd_sc_hd__inv_2
Xinput4 clk vss vss vdd vdd net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_74 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1195_ _0055_ vss vss vdd vdd _0579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0979_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0686_
+ sky130_fd_sc_hd__inv_2
X_2649_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ _0895_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_37_202 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1951_ clknet_4_7_0_prog_clk net200 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1882_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_7_129 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2434_ net35 _0680_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2365_ net28 _0611_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2503_ net36 _0749_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1316_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0098_ sky130_fd_sc_hd__clkbuf_1
X_2296_ net24 _0542_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1247_ _0063_ vss vss vdd vdd _0594_ sky130_fd_sc_hd__inv_2
X_1178_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0050_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_216 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_173 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2150_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out _0396_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_1032_ _0310_ vss vss vdd vdd _0724_ sky130_fd_sc_hd__clkbuf_1
X_2081_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
+ _0327_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ sky130_fd_sc_hd__ebufn_1
X_1101_ _0021_ vss vss vdd vdd _0754_ sky130_fd_sc_hd__clkbuf_1
X_1934_ clknet_4_12_0_prog_clk net205 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
X_1865_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ sky130_fd_sc_hd__inv_2
X_1796_ _0266_ vss vss vdd vdd _0892_ sky130_fd_sc_hd__buf_1
XFILLER_0_42_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2417_ net44 _0663_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2348_ net42 _0594_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2279_ net36 _0525_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_30_285 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1581_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0194_
+ sky130_fd_sc_hd__clkbuf_1
Xhold109 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd net176
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1650_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0218_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_230 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_2202_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out _0448_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2133_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out _0379_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_44_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1015_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_7 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_1917_ net4 vss vss vdd vdd _0011_ sky130_fd_sc_hd__inv_2
X_1848_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_8_63 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1779_ _0261_ vss vss vdd vdd _0665_ sky130_fd_sc_hd__clkbuf_1
X_1702_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd _0236_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_41 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1564_ _0187_ vss vss vdd vdd _0355_ sky130_fd_sc_hd__clkbuf_1
X_1633_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd _0212_
+ sky130_fd_sc_hd__buf_6
XTAP_299 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0161_
+ sky130_fd_sc_hd__clkbuf_1
Xfanout26 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net26 sky130_fd_sc_hd__buf_6
X_2116_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out _0362_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2047_ clknet_4_0_0_prog_clk net73 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ sky130_fd_sc_hd__dfxtp_1
Xfanout37 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out vss vss vdd vdd
+ net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1280_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q vss vss vdd vdd _0085_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_65 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_25_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0995_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q vss vss vdd vdd _0688_
+ sky130_fd_sc_hd__inv_2
X_1547_ net16 vss vss vdd vdd _0354_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1616_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0376_
+ sky130_fd_sc_hd__inv_2
X_2596_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ _0842_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_5_86 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1478_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q vss vss vdd vdd _0520_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_23_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1401_ _0128_ vss vss vdd vdd _0505_ sky130_fd_sc_hd__clkbuf_1
X_2381_ net22 _0627_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2450_ net21 _0696_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput5 left_width_0_height_0_subtile_0__pin_I_3_ vss vss vdd vdd net5 sky130_fd_sc_hd__clkbuf_1
X_1332_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0850_ sky130_fd_sc_hd__inv_2
X_1263_ _0079_ vss vss vdd vdd _0645_ sky130_fd_sc_hd__clkbuf_1
X_1194_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd _0055_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_225 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XTAP_94 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_166 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_0978_ _0288_ vss vss vdd vdd _0682_ sky130_fd_sc_hd__inv_2
X_2648_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ _0894_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_2579_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ _0825_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1950_ clknet_4_7_0_prog_clk net156 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1881_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_22_44 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2502_ net41 _0748_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1315_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ vss vss vdd vdd _0822_ sky130_fd_sc_hd__inv_2
X_2364_ net32 _0610_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_169 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2433_ net39 _0679_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2295_ net30 _0541_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1246_ _0073_ vss vss vdd vdd _0608_ sky130_fd_sc_hd__clkbuf_1
X_1177_ _0049_ vss vss vdd vdd _0590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2080_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
+ _0326_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_1100_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0021_
+ sky130_fd_sc_hd__clkbuf_1
X_1031_ _0307_ vss vss vdd vdd _0310_ sky130_fd_sc_hd__clkbuf_1
X_1933_ clknet_4_15_0_prog_clk net3 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_272 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_24_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_3_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1795_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ vss vss vdd vdd _0266_ sky130_fd_sc_hd__clkbuf_1
X_1864_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_35_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2416_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out _0662_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2347_ net46 _0593_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2278_ net40 _0524_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1229_ _0063_ vss vss vdd vdd _0597_ sky130_fd_sc_hd__inv_2
X_1580_ _0193_ vss vss vdd vdd _0395_ sky130_fd_sc_hd__clkbuf_1
X_2132_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out _0378_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2201_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out _0447_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1014_ _0277_ vss vss vdd vdd _0326_ sky130_fd_sc_hd__inv_2
X_1847_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
+ sky130_fd_sc_hd__inv_2
X_1916_ net4 vss vss vdd vdd _0008_ sky130_fd_sc_hd__inv_2
X_1778_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd _0261_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1701_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0433_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_38_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_14_89 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1563_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd _0187_
+ sky130_fd_sc_hd__clkbuf_1
X_1632_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0407_
+ sky130_fd_sc_hd__inv_2
XTAP_223 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _0160_ vss vss vdd vdd _0563_ sky130_fd_sc_hd__clkbuf_1
X_2115_ net26 _0361_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_289 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout38 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out vss vss vdd vdd
+ net38 sky130_fd_sc_hd__clkbuf_4
Xfanout27 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ vss vss vdd vdd net27 sky130_fd_sc_hd__buf_2
X_2046_ clknet_4_0_0_prog_clk net135 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_175 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_41_76 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0994_ _0288_ vss vss vdd vdd _0679_ sky130_fd_sc_hd__inv_2
X_1546_ _0180_ vss vss vdd vdd _0359_ sky130_fd_sc_hd__clkbuf_1
X_1615_ _0195_ vss vss vdd vdd _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1477_ _0146_ vss vss vdd vdd _0511_ sky130_fd_sc_hd__inv_2
X_2595_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ _0841_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_2029_ clknet_4_4_0_prog_clk net95 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_1_0_prog_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1400_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0128_
+ sky130_fd_sc_hd__clkbuf_1
X_1331_ _0103_ vss vss vdd vdd _0838_ sky130_fd_sc_hd__clkbuf_1
X_2380_ net24 _0626_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput6 left_width_0_height_0_subtile_0__pin_I_7_ vss vss vdd vdd net6 sky130_fd_sc_hd__clkbuf_1
X_1262_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0079_
+ sky130_fd_sc_hd__clkbuf_1
X_1193_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0572_
+ sky130_fd_sc_hd__inv_2
XTAP_95 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_112 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_134 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2647_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ _0893_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0977_ _0291_ vss vss vdd vdd _0696_ sky130_fd_sc_hd__clkbuf_1
X_1529_ _0173_ vss vss vdd vdd _0368_ sky130_fd_sc_hd__clkbuf_1
X_2578_ net65 _0824_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_2259__53 vss vss vdd vdd net53 _2259__53/LO sky130_fd_sc_hd__conb_1
XPHY_90 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1880_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__inv_2
X_2501_ net45 _0747_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2432_ net43 _0678_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2363_ net36 _0609_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1314_ _0096_ vss vss vdd vdd _0655_ sky130_fd_sc_hd__inv_2
X_2294_ net34 _0540_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1245_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd _0073_
+ sky130_fd_sc_hd__clkbuf_1
X_1176_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q vss vss vdd vdd _0049_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_259 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1030_ _0309_ vss vss vdd vdd _0728_ sky130_fd_sc_hd__clkbuf_1
X_1932_ clknet_4_11_0_prog_clk net151 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1863_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__inv_2
X_1794_ _0028_ vss vss vdd vdd _0766_ sky130_fd_sc_hd__inv_2
X_2415_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out _0661_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2346_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out _0592_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
X_1228_ _0067_ vss vss vdd vdd _0611_ sky130_fd_sc_hd__clkbuf_1
X_2277_ net44 _0523_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1159_ _0043_ vss vss vdd vdd _0589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_262 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_159 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2131_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out _0377_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2200_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out _0446_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_28_99 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_28_44 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_1013_ _0302_ vss vss vdd vdd _0902_ sky130_fd_sc_hd__buf_1
X_1846_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__inv_2
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_14_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1915_ net4 vss vss vdd vdd _0005_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_43 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_259 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1777_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0657_
+ sky130_fd_sc_hd__inv_2
X_2329_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out _0575_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1700_ _0228_ vss vss vdd vdd _0428_ sky130_fd_sc_hd__inv_2
X_1631_ _0211_ vss vss vdd vdd _0421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_56 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_39_76 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1562_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0348_
+ sky130_fd_sc_hd__inv_2
XTAP_257 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q vss vss vdd vdd _0160_
+ sky130_fd_sc_hd__clkbuf_1
X_2114_ net20 _0360_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_279 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ clknet_4_0_0_prog_clk net117 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ sky130_fd_sc_hd__dfxtp_1
Xfanout39 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out vss vss vdd vdd
+ net39 sky130_fd_sc_hd__clkbuf_2
Xfanout28 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out vss vss vdd vdd
+ net28 sky130_fd_sc_hd__clkbuf_4
X_1829_ _0176_ vss vss vdd vdd _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_198 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_35_165 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_25_34 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_41_11 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_78 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_0993_ _0296_ vss vss vdd vdd _0693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_179 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1614_ _0205_ vss vss vdd vdd _0384_ sky130_fd_sc_hd__clkbuf_1
X_2594_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ _0840_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1545_ _0176_ vss vss vdd vdd _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_66 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1476_ _0154_ vss vss vdd vdd _0525_ sky130_fd_sc_hd__clkbuf_1
X_2028_ clknet_4_4_0_prog_clk net86 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_121 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_23_135 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1330_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0103_ sky130_fd_sc_hd__clkbuf_1
X_1261_ _0078_ vss vss vdd vdd _0647_ sky130_fd_sc_hd__clkbuf_1
Xinput7 reset vss vss vdd vdd net7 sky130_fd_sc_hd__clkbuf_4
X_1192_ _0044_ vss vss vdd vdd _0566_ sky130_fd_sc_hd__inv_2
XTAP_96 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0976_ _0288_ vss vss vdd vdd _0291_ sky130_fd_sc_hd__clkbuf_1
X_2577_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ _0823_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_2646_ net67 _0892_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1528_ net16 vss vss vdd vdd _0173_ sky130_fd_sc_hd__clkbuf_1
X_1459_ _0146_ vss vss vdd vdd _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_91 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_80 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2431_ net46 _0677_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2500_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out _0746_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_2362_ net40 _0608_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1244_ _0072_ vss vss vdd vdd _0614_ sky130_fd_sc_hd__clkbuf_1
X_1313_ _0097_ vss vss vdd vdd _0669_ sky130_fd_sc_hd__clkbuf_1
X_2293_ net38 _0539_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1175_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q vss vss vdd vdd _0578_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_42_241 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0959_ _0277_ vss vss vdd vdd _0328_ sky130_fd_sc_hd__inv_2
X_2629_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ _0875_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_25_208 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_17_68 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_33_78 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput10 right_width_0_height_0_subtile_0__pin_I_9_ vss vss vdd vdd net10 sky130_fd_sc_hd__clkbuf_1
X_1793_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0855_ sky130_fd_sc_hd__inv_2
X_1931_ clknet_4_11_0_prog_clk net106 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1862_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__inv_2
X_2414_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out _0660_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1158_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0043_
+ sky130_fd_sc_hd__clkbuf_1
X_2345_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out _0591_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1227_ _0063_ vss vss vdd vdd _0067_ sky130_fd_sc_hd__clkbuf_1
X_2276_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out _0522_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_1089_ _0017_ vss vss vdd vdd _0758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_23 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_0_105 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_44_22 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2130_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out _0376_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_28_56 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1012_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0302_ sky130_fd_sc_hd__buf_1
XFILLER_0_44_77 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1914_ net4 vss vss vdd vdd _0002_ sky130_fd_sc_hd__inv_2
X_1845_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_8_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1776_ _0096_ vss vss vdd vdd _0652_ sky130_fd_sc_hd__inv_2
X_2328_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out _0574_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2259_ net53 _0505_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1630_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0211_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_13 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_39_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1561_ _0186_ vss vss vdd vdd _0356_ sky130_fd_sc_hd__clkbuf_1
XTAP_269 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _0159_ vss vss vdd vdd _0564_ sky130_fd_sc_hd__buf_1
X_2113_ net29 _0359_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2044_ clknet_4_0_0_prog_clk net115 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_7 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_44_122 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xfanout29 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out vss vss vdd vdd
+ net29 sky130_fd_sc_hd__buf_2
X_2231__52 vss vss vdd vdd net52 _2231__52/LO sky130_fd_sc_hd__conb_1
X_1828_ _0176_ vss vss vdd vdd _0343_ sky130_fd_sc_hd__inv_2
X_1759_ _0254_ vss vss vdd vdd _0672_ sky130_fd_sc_hd__clkbuf_1
X_2455__60 vss vss vdd vdd net60 _2455__60/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_46 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_41_67 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_0992_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd _0296_
+ sky130_fd_sc_hd__clkbuf_1
X_1544_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0350_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_41_169 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1613_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd _0205_
+ sky130_fd_sc_hd__clkbuf_1
X_2593_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ _0839_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_26_177 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1475_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd _0154_
+ sky130_fd_sc_hd__clkbuf_1
X_2027_ clknet_4_4_0_prog_clk net108 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_103 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_17_133 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_40_180 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1260_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q vss vss vdd vdd _0078_
+ sky130_fd_sc_hd__clkbuf_1
X_1191_ _0054_ vss vss vdd vdd _0580_ sky130_fd_sc_hd__clkbuf_1
Xinput8 right_width_0_height_0_subtile_0__pin_I_1_ vss vss vdd vdd net8 sky130_fd_sc_hd__buf_1
XFILLER_0_46_206 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_97 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ _0290_ vss vss vdd vdd _0700_ sky130_fd_sc_hd__clkbuf_1
X_1527_ _0172_ vss vss vdd vdd _0795_ sky130_fd_sc_hd__clkbuf_1
X_2576_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ _0822_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2645_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ _0891_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_1389_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0123_ sky130_fd_sc_hd__clkbuf_1
X_1458_ _0148_ vss vss vdd vdd _0532_ sky130_fd_sc_hd__clkbuf_1
XPHY_92 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_43_209 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_81 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_36_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_70 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2361_ net44 _0607_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2430_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out _0676_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1243_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0072_
+ sky130_fd_sc_hd__clkbuf_1
X_1312_ _0096_ vss vss vdd vdd _0097_ sky130_fd_sc_hd__clkbuf_1
X_1174_ _0044_ vss vss vdd vdd _0569_ sky130_fd_sc_hd__inv_2
X_2292_ net42 _0538_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0958_ _0283_ vss vss vdd vdd _0903_ sky130_fd_sc_hd__buf_1
X_2559_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ _0805_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
X_2628_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ _0874_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_18_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_33_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1930_ clknet_4_11_0_prog_clk net91 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1792_ _0265_ vss vss vdd vdd _0859_ sky130_fd_sc_hd__clkbuf_1
Xinput11 set vss vss vdd vdd net11 sky130_fd_sc_hd__clkbuf_2
X_1861_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__inv_2
X_2413_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out _0659_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2344_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out _0590_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1157_ _0042_ vss vss vdd vdd _0591_ sky130_fd_sc_hd__clkbuf_1
X_1226_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0602_
+ sky130_fd_sc_hd__inv_2
X_2275_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out _0521_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1088_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q vss vss vdd vdd _0017_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_191 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_278 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_44_56 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1011_ _0301_ vss vss vdd vdd _0896_ sky130_fd_sc_hd__clkbuf_1
X_1913_ _0176_ vss vss vdd vdd _0346_ sky130_fd_sc_hd__inv_2
X_1844_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__inv_2
X_1775_ _0260_ vss vss vdd vdd _0666_ sky130_fd_sc_hd__clkbuf_1
X_2258_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out _0504_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2327_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out _0573_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2189_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out _0435_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1209_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q vss vss vdd vdd _0060_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_186 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1560_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd _0186_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_89 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2112_ net33 _0358_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_259 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q vss vss vdd vdd _0159_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_215 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ clknet_4_0_0_prog_clk net121 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1827_ _0176_ vss vss vdd vdd _0344_ sky130_fd_sc_hd__inv_2
X_1689_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0434_
+ sky130_fd_sc_hd__inv_2
X_1758_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0254_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_69 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_167 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_26_101 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2661_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ _0907_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
X_0991_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0685_
+ sky130_fd_sc_hd__inv_2
X_1543_ _0179_ vss vss vdd vdd _0360_ sky130_fd_sc_hd__clkbuf_1
X_1612_ _0204_ vss vss vdd vdd _0390_ sky130_fd_sc_hd__clkbuf_1
X_2592_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ _0838_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_1474_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0517_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2026_ clknet_4_4_0_prog_clk net81 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_101 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_40_192 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_40_170 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput9 right_width_0_height_0_subtile_0__pin_I_5_ vss vss vdd vdd net9 sky130_fd_sc_hd__clkbuf_1
X_1190_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd _0054_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_98 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2644_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ _0890_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_0974_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0290_
+ sky130_fd_sc_hd__clkbuf_1
X_1526_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0172_ sky130_fd_sc_hd__clkbuf_1
X_2575_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ _0821_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1457_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0148_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_192 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1388_ _0099_ vss vss vdd vdd _0843_ sky130_fd_sc_hd__inv_2
X_2009_ clknet_4_7_0_prog_clk net109 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_295 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_82 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_71 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_60 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_28_218 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_93 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_22_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1311_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd _0096_
+ sky130_fd_sc_hd__buf_6
X_2360_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out _0606_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_2291_ net46 _0537_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1242_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q vss vss vdd vdd _0604_
+ sky130_fd_sc_hd__inv_2
X_1173_ _0048_ vss vss vdd vdd _0583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_221 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_0957_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0283_ sky130_fd_sc_hd__buf_1
X_2627_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ _0873_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_0_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_2558_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ _0804_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_1509_ _0165_ vss vss vdd vdd _0813_ sky130_fd_sc_hd__inv_2
X_2489_ net39 _0735_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1860_ net23 vss vss vdd vdd net19 sky130_fd_sc_hd__inv_2
XFILLER_0_33_25 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput12 top_width_0_height_0_subtile_0__pin_I_0_ vss vss vdd vdd net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1791_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_8 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2343_ net56 _0589_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2412_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out _0658_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2274_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out _0520_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1156_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q vss vss vdd vdd _0042_
+ sky130_fd_sc_hd__clkbuf_1
X_1225_ _0063_ vss vss vdd vdd _0598_ sky130_fd_sc_hd__inv_2
X_1087_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q vss vss vdd vdd _0746_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_15_232 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1989_ clknet_4_14_0_prog_clk net129 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1010_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0301_ sky130_fd_sc_hd__clkbuf_1
X_1843_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__inv_2
X_1912_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_8_79 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1774_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd _0260_
+ sky130_fd_sc_hd__clkbuf_1
X_2257_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out _0503_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_26_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1208_ _0059_ vss vss vdd vdd _0861_ sky130_fd_sc_hd__clkbuf_1
X_2326_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out _0572_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2188_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out _0434_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1139_ _0035_ vss vss vdd vdd _0870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_46 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1490_ _0099_ vss vss vdd vdd _0840_ sky130_fd_sc_hd__inv_2
XTAP_205 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ net37 _0357_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_249 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2042_ clknet_4_0_0_prog_clk net122 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ sky130_fd_sc_hd__dfxtp_1
Xhold1 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd net68 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1826_ _0176_ vss vss vdd vdd _0345_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_232 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1688_ _0228_ vss vss vdd vdd _0430_ sky130_fd_sc_hd__inv_2
X_1757_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q vss vss vdd vdd _0661_
+ sky130_fd_sc_hd__inv_2
X_2309_ net28 _0555_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_35_146 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_35_179 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_13_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1611_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0204_
+ sky130_fd_sc_hd__clkbuf_1
X_2660_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ _0906_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_0990_ _0288_ vss vss vdd vdd _0680_ sky130_fd_sc_hd__inv_2
X_1542_ _0176_ vss vss vdd vdd _0179_ sky130_fd_sc_hd__clkbuf_1
X_2591_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ _0837_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_1473_ _0146_ vss vss vdd vdd _0512_ sky130_fd_sc_hd__inv_2
X_2025_ clknet_4_5_0_prog_clk net71 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1809_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0769_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_157 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_28 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_36_69 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_99 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2574_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ _0820_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_8
X_2643_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ _0889_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_0973_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q vss vss vdd vdd _0689_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1525_ _0165_ vss vss vdd vdd _0810_ sky130_fd_sc_hd__inv_2
X_1387_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0849_ sky130_fd_sc_hd__inv_2
X_1456_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q vss vss vdd vdd _0521_
+ sky130_fd_sc_hd__inv_2
X_2008_ clknet_4_7_0_prog_clk net104 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_121 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_83 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_72 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_61 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_50 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_11_108 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_119 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1241_ _0063_ vss vss vdd vdd _0595_ sky130_fd_sc_hd__inv_2
X_1310_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0659_
+ sky130_fd_sc_hd__inv_2
X_2290_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out _0536_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_1172_ _0044_ vss vss vdd vdd _0048_ sky130_fd_sc_hd__clkbuf_1
X_0956_ _0282_ vss vss vdd vdd _0898_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_219 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2557_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ _0803_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_2626_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ _0872_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1508_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0165_ sky130_fd_sc_hd__buf_6
X_1439_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0141_ sky130_fd_sc_hd__clkbuf_1
X_2488_ net43 _0734_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xinput13 top_width_0_height_0_subtile_0__pin_I_4_ vss vss vdd vdd net13 sky130_fd_sc_hd__clkbuf_1
X_1790_ _0096_ vss vss vdd vdd _0649_ sky130_fd_sc_hd__inv_2
X_2411_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out _0657_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1224_ _0066_ vss vss vdd vdd _0612_ sky130_fd_sc_hd__clkbuf_1
X_2342_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out _0588_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2273_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out _0519_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1086_ _0012_ vss vss vdd vdd _0737_ sky130_fd_sc_hd__inv_2
X_1155_ _0041_ vss vss vdd vdd _0592_ sky130_fd_sc_hd__clkbuf_1
X_1988_ clknet_4_10_0_prog_clk net189 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_0939_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0338_ sky130_fd_sc_hd__inv_2
X_2609_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ _0855_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_21_225 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_208 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1842_ net27 vss vss vdd vdd net18 sky130_fd_sc_hd__inv_2
X_1911_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ sky130_fd_sc_hd__inv_2
X_1773_ _0259_ vss vss vdd vdd _0671_ sky130_fd_sc_hd__clkbuf_1
X_2187_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out _0433_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2256_ logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out _0502_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1207_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0059_ sky130_fd_sc_hd__clkbuf_1
X_2325_ net22 _0571_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1138_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0035_ sky130_fd_sc_hd__clkbuf_1
X_1069_ _0322_ vss vss vdd vdd _0759_ sky130_fd_sc_hd__clkbuf_1
XTAP_239 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ net40 _0356_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2041_ clknet_4_0_0_prog_clk net114 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ sky130_fd_sc_hd__dfxtp_1
Xhold2 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ vss vss vdd vdd net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_133 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_1756_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0821_ sky130_fd_sc_hd__inv_2
X_1825_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0889_ sky130_fd_sc_hd__inv_2
X_1687_ _0231_ vss vss vdd vdd _0444_ sky130_fd_sc_hd__clkbuf_1
X_2308_ net32 _0554_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2239_ net30 _0485_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_35_169 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_1610_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q vss vss vdd vdd _0380_
+ sky130_fd_sc_hd__inv_2
X_2590_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ _0836_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_26_158 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1541_ _0178_ vss vss vdd vdd _0364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_48 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_37 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1472_ _0153_ vss vss vdd vdd _0526_ sky130_fd_sc_hd__clkbuf_1
X_2024_ clknet_4_5_0_prog_clk net102 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_169 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_40_161 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1808_ _0028_ vss vss vdd vdd _0764_ sky130_fd_sc_hd__inv_2
X_1739_ _0162_ vss vss vdd vdd _0540_ sky130_fd_sc_hd__inv_2
X_0972_ _0288_ vss vss vdd vdd _0683_ sky130_fd_sc_hd__inv_2
X_1524_ _0171_ vss vss vdd vdd _0801_ sky130_fd_sc_hd__clkbuf_1
X_2573_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ _0819_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_4
X_2642_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ _0888_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
X_1386_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0852_ sky130_fd_sc_hd__inv_2
X_1455_ _0146_ vss vss vdd vdd _0515_ sky130_fd_sc_hd__inv_2
X_2007_ clknet_4_13_0_prog_clk net92 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_92 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_45_231 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_84 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_73 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_62 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_51 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_40 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1240_ _0071_ vss vss vdd vdd _0609_ sky130_fd_sc_hd__clkbuf_1
X_1171_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0574_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_27_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0955_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0282_ sky130_fd_sc_hd__clkbuf_1
X_2556_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ _0802_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_1507_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0817_ sky130_fd_sc_hd__inv_2
X_2487_ net47 _0733_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2625_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ _0871_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_175 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_186 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1369_ _0110_ vss vss vdd vdd _0456_ sky130_fd_sc_hd__inv_2
X_1438_ _0129_ vss vss vdd vdd _0481_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_253 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xinput14 top_width_0_height_0_subtile_0__pin_I_8_ vss vss vdd vdd net14 sky130_fd_sc_hd__clkbuf_1
X_2410_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out _0656_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2341_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out _0587_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1154_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q vss vss vdd vdd _0041_
+ sky130_fd_sc_hd__clkbuf_1
X_1223_ _0063_ vss vss vdd vdd _0066_ sky130_fd_sc_hd__clkbuf_1
X_2272_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out _0518_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1085_ _0016_ vss vss vdd vdd _0751_ sky130_fd_sc_hd__clkbuf_1
X_1987_ clknet_4_10_0_prog_clk net164 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_0938_ _0276_ vss vss vdd vdd _0891_ sky130_fd_sc_hd__clkbuf_1
X_2608_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ _0854_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
X_2539_ net63 _0785_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_44_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_44_15 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_28_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1910_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ sky130_fd_sc_hd__inv_2
X_1841_ net10 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out
+ sky130_fd_sc_hd__inv_2
X_1772_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0259_
+ sky130_fd_sc_hd__clkbuf_1
X_2324_ net24 _0570_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2186_ logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out _0432_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2255_ net26 _0501_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1137_ _0034_ vss vss vdd vdd _0866_ sky130_fd_sc_hd__clkbuf_1
X_1206_ _0033_ vss vss vdd vdd _0876_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_253 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1068_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q vss vss vdd vdd _0322_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2147__49 vss vss vdd vdd net49 _2147__49/LO sky130_fd_sc_hd__conb_1
XFILLER_0_11_281 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_229 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd net70 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ clknet_4_0_0_prog_clk net103 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_29_145 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1686_ _0228_ vss vss vdd vdd _0231_ sky130_fd_sc_hd__clkbuf_1
X_1824_ _0275_ vss vss vdd vdd _0893_ sky130_fd_sc_hd__clkbuf_1
X_1755_ _0253_ vss vss vdd vdd _0825_ sky130_fd_sc_hd__clkbuf_1
X_2238_ net34 _0484_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2307_ net36 _0553_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_91 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2169_ net28 _0415_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_41_16 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1540_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0178_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_27 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1471_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd _0153_
+ sky130_fd_sc_hd__clkbuf_1
X_2023_ clknet_4_5_0_prog_clk net97 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1807_ _0270_ vss vss vdd vdd _0778_ sky130_fd_sc_hd__clkbuf_1
X_1669_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0224_ sky130_fd_sc_hd__clkbuf_1
X_1738_ _0248_ vss vss vdd vdd _0554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_107 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_0971_ _0289_ vss vss vdd vdd _0697_ sky130_fd_sc_hd__clkbuf_1
X_1523_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0171_ sky130_fd_sc_hd__clkbuf_1
X_2572_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ _0818_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_2641_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ _0887_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_1454_ _0147_ vss vss vdd vdd _0529_ sky130_fd_sc_hd__clkbuf_1
X_1385_ _0122_ vss vss vdd vdd _0839_ sky130_fd_sc_hd__clkbuf_1
X_2006_ clknet_4_13_0_prog_clk net80 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ sky130_fd_sc_hd__dfxtp_1
XPHY_30 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_85 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_74 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_63 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_52 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1170_ _0044_ vss vss vdd vdd _0570_ sky130_fd_sc_hd__inv_2
X_2624_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ _0870_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_0954_ _0277_ vss vss vdd vdd _0329_ sky130_fd_sc_hd__inv_2
X_2555_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ _0801_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
X_1506_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0819_ sky130_fd_sc_hd__inv_2
X_1437_ _0140_ vss vss vdd vdd _0495_ sky130_fd_sc_hd__clkbuf_1
X_2486_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out _0732_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
X_1368_ _0117_ vss vss vdd vdd _0470_ sky130_fd_sc_hd__clkbuf_1
X_2646__67 vss vss vdd vdd net67 _2646__67/LO sky130_fd_sc_hd__conb_1
X_1299_ _0091_ vss vss vdd vdd _0635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_287 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_192 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_257 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_107 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2340_ logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out _0586_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2271_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out _0517_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1153_ _0040_ vss vss vdd vdd _0863_ sky130_fd_sc_hd__clkbuf_1
X_1222_ _0065_ vss vss vdd vdd _0616_ sky130_fd_sc_hd__clkbuf_1
X_1084_ _0012_ vss vss vdd vdd _0016_ sky130_fd_sc_hd__clkbuf_1
X_1986_ clknet_4_9_0_prog_clk net160 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2607_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ _0853_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_0937_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2538_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out _0784_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_195 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2469_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out _0715_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_21_249 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1840_ net14 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out
+ sky130_fd_sc_hd__inv_2
X_1771_ _0258_ vss vss vdd vdd _0674_ sky130_fd_sc_hd__clkbuf_1
X_2254_ net20 _0500_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2323_ net30 _0569_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2185_ net22 _0431_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1205_ _0058_ vss vss vdd vdd _0868_ sky130_fd_sc_hd__clkbuf_1
X_1136_ _0033_ vss vss vdd vdd _0034_ sky130_fd_sc_hd__clkbuf_1
X_1067_ _0321_ vss vss vdd vdd _0760_ sky130_fd_sc_hd__buf_1
X_1969_ clknet_4_2_0_prog_clk net74 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_157 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold4 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd net71 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_219 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1823_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0275_ sky130_fd_sc_hd__clkbuf_1
X_1685_ _0230_ vss vss vdd vdd _0448_ sky130_fd_sc_hd__clkbuf_1
X_1754_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0253_ sky130_fd_sc_hd__clkbuf_1
X_2237_ net38 _0483_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_24_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2306_ net40 _0552_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_81 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2099_ net30 _0345_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1119_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd _0028_
+ sky130_fd_sc_hd__buf_6
X_2168_ net32 _0414_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_290 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_26_127 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_26_105 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1470_ _0152_ vss vss vdd vdd _0531_ sky130_fd_sc_hd__clkbuf_1
X_2022_ clknet_4_5_0_prog_clk net123 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1806_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd _0270_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_138 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_17_149 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_40_152 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1599_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q vss vss vdd vdd _0200_
+ sky130_fd_sc_hd__clkbuf_1
X_1668_ _0212_ vss vss vdd vdd _0397_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_260 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1737_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd _0248_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_130 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2640_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ _0886_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_0970_ _0288_ vss vss vdd vdd _0289_ sky130_fd_sc_hd__clkbuf_1
X_1522_ _0170_ vss vss vdd vdd _0796_ sky130_fd_sc_hd__clkbuf_1
X_2571_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ _0817_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_2
X_1453_ _0146_ vss vss vdd vdd _0147_ sky130_fd_sc_hd__clkbuf_1
X_2005_ clknet_4_13_0_prog_clk net78 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1384_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_61 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_42_93 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_12_0_prog_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_93 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_64 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_31 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_42 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_86 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_75 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_105 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_42_236 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2554_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ _0800_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_2623_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ _0869_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0953_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0334_ sky130_fd_sc_hd__inv_2
X_1505_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0820_ sky130_fd_sc_hd__inv_2
X_1367_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd _0117_
+ sky130_fd_sc_hd__clkbuf_1
X_1436_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd _0140_
+ sky130_fd_sc_hd__clkbuf_1
X_2343__56 vss vss vdd vdd net56 _2343__56/LO sky130_fd_sc_hd__conb_1
X_2485_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out _0731_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1298_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd _0091_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_222 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1221_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0065_
+ sky130_fd_sc_hd__clkbuf_1
X_2270_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out _0516_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1152_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0040_ sky130_fd_sc_hd__clkbuf_1
X_1083_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q vss vss vdd vdd _0742_
+ sky130_fd_sc_hd__inv_2
X_0936_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ vss vss vdd vdd _0890_ sky130_fd_sc_hd__inv_2
X_1985_ clknet_4_11_0_prog_clk net77 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2537_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out _0783_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2606_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ _0852_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_1419_ _0134_ vss vss vdd vdd _0506_ sky130_fd_sc_hd__clkbuf_1
X_2399_ net58 _0645_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2468_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out _0714_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_28_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1770_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q vss vss vdd vdd _0258_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_17 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_2184_ net25 _0430_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2253_ net28 _0499_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1204_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0058_ sky130_fd_sc_hd__clkbuf_1
X_2322_ net34 _0568_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1135_ _0033_ vss vss vdd vdd _0881_ sky130_fd_sc_hd__inv_2
X_1066_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q vss vss vdd vdd _0321_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_222 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_233 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1899_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__inv_2
X_1968_ clknet_4_1_0_prog_clk net178 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_261 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_39_28 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold5 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd net72 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1822_ _0028_ vss vss vdd vdd _0761_ sky130_fd_sc_hd__inv_2
X_1753_ _0162_ vss vss vdd vdd _0537_ sky130_fd_sc_hd__inv_2
X_1684_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0230_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_50 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2236_ net42 _0482_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2167_ net36 _0413_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_29_94 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2305_ net44 _0551_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2098_ net35 _0344_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1118_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0771_
+ sky130_fd_sc_hd__inv_2
X_1049_ _0307_ vss vss vdd vdd _0707_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_51 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_60 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_117 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_34_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2021_ clknet_4_5_0_prog_clk net88 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1805_ _0269_ vss vss vdd vdd _0783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_194 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1736_ _0247_ vss vss vdd vdd _0559_ sky130_fd_sc_hd__clkbuf_1
X_1598_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q vss vss vdd vdd _0382_
+ sky130_fd_sc_hd__inv_2
X_1667_ _0223_ vss vss vdd vdd _0411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2219_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out _0465_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_39_242 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2570_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ _0816_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_39_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1521_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0170_ sky130_fd_sc_hd__clkbuf_1
X_1383_ _0110_ vss vss vdd vdd _0453_ sky130_fd_sc_hd__inv_2
X_1452_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd _0146_
+ sky130_fd_sc_hd__buf_6
X_2004_ clknet_4_15_0_prog_clk net72 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_40 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_45_267 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1719_ _0162_ vss vss vdd vdd _0543_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_87 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_76 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_65 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_54 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_32 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_43 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_0952_ _0281_ vss vss vdd vdd _0906_ sky130_fd_sc_hd__clkbuf_1
X_2553_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ _0799_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_1504_ _0164_ vss vss vdd vdd _0789_ sky130_fd_sc_hd__clkbuf_1
X_2622_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ _0868_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_1366_ _0116_ vss vss vdd vdd _0475_ sky130_fd_sc_hd__clkbuf_1
X_1435_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0488_
+ sky130_fd_sc_hd__inv_2
X_2484_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out _0730_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1297_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0628_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_5_172 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1151_ _0033_ vss vss vdd vdd _0878_ sky130_fd_sc_hd__inv_2
X_1220_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q vss vss vdd vdd _0605_
+ sky130_fd_sc_hd__inv_2
X_1082_ _0012_ vss vss vdd vdd _0738_ sky130_fd_sc_hd__inv_2
X_0935_ net7 vss vss vdd vdd _0000_ sky130_fd_sc_hd__inv_2
X_1984_ clknet_4_9_0_prog_clk net181 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_237 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_63 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_74 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2605_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ _0851_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_2536_ logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out _0782_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2467_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out _0713_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_23_270 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1349_ _0110_ vss vss vdd vdd _0111_ sky130_fd_sc_hd__clkbuf_1
X_1418_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q vss vss vdd vdd _0134_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_73 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2398_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out _0644_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_28_19 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_2321_ net38 _0567_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2183_ net30 _0429_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2252_ net32 _0498_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1203_ _0057_ vss vss vdd vdd _0862_ sky130_fd_sc_hd__clkbuf_1
X_1134_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0033_ sky130_fd_sc_hd__buf_6
X_1065_ _0320_ vss vss vdd vdd _0894_ sky130_fd_sc_hd__clkbuf_1
X_1898_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__inv_2
X_1967_ clknet_4_1_0_prog_clk net201 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2519_ net31 _0765_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold6 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ vss vss vdd vdd net73 sky130_fd_sc_hd__dlygate4sd3_1
X_1683_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q vss vss vdd vdd _0437_
+ sky130_fd_sc_hd__inv_2
X_1821_ _0274_ vss vss vdd vdd _0775_ sky130_fd_sc_hd__clkbuf_1
X_1752_ _0252_ vss vss vdd vdd _0551_ sky130_fd_sc_hd__clkbuf_1
X_2304_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out _0550_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2097_ net39 _0343_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2235_ net46 _0481_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2166_ net40 _0412_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1117_ _0027_ vss vss vdd vdd _0785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1048_ _0315_ vss vss vdd vdd _0721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_281 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_34_184 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2020_ clknet_4_5_0_prog_clk net93 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_107 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_17_129 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1804_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0269_
+ sky130_fd_sc_hd__clkbuf_1
X_1666_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd _0223_
+ sky130_fd_sc_hd__clkbuf_1
X_1735_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0247_
+ sky130_fd_sc_hd__clkbuf_1
X_1597_ _0195_ vss vss vdd vdd _0373_ sky130_fd_sc_hd__inv_2
X_2149_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out _0395_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2218_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out _0464_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_31_165 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1520_ _0165_ vss vss vdd vdd _0811_ sky130_fd_sc_hd__inv_2
X_1382_ _0121_ vss vss vdd vdd _0467_ sky130_fd_sc_hd__clkbuf_1
X_1451_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0519_
+ sky130_fd_sc_hd__inv_2
X_2003_ clknet_4_13_0_prog_clk net125 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1718_ _0241_ vss vss vdd vdd _0790_ sky130_fd_sc_hd__buf_1
X_1649_ _0217_ vss vss vdd vdd _0422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_121 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_88 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_77 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_66 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_55 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_33 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_44 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_42_205 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_27_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_76 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_0951_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0281_ sky130_fd_sc_hd__clkbuf_1
X_2552_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ _0798_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_1503_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0164_ sky130_fd_sc_hd__clkbuf_1
X_2621_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ _0867_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_2483_ net61 _0729_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1365_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0116_
+ sky130_fd_sc_hd__clkbuf_1
X_1434_ _0129_ vss vss vdd vdd _0482_ sky130_fd_sc_hd__inv_2
X_1296_ _0080_ vss vss vdd vdd _0622_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_213 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_190 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _0039_ vss vss vdd vdd _0869_ sky130_fd_sc_hd__clkbuf_1
X_1081_ _0015_ vss vss vdd vdd _0752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_42 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2604_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ _0850_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
X_0934_ _0009_ net11 vss vss vdd vdd _0001_ sky130_fd_sc_hd__nand2_1
X_1983_ clknet_4_9_0_prog_clk net185 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_249 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2535_ net27 _0781_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1417_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q vss vss vdd vdd _0494_
+ sky130_fd_sc_hd__inv_2
X_2466_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out _0712_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1348_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd _0110_
+ sky130_fd_sc_hd__buf_6
X_1279_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q vss vss vdd vdd _0634_
+ sky130_fd_sc_hd__inv_2
X_2397_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out _0643_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2251_ net36 _0497_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2320_ net42 _0566_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2182_ net34 _0428_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1133_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0885_ sky130_fd_sc_hd__inv_2
X_1202_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0057_ sky130_fd_sc_hd__clkbuf_1
X_1064_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0320_ sky130_fd_sc_hd__clkbuf_1
X_1966_ clknet_4_1_0_prog_clk net169 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1897_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__inv_2
X_2518_ net35 _0764_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_252 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2449_ net29 _0695_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold7 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q vss vss vdd vdd net74
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1820_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q vss vss vdd vdd _0274_
+ sky130_fd_sc_hd__clkbuf_1
X_1682_ _0228_ vss vss vdd vdd _0431_ sky130_fd_sc_hd__inv_2
X_1751_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q vss vss vdd vdd _0252_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_32 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2234_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out _0480_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
X_2303_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out _0549_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1116_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q vss vss vdd vdd _0027_
+ sky130_fd_sc_hd__clkbuf_1
X_2096_ net42 _0342_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2165_ net45 _0411_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_9_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1047_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd _0315_
+ sky130_fd_sc_hd__clkbuf_1
X_1949_ clknet_4_5_0_prog_clk net203 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_141 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_1803_ _0268_ vss vss vdd vdd _0786_ sky130_fd_sc_hd__clkbuf_1
X_1596_ _0199_ vss vss vdd vdd _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_166 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1665_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0404_
+ sky130_fd_sc_hd__inv_2
X_1734_ _0246_ vss vss vdd vdd _0562_ sky130_fd_sc_hd__clkbuf_1
X_2217_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out _0463_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_22_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2148_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out _0394_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2079_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
+ _0325_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_130 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_16_152 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_16_163 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_39_233 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1450_ _0145_ vss vss vdd vdd _0533_ sky130_fd_sc_hd__clkbuf_1
X_1381_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q vss vss vdd vdd _0121_
+ sky130_fd_sc_hd__clkbuf_1
X_2002_ clknet_4_13_0_prog_clk net87 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1579_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q vss vss vdd vdd _0193_
+ sky130_fd_sc_hd__clkbuf_1
X_1648_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q vss vss vdd vdd _0217_
+ sky130_fd_sc_hd__clkbuf_1
X_1717_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ vss vss vdd vdd _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_89 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_78 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_67 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_56 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_160 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_34 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_45 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_182 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_258 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_236 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_27_225 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_2620_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ _0866_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_0950_ _0280_ vss vss vdd vdd _0899_ sky130_fd_sc_hd__clkbuf_1
X_2551_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ _0797_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_1502_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd _0340_ sky130_fd_sc_hd__inv_2
X_1433_ _0139_ vss vss vdd vdd _0496_ sky130_fd_sc_hd__clkbuf_1
X_2482_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out _0728_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1364_ _0115_ vss vss vdd vdd _0478_ sky130_fd_sc_hd__clkbuf_1
X_1295_ _0090_ vss vss vdd vdd _0636_ sky130_fd_sc_hd__clkbuf_1
XTAP_180 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_11_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_1080_ _0012_ vss vss vdd vdd _0015_ sky130_fd_sc_hd__clkbuf_1
X_1982_ clknet_4_8_0_prog_clk net163 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2534_ net21 _0780_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2603_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
+ _0849_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_0933_ net7 vss vss vdd vdd _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_228 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_250 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1347_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0463_
+ sky130_fd_sc_hd__inv_2
X_1416_ _0129_ vss vss vdd vdd _0485_ sky130_fd_sc_hd__inv_2
X_2396_ logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out _0642_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2465_ net22 _0711_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1278_ _0080_ vss vss vdd vdd _0625_ sky130_fd_sc_hd__inv_2
X_2250_ net40 _0496_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1201_ _0033_ vss vss vdd vdd _0877_ sky130_fd_sc_hd__inv_2
X_2181_ net38 _0427_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1132_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0887_ sky130_fd_sc_hd__inv_2
X_1063_ _0277_ vss vss vdd vdd _0325_ sky130_fd_sc_hd__inv_2
X_1965_ clknet_4_1_0_prog_clk net206 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2517_ net39 _0763_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1896_ net24 vss vss vdd vdd net15 sky130_fd_sc_hd__inv_2
X_2448_ net33 _0694_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2379_ net30 _0625_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold8 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd net75 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q vss vss vdd vdd _0544_
+ sky130_fd_sc_hd__inv_2
X_1681_ _0229_ vss vss vdd vdd _0445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_66 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2233_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out _0479_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2164_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out _0410_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_2302_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out _0548_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2095_ net47 _0341_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1115_ _0026_ vss vss vdd vdd _0787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_65 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1046_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0713_
+ sky130_fd_sc_hd__inv_2
X_1948_ clknet_4_12_0_prog_clk net170 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1879_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_9_52 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2612__66 vss vss vdd vdd net66 _2612__66/LO sky130_fd_sc_hd__conb_1
XFILLER_0_43_197 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_34_164 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_31_98 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1802_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q vss vss vdd vdd _0268_
+ sky130_fd_sc_hd__clkbuf_1
X_1733_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q vss vss vdd vdd _0246_
+ sky130_fd_sc_hd__clkbuf_1
X_1595_ _0195_ vss vss vdd vdd _0199_ sky130_fd_sc_hd__clkbuf_1
X_1664_ _0212_ vss vss vdd vdd _0398_ sky130_fd_sc_hd__inv_2
X_2147_ net49 _0393_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2216_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out _0462_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2078_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
+ _0324_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1029_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0309_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_175 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_6 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1380_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0460_
+ sky130_fd_sc_hd__inv_2
X_2001_ clknet_4_13_0_prog_clk net89 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_106 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1716_ _0240_ vss vss vdd vdd _0791_ sky130_fd_sc_hd__clkbuf_1
X_1578_ _0192_ vss vss vdd vdd _0396_ sky130_fd_sc_hd__buf_1
X_1647_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q vss vss vdd vdd _0410_
+ sky130_fd_sc_hd__inv_2
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_46 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_79 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_68 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_57 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_150 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2550_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ _0796_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_35_281 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_248 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1363_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q vss vss vdd vdd _0115_
+ sky130_fd_sc_hd__clkbuf_1
X_1501_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ vss vss vdd vdd _0339_ sky130_fd_sc_hd__inv_2
X_1432_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q vss vss vdd vdd _0139_
+ sky130_fd_sc_hd__clkbuf_1
X_2481_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out _0727_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1294_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q vss vss vdd vdd _0090_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_284 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_170 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0009_ net11 vss vss vdd vdd _0004_ sky130_fd_sc_hd__nand2_1
X_1981_ clknet_4_9_0_prog_clk net154 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_99 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2533_ net29 _0779_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2602_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
+ _0848_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_1346_ _0109_ vss vss vdd vdd _0477_ sky130_fd_sc_hd__clkbuf_1
X_1415_ _0133_ vss vss vdd vdd _0499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_43 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_10 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2395_ net26 _0641_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2464_ net25 _0710_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1277_ _0084_ vss vss vdd vdd _0639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2180_ net42 _0426_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1200_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0883_ sky130_fd_sc_hd__inv_2
X_1062_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0332_ sky130_fd_sc_hd__inv_2
X_1131_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0888_ sky130_fd_sc_hd__inv_2
X_1895_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ sky130_fd_sc_hd__inv_2
X_1964_ clknet_4_6_0_prog_clk net159 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2516_ net43 _0762_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2447_ net37 _0693_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1329_ _0102_ vss vss vdd vdd _0831_ sky130_fd_sc_hd__clkbuf_1
X_2378_ net34 _0624_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_184 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold9 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q vss vss vdd vdd net76
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_107 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_184 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_29_129 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1680_ _0228_ vss vss vdd vdd _0229_ sky130_fd_sc_hd__clkbuf_1
X_2301_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out _0547_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2232_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out _0478_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2163_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out _0409_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1114_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q vss vss vdd vdd _0026_
+ sky130_fd_sc_hd__clkbuf_1
X_2094_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ _0340_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1045_ _0307_ vss vss vdd vdd _0708_ sky130_fd_sc_hd__inv_2
X_1878_ net20 vss vss vdd vdd net17 sky130_fd_sc_hd__inv_2
XFILLER_0_43_187 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1947_ clknet_4_12_0_prog_clk net192 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_195 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_184 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_31_66 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_31_33 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_25_198 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1663_ _0222_ vss vss vdd vdd _0412_ sky130_fd_sc_hd__clkbuf_1
X_1801_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q vss vss vdd vdd _0774_
+ sky130_fd_sc_hd__inv_2
X_1732_ logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q vss vss vdd vdd _0550_
+ sky130_fd_sc_hd__inv_2
X_1594_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q vss vss vdd vdd _0378_
+ sky130_fd_sc_hd__inv_2
X_2146_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out _0392_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2215_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out _0461_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1028_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q vss vss vdd vdd _0717_
+ sky130_fd_sc_hd__inv_2
X_2203__51 vss vss vdd vdd net51 _2203__51/LO sky130_fd_sc_hd__conb_1
XFILLER_0_31_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2000_ clknet_4_14_0_prog_clk net172 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_88 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1715_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0240_ sky130_fd_sc_hd__clkbuf_1
X_1646_ _0212_ vss vss vdd vdd _0401_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_330 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q vss vss vdd vdd _0192_
+ sky130_fd_sc_hd__clkbuf_1
X_2129_ net23 _0375_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_69 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_58 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_47 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_27_205 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1500_ _0163_ vss vss vdd vdd _0557_ sky130_fd_sc_hd__clkbuf_1
X_2480_ logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out _0726_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_116 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1362_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q vss vss vdd vdd _0466_
+ sky130_fd_sc_hd__inv_2
X_1431_ _0138_ vss vss vdd vdd _0502_ sky130_fd_sc_hd__clkbuf_1
X_1293_ _0089_ vss vss vdd vdd _0642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1629_ _0210_ vss vss vdd vdd _0423_ sky130_fd_sc_hd__clkbuf_1
XTAP_160 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ clknet_4_2_0_prog_clk net158 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_0931_ net7 vss vss vdd vdd _0006_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_67 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2601_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ _0847_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ sky130_fd_sc_hd__ebufn_1
X_2532_ net33 _0778_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2463_ net31 _0709_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1345_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q vss vss vdd vdd _0109_
+ sky130_fd_sc_hd__clkbuf_1
X_1414_ _0129_ vss vss vdd vdd _0133_ sky130_fd_sc_hd__clkbuf_1
X_1276_ _0080_ vss vss vdd vdd _0084_ sky130_fd_sc_hd__clkbuf_1
X_2394_ net21 _0640_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1130_ _0032_ vss vss vdd vdd _0857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_277 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1061_ _0319_ vss vss vdd vdd _0905_ sky130_fd_sc_hd__clkbuf_1
X_1894_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ sky130_fd_sc_hd__inv_2
X_1963_ clknet_4_3_0_prog_clk net196 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2515_ net47 _0761_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2446_ net41 _0692_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_222 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1328_ _0099_ vss vss vdd vdd _0102_ sky130_fd_sc_hd__clkbuf_1
X_1259_ _0077_ vss vss vdd vdd _0648_ sky130_fd_sc_hd__buf_1
X_2377_ net38 _0623_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_46_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_4_219 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2231_ net52 _0477_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2300_ logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out _0546_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_65 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2093_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
+ _0339_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_8
X_2162_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out _0408_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_1113_ _0025_ vss vss vdd vdd _0788_ sky130_fd_sc_hd__buf_1
X_1044_ _0314_ vss vss vdd vdd _0722_ sky130_fd_sc_hd__clkbuf_1
X_1877_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ sky130_fd_sc_hd__inv_2
X_1946_ clknet_4_6_0_prog_clk net183 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_2429_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out _0675_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_19_163 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1800_ _0028_ vss vss vdd vdd _0765_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_136 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1662_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q vss vss vdd vdd _0222_
+ sky130_fd_sc_hd__clkbuf_1
X_1731_ _0162_ vss vss vdd vdd _0541_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_188 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_0_200 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1593_ _0195_ vss vss vdd vdd _0374_ sky130_fd_sc_hd__inv_2
X_2214_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out _0460_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_222 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2145_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out _0391_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1027_ _0307_ vss vss vdd vdd _0711_ sky130_fd_sc_hd__inv_2
X_1929_ clknet_4_11_0_prog_clk net85 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_122 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_8_0_prog_clk sky130_fd_sc_hd__clkbuf_8
Xhold90 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ vss vss vdd vdd net157 sky130_fd_sc_hd__dlygate4sd3_1
X_1576_ _0191_ vss vss vdd vdd _0793_ sky130_fd_sc_hd__clkbuf_1
X_1714_ _0228_ vss vss vdd vdd _0425_ sky130_fd_sc_hd__inv_2
X_1645_ _0216_ vss vss vdd vdd _0415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_169 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_331 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ net24 _0374_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_59 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_48 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_37 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_44_272 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_44_250 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1430_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0138_
+ sky130_fd_sc_hd__clkbuf_1
X_1361_ _0110_ vss vss vdd vdd _0457_ sky130_fd_sc_hd__inv_2
X_1292_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0089_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_239 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1559_ _0185_ vss vss vdd vdd _0362_ sky130_fd_sc_hd__clkbuf_1
X_1628_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q vss vss vdd vdd _0210_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_150 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2600_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ _0846_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ sky130_fd_sc_hd__ebufn_1
X_0930_ _0009_ net11 vss vss vdd vdd _0007_ sky130_fd_sc_hd__nand2_1
X_2531_ net37 _0777_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1413_ logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q vss vss vdd vdd _0490_
+ sky130_fd_sc_hd__inv_2
X_2462_ net34 _0708_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2393_ net28 _0639_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1344_ _0108_ vss vss vdd vdd _0479_ sky130_fd_sc_hd__clkbuf_1
X_1275_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q vss vss vdd vdd _0630_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_90 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_212 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1060_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1962_ clknet_4_3_0_prog_clk net166 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1893_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ sky130_fd_sc_hd__inv_2
X_2376_ net43 _0622_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2445_ net44 _0691_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2514_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out _0760_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ sky130_fd_sc_hd__ebufn_8
X_1327_ _0099_ vss vss vdd vdd _0846_ sky130_fd_sc_hd__inv_2
X_1258_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q vss vss vdd vdd _0077_
+ sky130_fd_sc_hd__clkbuf_1
X_1189_ _0053_ vss vss vdd vdd _0586_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_10_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_2230_ logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out _0476_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_29_45 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2161_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out _0407_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1112_ logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q vss vss vdd vdd _0025_
+ sky130_fd_sc_hd__clkbuf_1
X_2092_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ _0338_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ sky130_fd_sc_hd__ebufn_2
X_1043_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd _0314_
+ sky130_fd_sc_hd__clkbuf_1
X_1945_ clknet_4_6_0_prog_clk net149 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_178 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1876_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_3_297 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2428_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out _0674_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_2359_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out _0605_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1592_ _0198_ vss vss vdd vdd _0388_ sky130_fd_sc_hd__clkbuf_1
X_1661_ _0221_ vss vss vdd vdd _0418_ sky130_fd_sc_hd__clkbuf_1
X_1730_ _0245_ vss vss vdd vdd _0555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_178 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2213_ net22 _0459_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2144_ logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out _0390_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_289 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_256 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_267 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1026_ _0308_ vss vss vdd vdd _0725_ sky130_fd_sc_hd__clkbuf_1
X_1859_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ sky130_fd_sc_hd__inv_2
X_1928_ clknet_4_10_0_prog_clk net69 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_189 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold91 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q vss vss vdd vdd net158
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q vss vss vdd vdd net147
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ _0239_ vss vss vdd vdd _0439_ sky130_fd_sc_hd__clkbuf_1
XTAP_332 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0191_ sky130_fd_sc_hd__clkbuf_1
XTAP_321 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1644_ _0212_ vss vss vdd vdd _0216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_148 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2127_ net31 _0373_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_49 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1009_ _0277_ vss vss vdd vdd _0327_ sky130_fd_sc_hd__inv_2
XPHY_38 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_44_240 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_35_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1360_ _0114_ vss vss vdd vdd _0471_ sky130_fd_sc_hd__clkbuf_1
X_1291_ logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q vss vss vdd vdd _0632_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_41_276 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_284 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1558_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0185_
+ sky130_fd_sc_hd__clkbuf_1
X_1627_ _0209_ vss vss vdd vdd _0424_ sky130_fd_sc_hd__buf_1
XTAP_140 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _0158_ vss vss vdd vdd _0833_ sky130_fd_sc_hd__clkbuf_1
XTAP_195 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_251 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2530_ net41 _0776_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1343_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q vss vss vdd vdd _0108_
+ sky130_fd_sc_hd__clkbuf_1
X_1412_ _0129_ vss vss vdd vdd _0486_ sky130_fd_sc_hd__inv_2
X_2461_ net39 _0707_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2392_ net32 _0638_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1274_ _0080_ vss vss vdd vdd _0626_ sky130_fd_sc_hd__inv_2
X_0989_ _0295_ vss vss vdd vdd _0694_ sky130_fd_sc_hd__clkbuf_1
X_2659_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ _0905_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_14_243 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_14_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_69 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1892_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ sky130_fd_sc_hd__inv_2
X_1961_ clknet_4_3_0_prog_clk net148 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_2513_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out _0759_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1326_ _0101_ vss vss vdd vdd _0836_ sky130_fd_sc_hd__clkbuf_1
X_2375_ net46 _0621_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2444_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out _0690_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_11_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1257_ _0076_ vss vss vdd vdd _0860_ sky130_fd_sc_hd__clkbuf_1
X_1188_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q vss vss vdd vdd _0053_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2160_ logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out _0406_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1111_ _0277_ vss vss vdd vdd _0324_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_47 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2091_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ _0337_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
+ sky130_fd_sc_hd__ebufn_1
X_1042_ _0313_ vss vss vdd vdd _0727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_113 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_43_102 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1944_ clknet_4_15_0_prog_clk net174 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1875_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_132 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2427_ net59 _0673_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1309_ _0095_ vss vss vdd vdd _0673_ sky130_fd_sc_hd__clkbuf_1
X_2358_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out _0604_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2289_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out _0535_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_25_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1591_ _0195_ vss vss vdd vdd _0198_ sky130_fd_sc_hd__clkbuf_1
X_1660_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0221_
+ sky130_fd_sc_hd__clkbuf_1
X_2143_ net27 _0389_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2212_ net25 _0458_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1025_ _0307_ vss vss vdd vdd _0308_ sky130_fd_sc_hd__clkbuf_1
X_1858_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
+ sky130_fd_sc_hd__inv_2
X_1927_ clknet_4_10_0_prog_clk net127 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1789_ _0264_ vss vss vdd vdd _0663_ sky130_fd_sc_hd__clkbuf_1
Xhold70 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q vss vss vdd vdd net148
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q vss vss vdd vdd net159
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1712_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q vss vss vdd vdd _0239_
+ sky130_fd_sc_hd__clkbuf_1
X_1643_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q vss vss vdd vdd _0406_
+ sky130_fd_sc_hd__inv_2
XANTENNA_1 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
+ vss vss vdd vdd sky130_fd_sc_hd__diode_2
XTAP_333 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _0165_ vss vss vdd vdd _0808_ sky130_fd_sc_hd__inv_2
XTAP_311 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2126_ net35 _0372_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2057_ clknet_4_8_0_prog_clk net204 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_28 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1008_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0333_ sky130_fd_sc_hd__inv_2
XPHY_39 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_44_263 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1290_ _0080_ vss vss vdd vdd _0623_ sky130_fd_sc_hd__inv_2
X_1626_ logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q vss vss vdd vdd _0209_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1557_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q vss vss vdd vdd _0352_
+ sky130_fd_sc_hd__inv_2
X_1488_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0158_ sky130_fd_sc_hd__clkbuf_1
XTAP_130 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ net45 _0355_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_241 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_23_48 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2460_ net43 _0706_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1342_ _0107_ vss vss vdd vdd _0480_ sky130_fd_sc_hd__clkbuf_1
X_1411_ _0132_ vss vss vdd vdd _0500_ sky130_fd_sc_hd__clkbuf_1
X_2391_ net36 _0637_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1273_ _0083_ vss vss vdd vdd _0640_ sky130_fd_sc_hd__clkbuf_1
X_0988_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd _0295_
+ sky130_fd_sc_hd__clkbuf_1
X_1609_ _0195_ vss vss vdd vdd _0371_ sky130_fd_sc_hd__inv_2
X_2589_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ _0835_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
X_2658_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
+ _0904_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_1960_ clknet_4_6_0_prog_clk net190 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1891_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_11_236 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2443_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out _0689_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_4
X_2512_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out _0758_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1325_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0101_ sky130_fd_sc_hd__clkbuf_1
X_1256_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0076_ sky130_fd_sc_hd__clkbuf_1
X_2374_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out _0620_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_0_46_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1187_ logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q vss vss vdd vdd _0576_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_40_90 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_166 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_37_122 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_2090_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ _0336_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
+ sky130_fd_sc_hd__ebufn_1
X_1110_ _0024_ vss vss vdd vdd _0901_ sky130_fd_sc_hd__clkbuf_1
X_1041_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0313_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_147 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1874_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ sky130_fd_sc_hd__inv_2
X_1943_ clknet_4_15_0_prog_clk net182 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_35 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2426_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out _0672_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1308_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0095_
+ sky130_fd_sc_hd__clkbuf_1
X_1239_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q vss vss vdd vdd _0071_
+ sky130_fd_sc_hd__clkbuf_1
X_2357_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out _0603_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2288_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out _0534_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_155 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_177 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2119__48 vss vss vdd vdd net48 _2119__48/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_169 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_136 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1590_ _0197_ vss vss vdd vdd _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_180 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_2211_ net30 _0457_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2142_ net20 _0388_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1024_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q vss vss vdd vdd _0307_
+ sky130_fd_sc_hd__buf_6
XFILLER_0_16_103 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1857_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
+ sky130_fd_sc_hd__inv_2
X_1788_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q vss vss vdd vdd _0264_
+ sky130_fd_sc_hd__clkbuf_1
X_1926_ clknet_4_10_0_prog_clk net98 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
+ sky130_fd_sc_hd__dfxtp_1
X_2409_ net23 _0655_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_30_194 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_22_117 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold82 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q vss vss vdd vdd net149
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ vss vss vdd vdd net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_48 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold60 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
+ vss vss vdd vdd net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd net160
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1711_ logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q vss vss vdd vdd _0432_
+ sky130_fd_sc_hd__inv_2
X_1642_ _0212_ vss vss vdd vdd _0402_ sky130_fd_sc_hd__inv_2
XANTENNA_2 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
+ vss vss vdd vdd sky130_fd_sc_hd__diode_2
XFILLER_0_13_128 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_334 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _0190_ vss vss vdd vdd _0800_ sky130_fd_sc_hd__clkbuf_1
XTAP_301 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ net39 _0371_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2056_ clknet_4_8_0_prog_clk net134 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_1007_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
+ vss vss vdd vdd _0336_ sky130_fd_sc_hd__inv_2
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_44_220 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_100 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1909_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_35_242 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_253 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_18_209 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_41_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1625_ _0208_ vss vss vdd vdd _0792_ sky130_fd_sc_hd__clkbuf_1
X_1556_ _0184_ vss vss vdd vdd _0357_ sky130_fd_sc_hd__clkbuf_1
XTAP_120 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _0146_ vss vss vdd vdd _0509_ sky130_fd_sc_hd__inv_2
XTAP_197 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out _0354_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_4_7_0_prog_clk sky130_fd_sc_hd__clkbuf_8
X_2039_ clknet_4_0_0_prog_clk net96 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1410_ _0129_ vss vss vdd vdd _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_128 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1341_ logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q vss vss vdd vdd _0107_
+ sky130_fd_sc_hd__clkbuf_1
X_2390_ net41 _0636_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1272_ _0080_ vss vss vdd vdd _0083_ sky130_fd_sc_hd__clkbuf_1
X_0987_ _0294_ vss vss vdd vdd _0699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1539_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q vss vss vdd vdd _0353_
+ sky130_fd_sc_hd__inv_2
X_1608_ _0203_ vss vss vdd vdd _0385_ sky130_fd_sc_hd__clkbuf_1
X_2588_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ _0834_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_2657_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
+ _0903_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_34_59 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1890_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ sky130_fd_sc_hd__inv_2
X_2442_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out _0688_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2373_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out _0619_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2511_ net62 _0757_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_45_8 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_1324_ _0100_ vss vss vdd vdd _0832_ sky130_fd_sc_hd__clkbuf_1
X_1255_ _0033_ vss vss vdd vdd _0875_ sky130_fd_sc_hd__inv_2
X_1186_ _0044_ vss vss vdd vdd _0567_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_156 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_92 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_292 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1040_ _0312_ vss vss vdd vdd _0730_ sky130_fd_sc_hd__clkbuf_1
X_1942_ clknet_4_13_0_prog_clk net152 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_1873_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_3_223 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2425_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out _0671_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2356_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out _0602_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1307_ _0094_ vss vss vdd vdd _0675_ sky130_fd_sc_hd__clkbuf_1
X_1238_ logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q vss vss vdd vdd _0601_
+ sky130_fd_sc_hd__inv_2
X_1169_ _0047_ vss vss vdd vdd _0584_ sky130_fd_sc_hd__clkbuf_1
X_2287_ net54 _0533_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_19_167 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_104 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2210_ net34 _0456_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2141_ net29 _0387_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1023_ logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q vss vss vdd vdd _0715_
+ sky130_fd_sc_hd__inv_2
X_1925_ clknet_4_10_0_prog_clk net111 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1856_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
+ sky130_fd_sc_hd__inv_2
X_1787_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q vss vss vdd vdd _0656_
+ sky130_fd_sc_hd__inv_2
X_2339_ net26 _0585_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2408_ net24 _0654_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_92 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold61 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
+ vss vss vdd vdd net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q vss vss vdd vdd net139
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q vss vss vdd vdd net150
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
+ vss vss vdd vdd net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q vss vss vdd vdd net161
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_251 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1572_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0190_ sky130_fd_sc_hd__clkbuf_1
X_1710_ _0228_ vss vss vdd vdd _0426_ sky130_fd_sc_hd__inv_2
X_1641_ _0215_ vss vss vdd vdd _0416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_37 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XANTENNA_3 right_width_0_height_0_subtile_0__pin_I_5_ vss vss vdd vdd sky130_fd_sc_hd__diode_2
XTAP_335 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ net42 _0370_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1006_ _0300_ vss vss vdd vdd _0907_ sky130_fd_sc_hd__clkbuf_1
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_2055_ _0011_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
+ _0009_ _0010_ vss vss vdd vdd _2055_/Q logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
+ sky130_fd_sc_hd__dfbbn_1
XFILLER_0_44_276 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1839_ net6 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out
+ sky130_fd_sc_hd__inv_2
X_1908_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ sky130_fd_sc_hd__inv_2
XFILLER_0_12_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1624_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
+ vss vss vdd vdd _0208_ sky130_fd_sc_hd__clkbuf_1
X_1555_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q vss vss vdd vdd _0184_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_121 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out _0353_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_143 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _0157_ vss vss vdd vdd _0523_ sky130_fd_sc_hd__clkbuf_1
XTAP_198 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2038_ clknet_4_1_0_prog_clk net137 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_268 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_298 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_202 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1340_ _0106_ vss vss vdd vdd _0829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_1271_ _0082_ vss vss vdd vdd _0644_ sky130_fd_sc_hd__clkbuf_1
X_2656_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
+ _0902_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
+ sky130_fd_sc_hd__ebufn_1
X_0986_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q vss vss vdd vdd _0294_
+ sky130_fd_sc_hd__clkbuf_1
X_1538_ _0176_ vss vss vdd vdd _0347_ sky130_fd_sc_hd__inv_2
X_1607_ logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q vss vss vdd vdd _0203_
+ sky130_fd_sc_hd__clkbuf_1
X_1469_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q vss vss vdd vdd _0152_
+ sky130_fd_sc_hd__clkbuf_1
X_2587_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
+ _0833_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
+ sky130_fd_sc_hd__ebufn_1
X_2315__55 vss vss vdd vdd net55 _2315__55/LO sky130_fd_sc_hd__conb_1
XFILLER_0_9_284 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2539__63 vss vss vdd vdd net63 _2539__63/LO sky130_fd_sc_hd__conb_1
X_2510_ logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out _0756_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1323_ _0099_ vss vss vdd vdd _0100_ sky130_fd_sc_hd__clkbuf_1
X_2372_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out _0618_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2441_ logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out _0687_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1254_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
+ vss vss vdd vdd _0882_ sky130_fd_sc_hd__inv_2
X_1185_ _0052_ vss vss vdd vdd _0581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2639_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
+ _0885_ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
+ sky130_fd_sc_hd__ebufn_1
X_0969_ logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q vss vss vdd vdd _0288_
+ sky130_fd_sc_hd__buf_6
X_1872_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
+ sky130_fd_sc_hd__inv_2
X_1941_ clknet_4_12_0_prog_clk net139 vss vss vdd vdd logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_157 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_28_124 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_3_279 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_202 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_43_6 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2424_ logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out _0670_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1306_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q vss vss vdd vdd _0094_
+ sky130_fd_sc_hd__clkbuf_1
X_2355_ logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out _0601_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2286_ logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out _0532_
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1237_ _0063_ vss vss vdd vdd _0596_ sky130_fd_sc_hd__inv_2
X_1168_ _0044_ vss vss vdd vdd _0047_ sky130_fd_sc_hd__clkbuf_1
X_1099_ logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q vss vss vdd vdd _0744_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_42_171 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_190 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2140_ net33 _0386_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_1022_ _0306_ vss vss vdd vdd _0729_ sky130_fd_sc_hd__clkbuf_1
X_1855_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
+ sky130_fd_sc_hd__inv_2
X_1924_ clknet_4_10_0_prog_clk net119 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_24_182 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1786_ _0096_ vss vss vdd vdd _0650_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_2338_ net20 _0584_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2407_ net31 _0653_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_2269_ net23 _0515_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_30_163 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_30_152 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold40 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
+ vss vss vdd vdd net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ vss vss vdd vdd net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q vss vss vdd vdd net140
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
+ vss vss vdd vdd net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q vss vss vdd vdd net162
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q vss vss vdd vdd net129
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_285 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1571_ _0189_ vss vss vdd vdd _0794_ sky130_fd_sc_hd__clkbuf_1
XTAP_314 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _0212_ vss vss vdd vdd _0215_ sky130_fd_sc_hd__clkbuf_1
XTAP_336 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ net47 _0369_ vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_29_263 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_2054_ clknet_4_8_0_prog_clk net141 vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
+ sky130_fd_sc_hd__dfxtp_1
X_1005_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
+ vss vss vdd vdd _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_94 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_44_211 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_32_71 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_1838_ net2 vss vss vdd vdd logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out
+ sky130_fd_sc_hd__inv_2
X_1907_ logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
+ vss vss vdd vdd logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
+ sky130_fd_sc_hd__inv_2
X_1769_ logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q vss vss vdd vdd _0662_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_12_152 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_41_203 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_1623_ _0165_ vss vss vdd vdd _0807_ sky130_fd_sc_hd__inv_2
X_1554_ logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q vss vss vdd vdd _0349_
+ sky130_fd_sc_hd__inv_2
XTAP_122 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q vss vss vdd vdd _0157_
+ sky130_fd_sc_hd__clkbuf_1
.ends

