magic
tech sky130A
magscale 1 2
timestamp 1708041393
<< viali >>
rect 2421 21641 2455 21675
rect 3065 21641 3099 21675
rect 3341 21641 3375 21675
rect 4997 21641 5031 21675
rect 5917 21641 5951 21675
rect 7573 21641 7607 21675
rect 7849 21641 7883 21675
rect 8493 21641 8527 21675
rect 9321 21641 9355 21675
rect 10057 21641 10091 21675
rect 10793 21641 10827 21675
rect 11713 21641 11747 21675
rect 14105 21641 14139 21675
rect 2697 21573 2731 21607
rect 8401 21573 8435 21607
rect 11621 21573 11655 21607
rect 1685 21505 1719 21539
rect 1777 21505 1811 21539
rect 2145 21505 2179 21539
rect 2881 21505 2915 21539
rect 3157 21505 3191 21539
rect 3617 21505 3651 21539
rect 3801 21505 3835 21539
rect 4353 21505 4387 21539
rect 4629 21505 4663 21539
rect 4905 21505 4939 21539
rect 5181 21505 5215 21539
rect 5641 21505 5675 21539
rect 5733 21505 5767 21539
rect 6009 21505 6043 21539
rect 6377 21505 6411 21539
rect 7021 21505 7055 21539
rect 7113 21505 7147 21539
rect 7389 21505 7423 21539
rect 7757 21505 7791 21539
rect 9229 21505 9263 21539
rect 9965 21505 9999 21539
rect 10701 21505 10735 21539
rect 11345 21505 11379 21539
rect 12081 21505 12115 21539
rect 14289 21505 14323 21539
rect 4261 21437 4295 21471
rect 6929 21437 6963 21471
rect 12449 21437 12483 21471
rect 12633 21437 12667 21471
rect 13185 21437 13219 21471
rect 3525 21369 3559 21403
rect 4537 21369 4571 21403
rect 6561 21369 6595 21403
rect 13093 21369 13127 21403
rect 1593 21301 1627 21335
rect 3985 21301 4019 21335
rect 4813 21301 4847 21335
rect 5365 21301 5399 21335
rect 5457 21301 5491 21335
rect 6101 21301 6135 21335
rect 7205 21301 7239 21335
rect 11253 21301 11287 21335
rect 12265 21301 12299 21335
rect 13829 21301 13863 21335
rect 1501 21097 1535 21131
rect 4997 21097 5031 21131
rect 7205 21097 7239 21131
rect 7941 21097 7975 21131
rect 8493 21097 8527 21131
rect 8769 21097 8803 21131
rect 3893 21029 3927 21063
rect 13829 21029 13863 21063
rect 3525 20961 3559 20995
rect 6745 20961 6779 20995
rect 8125 20961 8159 20995
rect 11897 20961 11931 20995
rect 13277 20961 13311 20995
rect 2513 20893 2547 20927
rect 2697 20893 2731 20927
rect 2973 20893 3007 20927
rect 4077 20893 4111 20927
rect 4169 20893 4203 20927
rect 4905 20893 4939 20927
rect 5181 20893 5215 20927
rect 5825 20893 5859 20927
rect 6561 20893 6595 20927
rect 7297 20893 7331 20927
rect 7481 20893 7515 20927
rect 8217 20893 8251 20927
rect 8309 20893 8343 20927
rect 8585 20893 8619 20927
rect 8953 20893 8987 20927
rect 10609 20893 10643 20927
rect 11253 20893 11287 20927
rect 11713 20893 11747 20927
rect 11989 20893 12023 20927
rect 12173 20893 12207 20927
rect 12909 20893 12943 20927
rect 14289 20893 14323 20927
rect 1777 20825 1811 20859
rect 5549 20825 5583 20859
rect 5733 20825 5767 20859
rect 9198 20825 9232 20859
rect 13369 20825 13403 20859
rect 2053 20757 2087 20791
rect 2329 20757 2363 20791
rect 2881 20757 2915 20791
rect 4813 20757 4847 20791
rect 5365 20757 5399 20791
rect 6469 20757 6503 20791
rect 10333 20757 10367 20791
rect 11161 20757 11195 20791
rect 12633 20757 12667 20791
rect 12725 20757 12759 20791
rect 14105 20757 14139 20791
rect 2237 20553 2271 20587
rect 2329 20553 2363 20587
rect 3985 20553 4019 20587
rect 6193 20553 6227 20587
rect 10517 20553 10551 20587
rect 1777 20485 1811 20519
rect 4344 20485 4378 20519
rect 6622 20485 6656 20519
rect 13360 20485 13394 20519
rect 2053 20417 2087 20451
rect 2513 20417 2547 20451
rect 2605 20417 2639 20451
rect 2872 20417 2906 20451
rect 5733 20417 5767 20451
rect 7941 20417 7975 20451
rect 8861 20417 8895 20451
rect 9873 20417 9907 20451
rect 10609 20417 10643 20451
rect 11253 20417 11287 20451
rect 11529 20417 11563 20451
rect 11785 20417 11819 20451
rect 13093 20417 13127 20451
rect 4077 20349 4111 20383
rect 5549 20349 5583 20383
rect 6377 20349 6411 20383
rect 8125 20349 8159 20383
rect 8953 20349 8987 20383
rect 9597 20349 9631 20383
rect 9781 20349 9815 20383
rect 10057 20349 10091 20383
rect 1501 20213 1535 20247
rect 5457 20213 5491 20247
rect 7757 20213 7791 20247
rect 8585 20213 8619 20247
rect 9137 20213 9171 20247
rect 10793 20213 10827 20247
rect 11161 20213 11195 20247
rect 12909 20213 12943 20247
rect 14473 20213 14507 20247
rect 6285 20009 6319 20043
rect 8309 20009 8343 20043
rect 9965 20009 9999 20043
rect 10517 20009 10551 20043
rect 10885 20009 10919 20043
rect 11345 20009 11379 20043
rect 1777 19941 1811 19975
rect 3525 19941 3559 19975
rect 8677 19941 8711 19975
rect 3157 19873 3191 19907
rect 6653 19873 6687 19907
rect 9137 19873 9171 19907
rect 11529 19873 11563 19907
rect 12633 19873 12667 19907
rect 1685 19805 1719 19839
rect 3433 19805 3467 19839
rect 3985 19805 4019 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 6101 19805 6135 19839
rect 8401 19805 8435 19839
rect 8493 19805 8527 19839
rect 8953 19805 8987 19839
rect 10057 19805 10091 19839
rect 10333 19805 10367 19839
rect 10609 19805 10643 19839
rect 10701 19805 10735 19839
rect 11713 19805 11747 19839
rect 12173 19805 12207 19839
rect 12449 19805 12483 19839
rect 14105 19805 14139 19839
rect 2912 19737 2946 19771
rect 4261 19737 4295 19771
rect 4813 19737 4847 19771
rect 4905 19737 4939 19771
rect 5089 19737 5123 19771
rect 6920 19737 6954 19771
rect 11069 19737 11103 19771
rect 13093 19737 13127 19771
rect 13277 19737 13311 19771
rect 13369 19737 13403 19771
rect 13921 19737 13955 19771
rect 1593 19669 1627 19703
rect 4169 19669 4203 19703
rect 8033 19669 8067 19703
rect 9597 19669 9631 19703
rect 10149 19669 10183 19703
rect 14289 19669 14323 19703
rect 2513 19465 2547 19499
rect 4537 19465 4571 19499
rect 6101 19465 6135 19499
rect 7021 19465 7055 19499
rect 7205 19465 7239 19499
rect 7665 19465 7699 19499
rect 7941 19465 7975 19499
rect 9413 19465 9447 19499
rect 9689 19465 9723 19499
rect 12357 19465 12391 19499
rect 13277 19465 13311 19499
rect 14013 19465 14047 19499
rect 14197 19465 14231 19499
rect 3801 19397 3835 19431
rect 5273 19397 5307 19431
rect 8309 19397 8343 19431
rect 10517 19397 10551 19431
rect 1777 19329 1811 19363
rect 1961 19329 1995 19363
rect 2329 19329 2363 19363
rect 2605 19329 2639 19363
rect 2697 19329 2731 19363
rect 3065 19329 3099 19363
rect 5181 19329 5215 19363
rect 6009 19329 6043 19363
rect 7389 19329 7423 19363
rect 7481 19329 7515 19363
rect 7757 19329 7791 19363
rect 8033 19329 8067 19363
rect 8125 19329 8159 19363
rect 8953 19329 8987 19363
rect 9229 19329 9263 19363
rect 9505 19329 9539 19363
rect 10609 19329 10643 19363
rect 10977 19329 11011 19363
rect 11529 19329 11563 19363
rect 12449 19329 12483 19363
rect 12633 19329 12667 19363
rect 13369 19329 13403 19363
rect 14105 19329 14139 19363
rect 2881 19261 2915 19295
rect 3525 19261 3559 19295
rect 3709 19261 3743 19295
rect 4353 19261 4387 19295
rect 4997 19261 5031 19295
rect 5917 19261 5951 19295
rect 6377 19261 6411 19295
rect 8769 19261 8803 19295
rect 9873 19261 9907 19295
rect 10057 19261 10091 19295
rect 11713 19261 11747 19295
rect 12817 19261 12851 19295
rect 13553 19261 13587 19295
rect 11161 19193 11195 19227
rect 1501 19125 1535 19159
rect 2145 19125 2179 19159
rect 10701 19125 10735 19159
rect 12173 19125 12207 19159
rect 1593 18921 1627 18955
rect 3433 18921 3467 18955
rect 4169 18921 4203 18955
rect 4445 18921 4479 18955
rect 9689 18921 9723 18955
rect 10517 18921 10551 18955
rect 11621 18921 11655 18955
rect 12449 18921 12483 18955
rect 13001 18921 13035 18955
rect 13829 18921 13863 18955
rect 4629 18853 4663 18887
rect 4997 18853 5031 18887
rect 5273 18853 5307 18887
rect 7573 18853 7607 18887
rect 7941 18853 7975 18887
rect 8217 18853 8251 18887
rect 8493 18853 8527 18887
rect 2053 18785 2087 18819
rect 5549 18785 5583 18819
rect 6193 18785 6227 18819
rect 9229 18785 9263 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 1409 18717 1443 18751
rect 1869 18717 1903 18751
rect 2789 18717 2823 18751
rect 2973 18717 3007 18751
rect 3985 18717 4019 18751
rect 4261 18717 4295 18751
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 5089 18717 5123 18751
rect 5365 18717 5399 18751
rect 6929 18717 6963 18751
rect 7205 18717 7239 18751
rect 7481 18717 7515 18751
rect 7757 18717 7791 18751
rect 8033 18717 8067 18751
rect 8309 18717 8343 18751
rect 8585 18717 8619 18751
rect 8677 18717 8711 18751
rect 9045 18717 9079 18751
rect 9873 18717 9907 18751
rect 10425 18717 10459 18751
rect 10977 18717 11011 18751
rect 11161 18717 11195 18751
rect 11253 18717 11287 18751
rect 12173 18717 12207 18751
rect 13553 18717 13587 18751
rect 14105 18717 14139 18751
rect 6285 18649 6319 18683
rect 6837 18649 6871 18683
rect 12909 18649 12943 18683
rect 2513 18581 2547 18615
rect 6009 18581 6043 18615
rect 7113 18581 7147 18615
rect 7389 18581 7423 18615
rect 14289 18581 14323 18615
rect 2329 18377 2363 18411
rect 5089 18377 5123 18411
rect 5365 18377 5399 18411
rect 8769 18377 8803 18411
rect 11621 18377 11655 18411
rect 6469 18309 6503 18343
rect 6561 18309 6595 18343
rect 13921 18309 13955 18343
rect 14105 18309 14139 18343
rect 1409 18241 1443 18275
rect 1869 18241 1903 18275
rect 2605 18241 2639 18275
rect 3341 18241 3375 18275
rect 3689 18241 3723 18275
rect 4905 18241 4939 18275
rect 5273 18241 5307 18275
rect 6101 18241 6135 18275
rect 7389 18241 7423 18275
rect 8125 18241 8159 18275
rect 8401 18241 8435 18275
rect 8677 18241 8711 18275
rect 9137 18241 9171 18275
rect 9597 18241 9631 18275
rect 9965 18241 9999 18275
rect 11529 18241 11563 18275
rect 12173 18241 12207 18275
rect 12449 18241 12483 18275
rect 13553 18241 13587 18275
rect 1685 18173 1719 18207
rect 2421 18173 2455 18207
rect 3433 18173 3467 18207
rect 7205 18173 7239 18207
rect 10149 18173 10183 18207
rect 10701 18173 10735 18207
rect 10885 18173 10919 18207
rect 12725 18173 12759 18207
rect 12909 18173 12943 18207
rect 4813 18105 4847 18139
rect 7021 18105 7055 18139
rect 8217 18105 8251 18139
rect 9229 18105 9263 18139
rect 12265 18105 12299 18139
rect 1593 18037 1627 18071
rect 2789 18037 2823 18071
rect 3249 18037 3283 18071
rect 5549 18037 5583 18071
rect 7573 18037 7607 18071
rect 7941 18037 7975 18071
rect 9781 18037 9815 18071
rect 10609 18037 10643 18071
rect 11345 18037 11379 18071
rect 12081 18037 12115 18071
rect 13369 18037 13403 18071
rect 14381 18037 14415 18071
rect 2421 17833 2455 17867
rect 8585 17833 8619 17867
rect 9413 17833 9447 17867
rect 9965 17833 9999 17867
rect 10701 17833 10735 17867
rect 10885 17833 10919 17867
rect 12541 17833 12575 17867
rect 13001 17833 13035 17867
rect 13461 17833 13495 17867
rect 7113 17765 7147 17799
rect 9505 17765 9539 17799
rect 10517 17765 10551 17799
rect 11345 17765 11379 17799
rect 11437 17765 11471 17799
rect 2605 17697 2639 17731
rect 5181 17697 5215 17731
rect 7389 17697 7423 17731
rect 7941 17697 7975 17731
rect 12081 17697 12115 17731
rect 12817 17697 12851 17731
rect 1409 17629 1443 17663
rect 2789 17629 2823 17663
rect 3433 17629 3467 17663
rect 3893 17629 3927 17663
rect 4813 17629 4847 17663
rect 6929 17629 6963 17663
rect 7205 17629 7239 17663
rect 8125 17629 8159 17663
rect 8953 17629 8987 17663
rect 9229 17629 9263 17663
rect 9689 17629 9723 17663
rect 9781 17629 9815 17663
rect 10057 17629 10091 17663
rect 10333 17629 10367 17663
rect 10793 17629 10827 17663
rect 11069 17629 11103 17663
rect 11161 17629 11195 17663
rect 11621 17629 11655 17663
rect 11897 17629 11931 17663
rect 12633 17629 12667 17663
rect 13553 17629 13587 17663
rect 13645 17629 13679 17663
rect 14289 17629 14323 17663
rect 1777 17561 1811 17595
rect 5448 17561 5482 17595
rect 2881 17493 2915 17527
rect 3985 17493 4019 17527
rect 4261 17493 4295 17527
rect 6561 17493 6595 17527
rect 7849 17493 7883 17527
rect 9137 17493 9171 17527
rect 10241 17493 10275 17527
rect 13737 17493 13771 17527
rect 14105 17493 14139 17527
rect 1961 17289 1995 17323
rect 5733 17289 5767 17323
rect 6101 17289 6135 17323
rect 7573 17289 7607 17323
rect 8861 17289 8895 17323
rect 13369 17289 13403 17323
rect 4414 17221 4448 17255
rect 9873 17221 9907 17255
rect 10425 17221 10459 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2421 17153 2455 17187
rect 2697 17153 2731 17187
rect 2964 17153 2998 17187
rect 5917 17153 5951 17187
rect 6009 17153 6043 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 7021 17153 7055 17187
rect 7757 17153 7791 17187
rect 7941 17153 7975 17187
rect 9137 17153 9171 17187
rect 9505 17153 9539 17187
rect 9965 17153 9999 17187
rect 10057 17153 10091 17187
rect 10333 17153 10367 17187
rect 10609 17153 10643 17187
rect 11069 17153 11103 17187
rect 11161 17153 11195 17187
rect 11537 17153 11571 17187
rect 14197 17153 14231 17187
rect 4169 17085 4203 17119
rect 6837 17085 6871 17119
rect 8217 17085 8251 17119
rect 8401 17085 8435 17119
rect 11897 17085 11931 17119
rect 12081 17085 12115 17119
rect 12633 17085 12667 17119
rect 12817 17085 12851 17119
rect 13829 17085 13863 17119
rect 14013 17085 14047 17119
rect 5549 17017 5583 17051
rect 8125 17017 8159 17051
rect 8953 17017 8987 17051
rect 9597 17017 9631 17051
rect 10793 17017 10827 17051
rect 10885 17017 10919 17051
rect 12541 17017 12575 17051
rect 13001 17017 13035 17051
rect 1501 16949 1535 16983
rect 2237 16949 2271 16983
rect 4077 16949 4111 16983
rect 7205 16949 7239 16983
rect 10241 16949 10275 16983
rect 11253 16949 11287 16983
rect 11713 16949 11747 16983
rect 14381 16949 14415 16983
rect 12725 16745 12759 16779
rect 13369 16745 13403 16779
rect 5733 16677 5767 16711
rect 11253 16677 11287 16711
rect 2789 16609 2823 16643
rect 4353 16609 4387 16643
rect 6561 16609 6595 16643
rect 8677 16609 8711 16643
rect 9137 16609 9171 16643
rect 12081 16609 12115 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 3893 16541 3927 16575
rect 4169 16541 4203 16575
rect 4905 16541 4939 16575
rect 5365 16541 5399 16575
rect 5549 16541 5583 16575
rect 5825 16541 5859 16575
rect 6285 16541 6319 16575
rect 6377 16541 6411 16575
rect 7021 16541 7055 16575
rect 7297 16541 7331 16575
rect 8125 16541 8159 16575
rect 8401 16541 8435 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 9873 16541 9907 16575
rect 12265 16541 12299 16575
rect 12541 16541 12575 16575
rect 12817 16541 12851 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 14105 16541 14139 16575
rect 2522 16473 2556 16507
rect 3525 16473 3559 16507
rect 10140 16473 10174 16507
rect 12909 16473 12943 16507
rect 1409 16405 1443 16439
rect 4077 16405 4111 16439
rect 4813 16405 4847 16439
rect 4997 16405 5031 16439
rect 5181 16405 5215 16439
rect 5917 16405 5951 16439
rect 6101 16405 6135 16439
rect 7389 16405 7423 16439
rect 7941 16405 7975 16439
rect 8217 16405 8251 16439
rect 9597 16405 9631 16439
rect 11529 16405 11563 16439
rect 12357 16405 12391 16439
rect 13829 16405 13863 16439
rect 14289 16405 14323 16439
rect 3249 16201 3283 16235
rect 4537 16201 4571 16235
rect 7205 16201 7239 16235
rect 8769 16201 8803 16235
rect 11253 16201 11287 16235
rect 4813 16133 4847 16167
rect 5549 16133 5583 16167
rect 5641 16133 5675 16167
rect 1777 16065 1811 16099
rect 2781 16065 2815 16099
rect 3065 16065 3099 16099
rect 3341 16065 3375 16099
rect 3617 16065 3651 16099
rect 3893 16065 3927 16099
rect 6469 16065 6503 16099
rect 7665 16065 7699 16099
rect 8125 16065 8159 16099
rect 10342 16065 10376 16099
rect 10609 16065 10643 16099
rect 10885 16065 10919 16099
rect 11161 16065 11195 16099
rect 11529 16065 11563 16099
rect 11796 16065 11830 16099
rect 13921 16065 13955 16099
rect 14197 16065 14231 16099
rect 2421 15997 2455 16031
rect 2605 15997 2639 16031
rect 4077 15997 4111 16031
rect 4721 15997 4755 16031
rect 6653 15997 6687 16031
rect 7849 15997 7883 16031
rect 8309 15997 8343 16031
rect 10793 15997 10827 16031
rect 13093 15997 13127 16031
rect 3433 15929 3467 15963
rect 5273 15929 5307 15963
rect 6101 15929 6135 15963
rect 13737 15929 13771 15963
rect 1501 15861 1535 15895
rect 2237 15861 2271 15895
rect 2881 15861 2915 15895
rect 3709 15861 3743 15895
rect 7021 15861 7055 15895
rect 9229 15861 9263 15895
rect 12909 15861 12943 15895
rect 13645 15861 13679 15895
rect 14381 15861 14415 15895
rect 2605 15657 2639 15691
rect 3525 15657 3559 15691
rect 3801 15657 3835 15691
rect 4077 15657 4111 15691
rect 4813 15657 4847 15691
rect 5733 15657 5767 15691
rect 7021 15657 7055 15691
rect 8033 15657 8067 15691
rect 1869 15589 1903 15623
rect 3341 15589 3375 15623
rect 10793 15589 10827 15623
rect 12817 15589 12851 15623
rect 2881 15521 2915 15555
rect 4537 15521 4571 15555
rect 5917 15521 5951 15555
rect 6561 15521 6595 15555
rect 7573 15521 7607 15555
rect 9965 15521 9999 15555
rect 12265 15521 12299 15555
rect 12633 15521 12667 15555
rect 13277 15521 13311 15555
rect 1409 15453 1443 15487
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 2697 15453 2731 15487
rect 3617 15453 3651 15487
rect 3985 15453 4019 15487
rect 4721 15453 4755 15487
rect 4997 15453 5031 15487
rect 5549 15453 5583 15487
rect 6009 15453 6043 15487
rect 6285 15453 6319 15487
rect 6377 15453 6411 15487
rect 7389 15453 7423 15487
rect 8125 15453 8159 15487
rect 8309 15453 8343 15487
rect 9137 15453 9171 15487
rect 11161 15453 11195 15487
rect 11253 15453 11287 15487
rect 12357 15453 12391 15487
rect 12449 15453 12483 15487
rect 14289 15453 14323 15487
rect 8769 15385 8803 15419
rect 10241 15385 10275 15419
rect 10333 15385 10367 15419
rect 13369 15385 13403 15419
rect 13921 15385 13955 15419
rect 1593 15317 1627 15351
rect 6101 15317 6135 15351
rect 8953 15317 8987 15351
rect 9321 15317 9355 15351
rect 10977 15317 11011 15351
rect 11437 15317 11471 15351
rect 14197 15317 14231 15351
rect 1593 15113 1627 15147
rect 3433 15113 3467 15147
rect 8309 15113 8343 15147
rect 9965 15113 9999 15147
rect 12173 15113 12207 15147
rect 9229 15045 9263 15079
rect 10609 15045 10643 15079
rect 11161 15045 11195 15079
rect 13654 15045 13688 15079
rect 1685 14977 1719 15011
rect 1777 14977 1811 15011
rect 2513 14977 2547 15011
rect 2789 14977 2823 15011
rect 2973 14977 3007 15011
rect 3525 14977 3559 15011
rect 3985 14977 4019 15011
rect 4077 14977 4111 15011
rect 4537 14977 4571 15011
rect 7665 14977 7699 15011
rect 9321 14977 9355 15011
rect 10149 14977 10183 15011
rect 11529 14977 11563 15011
rect 12449 14977 12483 15011
rect 13921 14977 13955 15011
rect 14197 14977 14231 15011
rect 1961 14909 1995 14943
rect 7205 14909 7239 14943
rect 7849 14909 7883 14943
rect 8585 14909 8619 14943
rect 9505 14909 9539 14943
rect 11253 14909 11287 14943
rect 11713 14909 11747 14943
rect 12357 14909 12391 14943
rect 3801 14841 3835 14875
rect 2421 14773 2455 14807
rect 3709 14773 3743 14807
rect 4169 14773 4203 14807
rect 4721 14773 4755 14807
rect 6653 14773 6687 14807
rect 10333 14773 10367 14807
rect 12541 14773 12575 14807
rect 14381 14773 14415 14807
rect 2697 14569 2731 14603
rect 4445 14569 4479 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 9045 14569 9079 14603
rect 10149 14569 10183 14603
rect 12173 14569 12207 14603
rect 12817 14569 12851 14603
rect 13829 14501 13863 14535
rect 4261 14433 4295 14467
rect 7665 14433 7699 14467
rect 10977 14433 11011 14467
rect 11713 14433 11747 14467
rect 12633 14433 12667 14467
rect 13277 14433 13311 14467
rect 1409 14365 1443 14399
rect 2329 14365 2363 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 5457 14365 5491 14399
rect 6929 14365 6963 14399
rect 7481 14365 7515 14399
rect 8125 14365 8159 14399
rect 8585 14365 8619 14399
rect 9229 14365 9263 14399
rect 9965 14365 9999 14399
rect 10241 14365 10275 14399
rect 11069 14365 11103 14399
rect 11529 14365 11563 14399
rect 12449 14365 12483 14399
rect 14289 14365 14323 14399
rect 1777 14297 1811 14331
rect 2237 14297 2271 14331
rect 6684 14297 6718 14331
rect 10333 14297 10367 14331
rect 13369 14297 13403 14331
rect 2421 14229 2455 14263
rect 3341 14229 3375 14263
rect 3525 14229 3559 14263
rect 3985 14229 4019 14263
rect 4813 14229 4847 14263
rect 5549 14229 5583 14263
rect 7021 14229 7055 14263
rect 9321 14229 9355 14263
rect 11253 14229 11287 14263
rect 14105 14229 14139 14263
rect 1593 14025 1627 14059
rect 2513 14025 2547 14059
rect 2881 14025 2915 14059
rect 7297 14025 7331 14059
rect 7573 14025 7607 14059
rect 9137 14025 9171 14059
rect 10609 14025 10643 14059
rect 11345 14025 11379 14059
rect 11529 14025 11563 14059
rect 12633 14025 12667 14059
rect 12725 14025 12759 14059
rect 13737 14025 13771 14059
rect 4005 13957 4039 13991
rect 1777 13889 1811 13923
rect 4261 13889 4295 13923
rect 4537 13889 4571 13923
rect 5273 13889 5307 13923
rect 5457 13889 5491 13923
rect 5733 13889 5767 13923
rect 7113 13889 7147 13923
rect 7665 13889 7699 13923
rect 7757 13889 7791 13923
rect 8024 13889 8058 13923
rect 9229 13889 9263 13923
rect 9485 13889 9519 13923
rect 10885 13889 10919 13923
rect 11713 13889 11747 13923
rect 13921 13889 13955 13923
rect 14105 13889 14139 13923
rect 1869 13821 1903 13855
rect 2053 13821 2087 13855
rect 4629 13821 4663 13855
rect 5549 13821 5583 13855
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 10701 13821 10735 13855
rect 11989 13821 12023 13855
rect 12173 13821 12207 13855
rect 13185 13821 13219 13855
rect 13369 13821 13403 13855
rect 4905 13753 4939 13787
rect 5917 13753 5951 13787
rect 6377 13753 6411 13787
rect 14381 13685 14415 13719
rect 1685 13481 1719 13515
rect 2421 13481 2455 13515
rect 3617 13481 3651 13515
rect 4261 13481 4295 13515
rect 7205 13481 7239 13515
rect 9045 13481 9079 13515
rect 9965 13481 9999 13515
rect 10977 13481 11011 13515
rect 12909 13481 12943 13515
rect 13277 13481 13311 13515
rect 12173 13413 12207 13447
rect 2237 13345 2271 13379
rect 7389 13345 7423 13379
rect 10149 13345 10183 13379
rect 10517 13345 10551 13379
rect 13369 13345 13403 13379
rect 1777 13277 1811 13311
rect 2053 13277 2087 13311
rect 3065 13277 3099 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 4537 13277 4571 13311
rect 4997 13277 5031 13311
rect 7021 13277 7055 13311
rect 7113 13277 7147 13311
rect 8953 13277 8987 13311
rect 9413 13277 9447 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 12541 13277 12575 13311
rect 12817 13277 12851 13311
rect 13093 13277 13127 13311
rect 14289 13277 14323 13311
rect 7656 13209 7690 13243
rect 4721 13141 4755 13175
rect 5089 13141 5123 13175
rect 5549 13141 5583 13175
rect 8769 13141 8803 13175
rect 9229 13141 9263 13175
rect 9689 13141 9723 13175
rect 11713 13141 11747 13175
rect 12725 13141 12759 13175
rect 14105 13141 14139 13175
rect 1961 12937 1995 12971
rect 2237 12937 2271 12971
rect 3433 12937 3467 12971
rect 4169 12937 4203 12971
rect 5641 12937 5675 12971
rect 5917 12937 5951 12971
rect 6193 12937 6227 12971
rect 7573 12937 7607 12971
rect 9321 12937 9355 12971
rect 10793 12937 10827 12971
rect 11529 12937 11563 12971
rect 13829 12937 13863 12971
rect 6929 12869 6963 12903
rect 7021 12869 7055 12903
rect 7849 12869 7883 12903
rect 10977 12869 11011 12903
rect 14105 12869 14139 12903
rect 1593 12801 1627 12835
rect 1869 12801 1903 12835
rect 2145 12801 2179 12835
rect 2697 12801 2731 12835
rect 3157 12801 3191 12835
rect 3249 12801 3283 12835
rect 3525 12801 3559 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 6009 12801 6043 12835
rect 7297 12801 7331 12835
rect 7757 12801 7791 12835
rect 9689 12801 9723 12835
rect 10149 12801 10183 12835
rect 10885 12801 10919 12835
rect 11713 12801 11747 12835
rect 11805 12801 11839 12835
rect 12541 12801 12575 12835
rect 13553 12801 13587 12835
rect 13645 12801 13679 12835
rect 3065 12733 3099 12767
rect 3709 12733 3743 12767
rect 4445 12733 4479 12767
rect 6745 12733 6779 12767
rect 10333 12733 10367 12767
rect 1777 12665 1811 12699
rect 2881 12597 2915 12631
rect 4629 12597 4663 12631
rect 5181 12597 5215 12631
rect 7389 12597 7423 12631
rect 9873 12597 9907 12631
rect 11897 12597 11931 12631
rect 12725 12597 12759 12631
rect 13461 12597 13495 12631
rect 14381 12597 14415 12631
rect 1593 12393 1627 12427
rect 12633 12393 12667 12427
rect 14105 12393 14139 12427
rect 4169 12325 4203 12359
rect 4629 12325 4663 12359
rect 6009 12325 6043 12359
rect 7849 12325 7883 12359
rect 10057 12325 10091 12359
rect 10425 12325 10459 12359
rect 2053 12257 2087 12291
rect 2973 12257 3007 12291
rect 4813 12257 4847 12291
rect 6377 12257 6411 12291
rect 8309 12257 8343 12291
rect 8493 12257 8527 12291
rect 9045 12257 9079 12291
rect 10977 12257 11011 12291
rect 1409 12189 1443 12223
rect 1777 12189 1811 12223
rect 2237 12189 2271 12223
rect 3157 12189 3191 12223
rect 3801 12189 3835 12223
rect 4077 12189 4111 12223
rect 4997 12189 5031 12223
rect 6193 12189 6227 12223
rect 6633 12189 6667 12223
rect 8769 12189 8803 12223
rect 9873 12189 9907 12223
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 11244 12189 11278 12223
rect 12449 12189 12483 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 1869 12121 1903 12155
rect 5181 12121 5215 12155
rect 5273 12121 5307 12155
rect 5825 12121 5859 12155
rect 9137 12121 9171 12155
rect 9689 12121 9723 12155
rect 13461 12121 13495 12155
rect 2697 12053 2731 12087
rect 3617 12053 3651 12087
rect 3985 12053 4019 12087
rect 7757 12053 7791 12087
rect 8677 12053 8711 12087
rect 12357 12053 12391 12087
rect 13645 12053 13679 12087
rect 2973 11849 3007 11883
rect 4169 11849 4203 11883
rect 7665 11849 7699 11883
rect 11253 11849 11287 11883
rect 11897 11849 11931 11883
rect 12633 11849 12667 11883
rect 13553 11849 13587 11883
rect 7757 11781 7791 11815
rect 1501 11713 1535 11747
rect 1777 11713 1811 11747
rect 2053 11713 2087 11747
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 3341 11713 3375 11747
rect 4261 11713 4295 11747
rect 5845 11713 5879 11747
rect 6101 11713 6135 11747
rect 6377 11713 6411 11747
rect 6929 11713 6963 11747
rect 9597 11713 9631 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 12265 11713 12299 11747
rect 12541 11713 12575 11747
rect 13093 11713 13127 11747
rect 13737 11713 13771 11747
rect 13921 11713 13955 11747
rect 2237 11645 2271 11679
rect 3525 11645 3559 11679
rect 7021 11645 7055 11679
rect 10885 11645 10919 11679
rect 12909 11645 12943 11679
rect 3249 11577 3283 11611
rect 6561 11577 6595 11611
rect 9045 11577 9079 11611
rect 12449 11577 12483 11611
rect 1685 11509 1719 11543
rect 1869 11509 1903 11543
rect 2421 11509 2455 11543
rect 3709 11509 3743 11543
rect 4721 11509 4755 11543
rect 6837 11509 6871 11543
rect 10241 11509 10275 11543
rect 10333 11509 10367 11543
rect 11529 11509 11563 11543
rect 14105 11509 14139 11543
rect 1961 11305 1995 11339
rect 8769 11305 8803 11339
rect 10425 11305 10459 11339
rect 11989 11305 12023 11339
rect 14381 11305 14415 11339
rect 4629 11237 4663 11271
rect 6837 11237 6871 11271
rect 11805 11237 11839 11271
rect 2329 11169 2363 11203
rect 2973 11169 3007 11203
rect 4997 11169 5031 11203
rect 7389 11169 7423 11203
rect 10885 11169 10919 11203
rect 11161 11169 11195 11203
rect 11345 11169 11379 11203
rect 12265 11169 12299 11203
rect 13277 11169 13311 11203
rect 1685 11101 1719 11135
rect 1777 11101 1811 11135
rect 2145 11101 2179 11135
rect 3157 11101 3191 11135
rect 4813 11101 4847 11135
rect 5181 11101 5215 11135
rect 5273 11101 5307 11135
rect 5457 11101 5491 11135
rect 7113 11101 7147 11135
rect 7656 11101 7690 11135
rect 10077 11101 10111 11135
rect 10333 11101 10367 11135
rect 11069 11101 11103 11135
rect 11897 11101 11931 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 13461 11101 13495 11135
rect 14197 11101 14231 11135
rect 2789 11033 2823 11067
rect 5724 11033 5758 11067
rect 13921 11033 13955 11067
rect 1593 10965 1627 10999
rect 3617 10965 3651 10999
rect 6929 10965 6963 10999
rect 8953 10965 8987 10999
rect 13185 10965 13219 10999
rect 1777 10761 1811 10795
rect 2697 10761 2731 10795
rect 3525 10761 3559 10795
rect 5365 10761 5399 10795
rect 6653 10761 6687 10795
rect 10425 10761 10459 10795
rect 14105 10761 14139 10795
rect 6929 10693 6963 10727
rect 7757 10693 7791 10727
rect 9137 10693 9171 10727
rect 1593 10625 1627 10659
rect 3249 10625 3283 10659
rect 3617 10625 3651 10659
rect 3893 10625 3927 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 4813 10625 4847 10659
rect 5641 10625 5675 10659
rect 6469 10625 6503 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 9965 10625 9999 10659
rect 10609 10625 10643 10659
rect 11161 10625 11195 10659
rect 11529 10625 11563 10659
rect 12265 10625 12299 10659
rect 13185 10625 13219 10659
rect 13461 10625 13495 10659
rect 13645 10625 13679 10659
rect 14197 10625 14231 10659
rect 2053 10557 2087 10591
rect 2237 10557 2271 10591
rect 2789 10557 2823 10591
rect 6837 10557 6871 10591
rect 7665 10557 7699 10591
rect 9045 10557 9079 10591
rect 9413 10557 9447 10591
rect 11713 10557 11747 10591
rect 12449 10557 12483 10591
rect 7389 10489 7423 10523
rect 8217 10489 8251 10523
rect 8861 10489 8895 10523
rect 11345 10489 11379 10523
rect 13001 10489 13035 10523
rect 3065 10421 3099 10455
rect 3801 10421 3835 10455
rect 4077 10421 4111 10455
rect 4353 10421 4387 10455
rect 5457 10421 5491 10455
rect 8401 10421 8435 10455
rect 9873 10421 9907 10455
rect 12173 10421 12207 10455
rect 12817 10421 12851 10455
rect 14381 10421 14415 10455
rect 1685 10217 1719 10251
rect 3617 10217 3651 10251
rect 4169 10217 4203 10251
rect 5917 10217 5951 10251
rect 6285 10217 6319 10251
rect 8493 10217 8527 10251
rect 11161 10217 11195 10251
rect 11621 10217 11655 10251
rect 12173 10217 12207 10251
rect 14105 10217 14139 10251
rect 4537 10149 4571 10183
rect 5181 10149 5215 10183
rect 5457 10081 5491 10115
rect 7205 10081 7239 10115
rect 7389 10081 7423 10115
rect 9689 10081 9723 10115
rect 1409 10013 1443 10047
rect 1869 10013 1903 10047
rect 1961 10013 1995 10047
rect 2237 10013 2271 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4721 10013 4755 10047
rect 4997 10013 5031 10047
rect 5273 10013 5307 10047
rect 6469 10013 6503 10047
rect 6653 10013 6687 10047
rect 6745 10013 6779 10047
rect 8125 10013 8159 10047
rect 8309 10013 8343 10047
rect 8401 10013 8435 10047
rect 8677 10013 8711 10047
rect 9229 10013 9263 10047
rect 9505 10013 9539 10047
rect 10241 10013 10275 10047
rect 10425 10013 10459 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 12265 10013 12299 10047
rect 13829 10013 13863 10047
rect 14289 10013 14323 10047
rect 2504 9945 2538 9979
rect 7481 9945 7515 9979
rect 13562 9945 13596 9979
rect 1593 9877 1627 9911
rect 2053 9877 2087 9911
rect 9413 9877 9447 9911
rect 10149 9877 10183 9911
rect 10885 9877 10919 9911
rect 12449 9877 12483 9911
rect 2973 9673 3007 9707
rect 3893 9673 3927 9707
rect 6009 9673 6043 9707
rect 6929 9673 6963 9707
rect 7113 9673 7147 9707
rect 8401 9673 8435 9707
rect 9597 9673 9631 9707
rect 10057 9673 10091 9707
rect 12909 9673 12943 9707
rect 1685 9537 1719 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 3709 9537 3743 9571
rect 4077 9537 4111 9571
rect 4169 9537 4203 9571
rect 4353 9537 4387 9571
rect 4629 9537 4663 9571
rect 4905 9537 4939 9571
rect 5917 9537 5951 9571
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 7021 9537 7055 9571
rect 7665 9537 7699 9571
rect 9045 9537 9079 9571
rect 9321 9537 9355 9571
rect 9781 9537 9815 9571
rect 10241 9537 10275 9571
rect 11713 9537 11747 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 12725 9537 12759 9571
rect 14381 9537 14415 9571
rect 1409 9469 1443 9503
rect 2329 9469 2363 9503
rect 2513 9469 2547 9503
rect 3157 9469 3191 9503
rect 5181 9469 5215 9503
rect 5365 9469 5399 9503
rect 5825 9469 5859 9503
rect 7481 9469 7515 9503
rect 8125 9469 8159 9503
rect 8861 9469 8895 9503
rect 10425 9469 10459 9503
rect 13461 9469 13495 9503
rect 13645 9469 13679 9503
rect 14197 9469 14231 9503
rect 3617 9401 3651 9435
rect 4537 9401 4571 9435
rect 4813 9401 4847 9435
rect 9137 9401 9171 9435
rect 12265 9401 12299 9435
rect 4997 9333 5031 9367
rect 6377 9333 6411 9367
rect 10701 9333 10735 9367
rect 11897 9333 11931 9367
rect 12633 9333 12667 9367
rect 13277 9333 13311 9367
rect 13737 9333 13771 9367
rect 2145 9129 2179 9163
rect 3433 9129 3467 9163
rect 5641 9129 5675 9163
rect 8309 9129 8343 9163
rect 10517 9129 10551 9163
rect 14289 9129 14323 9163
rect 3157 9061 3191 9095
rect 3801 9061 3835 9095
rect 6837 9061 6871 9095
rect 7297 9061 7331 9095
rect 11437 9061 11471 9095
rect 11713 9061 11747 9095
rect 2513 8993 2547 9027
rect 5365 8993 5399 9027
rect 6193 8993 6227 9027
rect 6377 8993 6411 9027
rect 7849 8993 7883 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 13185 8993 13219 9027
rect 13369 8993 13403 9027
rect 1777 8925 1811 8959
rect 2329 8925 2363 8959
rect 2789 8925 2823 8959
rect 2881 8925 2915 8959
rect 3341 8925 3375 8959
rect 3617 8925 3651 8959
rect 3985 8925 4019 8959
rect 4629 8925 4663 8959
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 5181 8925 5215 8959
rect 6101 8925 6135 8959
rect 6929 8925 6963 8959
rect 7113 8925 7147 8959
rect 7665 8925 7699 8959
rect 9413 8925 9447 8959
rect 9873 8925 9907 8959
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 13093 8925 13127 8959
rect 14105 8925 14139 8959
rect 4997 8857 5031 8891
rect 6009 8857 6043 8891
rect 10885 8857 10919 8891
rect 10977 8857 11011 8891
rect 12173 8857 12207 8891
rect 12265 8857 12299 8891
rect 13829 8857 13863 8891
rect 1685 8789 1719 8823
rect 2605 8789 2639 8823
rect 2973 8789 3007 8823
rect 4169 8789 4203 8823
rect 8401 8789 8435 8823
rect 8953 8789 8987 8823
rect 10241 8789 10275 8823
rect 12449 8789 12483 8823
rect 2973 8585 3007 8619
rect 4353 8585 4387 8619
rect 4629 8585 4663 8619
rect 5733 8585 5767 8619
rect 6009 8585 6043 8619
rect 6561 8585 6595 8619
rect 8585 8585 8619 8619
rect 10701 8585 10735 8619
rect 11069 8585 11103 8619
rect 11805 8585 11839 8619
rect 14289 8585 14323 8619
rect 7757 8517 7791 8551
rect 1685 8449 1719 8483
rect 2421 8449 2455 8483
rect 2697 8449 2731 8483
rect 4445 8449 4479 8483
rect 4721 8449 4755 8483
rect 4813 8449 4847 8483
rect 5181 8449 5215 8483
rect 5917 8449 5951 8483
rect 6193 8449 6227 8483
rect 6377 8449 6411 8483
rect 6837 8449 6871 8483
rect 7113 8449 7147 8483
rect 7389 8449 7423 8483
rect 7665 8449 7699 8483
rect 7941 8449 7975 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 10977 8449 11011 8483
rect 11253 8449 11287 8483
rect 11713 8449 11747 8483
rect 12265 8449 12299 8483
rect 12633 8449 12667 8483
rect 12725 8449 12759 8483
rect 12817 8449 12851 8483
rect 12909 8449 12943 8483
rect 13369 8449 13403 8483
rect 13921 8449 13955 8483
rect 14197 8449 14231 8483
rect 1409 8381 1443 8415
rect 3525 8381 3559 8415
rect 3709 8381 3743 8415
rect 3893 8381 3927 8415
rect 4997 8381 5031 8415
rect 5641 8381 5675 8415
rect 8125 8381 8159 8415
rect 10057 8381 10091 8415
rect 10241 8381 10275 8415
rect 10885 8381 10919 8415
rect 12449 8381 12483 8415
rect 13185 8381 13219 8415
rect 2881 8313 2915 8347
rect 6653 8313 6687 8347
rect 7297 8313 7331 8347
rect 7573 8313 7607 8347
rect 9689 8313 9723 8347
rect 11529 8313 11563 8347
rect 2605 8245 2639 8279
rect 9321 8245 9355 8279
rect 13553 8245 13587 8279
rect 14105 8245 14139 8279
rect 3525 8041 3559 8075
rect 5089 8041 5123 8075
rect 5549 8041 5583 8075
rect 10057 8041 10091 8075
rect 12357 8041 12391 8075
rect 12541 8041 12575 8075
rect 4629 7973 4663 8007
rect 8125 7973 8159 8007
rect 9137 7973 9171 8007
rect 3065 7905 3099 7939
rect 9413 7905 9447 7939
rect 12081 7905 12115 7939
rect 12817 7905 12851 7939
rect 3157 7837 3191 7871
rect 3433 7837 3467 7871
rect 3801 7837 3835 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 11437 7837 11471 7871
rect 12265 7837 12299 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 13553 7837 13587 7871
rect 14289 7837 14323 7871
rect 2820 7769 2854 7803
rect 3249 7769 3283 7803
rect 4353 7769 4387 7803
rect 4445 7769 4479 7803
rect 7021 7769 7055 7803
rect 11192 7769 11226 7803
rect 1593 7701 1627 7735
rect 1685 7701 1719 7735
rect 7849 7701 7883 7735
rect 8493 7701 8527 7735
rect 9873 7701 9907 7735
rect 11529 7701 11563 7735
rect 13461 7701 13495 7735
rect 13737 7701 13771 7735
rect 14105 7701 14139 7735
rect 1409 7497 1443 7531
rect 6377 7497 6411 7531
rect 6929 7497 6963 7531
rect 11253 7497 11287 7531
rect 12633 7497 12667 7531
rect 13093 7497 13127 7531
rect 13369 7497 13403 7531
rect 3065 7429 3099 7463
rect 7849 7429 7883 7463
rect 9597 7429 9631 7463
rect 2533 7361 2567 7395
rect 2789 7361 2823 7395
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 4629 7361 4663 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 9873 7361 9907 7395
rect 10140 7361 10174 7395
rect 12081 7361 12115 7395
rect 12265 7361 12299 7395
rect 12541 7361 12575 7395
rect 13001 7361 13035 7395
rect 13277 7361 13311 7395
rect 13829 7361 13863 7395
rect 14289 7361 14323 7395
rect 2973 7293 3007 7327
rect 4353 7293 4387 7327
rect 5733 7293 5767 7327
rect 5917 7293 5951 7327
rect 14013 7293 14047 7327
rect 5273 7225 5307 7259
rect 7113 7225 7147 7259
rect 11529 7225 11563 7259
rect 3709 7157 3743 7191
rect 4813 7157 4847 7191
rect 6193 7157 6227 7191
rect 7665 7157 7699 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 14105 7157 14139 7191
rect 3065 6953 3099 6987
rect 4261 6953 4295 6987
rect 7849 6953 7883 6987
rect 9781 6953 9815 6987
rect 11069 6953 11103 6987
rect 13461 6953 13495 6987
rect 10333 6885 10367 6919
rect 11345 6885 11379 6919
rect 1409 6817 1443 6851
rect 1685 6817 1719 6851
rect 2421 6817 2455 6851
rect 3801 6817 3835 6851
rect 5273 6817 5307 6851
rect 6377 6817 6411 6851
rect 6837 6817 6871 6851
rect 7113 6817 7147 6851
rect 8309 6817 8343 6851
rect 9137 6817 9171 6851
rect 9321 6817 9355 6851
rect 11897 6817 11931 6851
rect 13645 6817 13679 6851
rect 13829 6817 13863 6851
rect 3341 6749 3375 6783
rect 3985 6749 4019 6783
rect 5089 6749 5123 6783
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 7297 6749 7331 6783
rect 8493 6749 8527 6783
rect 8609 6749 8643 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 11529 6749 11563 6783
rect 11621 6749 11655 6783
rect 12081 6749 12115 6783
rect 12725 6749 12759 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 14289 6749 14323 6783
rect 4629 6681 4663 6715
rect 5365 6681 5399 6715
rect 3525 6613 3559 6647
rect 7757 6613 7791 6647
rect 8677 6613 8711 6647
rect 9965 6613 9999 6647
rect 10517 6613 10551 6647
rect 10885 6613 10919 6647
rect 11805 6613 11839 6647
rect 12541 6613 12575 6647
rect 13093 6613 13127 6647
rect 14105 6613 14139 6647
rect 1961 6409 1995 6443
rect 2789 6409 2823 6443
rect 4077 6409 4111 6443
rect 6377 6409 6411 6443
rect 9965 6409 9999 6443
rect 2697 6341 2731 6375
rect 4261 6341 4295 6375
rect 13001 6341 13035 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 2053 6273 2087 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 4169 6273 4203 6307
rect 4445 6273 4479 6307
rect 5937 6273 5971 6307
rect 6193 6273 6227 6307
rect 8033 6273 8067 6307
rect 8677 6273 8711 6307
rect 8953 6273 8987 6307
rect 9689 6273 9723 6307
rect 11078 6273 11112 6307
rect 11345 6273 11379 6307
rect 12449 6273 12483 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 14105 6273 14139 6307
rect 2237 6205 2271 6239
rect 6837 6205 6871 6239
rect 7021 6205 7055 6239
rect 7757 6205 7791 6239
rect 7941 6205 7975 6239
rect 9137 6205 9171 6239
rect 11529 6205 11563 6239
rect 11713 6205 11747 6239
rect 13093 6205 13127 6239
rect 3801 6137 3835 6171
rect 4629 6137 4663 6171
rect 9781 6137 9815 6171
rect 11897 6137 11931 6171
rect 13645 6137 13679 6171
rect 1593 6069 1627 6103
rect 4813 6069 4847 6103
rect 7573 6069 7607 6103
rect 9321 6069 9355 6103
rect 14197 6069 14231 6103
rect 2697 5865 2731 5899
rect 3893 5865 3927 5899
rect 6285 5865 6319 5899
rect 6653 5865 6687 5899
rect 7205 5865 7239 5899
rect 7481 5865 7515 5899
rect 8125 5865 8159 5899
rect 11529 5865 11563 5899
rect 12725 5865 12759 5899
rect 13369 5865 13403 5899
rect 7849 5797 7883 5831
rect 8217 5797 8251 5831
rect 9689 5797 9723 5831
rect 10149 5797 10183 5831
rect 10885 5797 10919 5831
rect 12541 5797 12575 5831
rect 1685 5729 1719 5763
rect 3065 5729 3099 5763
rect 3249 5729 3283 5763
rect 5273 5729 5307 5763
rect 8677 5729 8711 5763
rect 9229 5729 9263 5763
rect 11161 5729 11195 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 3617 5661 3651 5695
rect 5365 5661 5399 5695
rect 5641 5661 5675 5695
rect 5825 5661 5859 5695
rect 6837 5661 6871 5695
rect 7021 5661 7055 5695
rect 7113 5661 7147 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 9045 5661 9079 5695
rect 9781 5661 9815 5695
rect 9965 5661 9999 5695
rect 10701 5661 10735 5695
rect 10977 5661 11011 5695
rect 11897 5661 11931 5695
rect 12081 5661 12115 5695
rect 12817 5661 12851 5695
rect 13553 5661 13587 5695
rect 13737 5661 13771 5695
rect 14289 5661 14323 5695
rect 5028 5593 5062 5627
rect 1593 5525 1627 5559
rect 2329 5525 2363 5559
rect 3433 5525 3467 5559
rect 5549 5525 5583 5559
rect 14105 5525 14139 5559
rect 2421 5321 2455 5355
rect 3617 5321 3651 5355
rect 4445 5321 4479 5355
rect 5917 5321 5951 5355
rect 8125 5321 8159 5355
rect 8493 5321 8527 5355
rect 8769 5321 8803 5355
rect 11069 5321 11103 5355
rect 11713 5321 11747 5355
rect 12357 5253 12391 5287
rect 12449 5253 12483 5287
rect 13277 5253 13311 5287
rect 13369 5253 13403 5287
rect 1685 5185 1719 5219
rect 3065 5185 3099 5219
rect 3341 5185 3375 5219
rect 3801 5185 3835 5219
rect 3893 5185 3927 5219
rect 4353 5185 4387 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 6009 5185 6043 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 8309 5185 8343 5219
rect 8585 5185 8619 5219
rect 9597 5185 9631 5219
rect 10333 5185 10367 5219
rect 11253 5185 11287 5219
rect 11529 5185 11563 5219
rect 12633 5185 12667 5219
rect 13829 5185 13863 5219
rect 14013 5185 14047 5219
rect 14381 5185 14415 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 4905 5117 4939 5151
rect 5089 5117 5123 5151
rect 5549 5117 5583 5151
rect 6929 5117 6963 5151
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 8861 5117 8895 5151
rect 9413 5117 9447 5151
rect 9781 5117 9815 5151
rect 10517 5117 10551 5151
rect 11989 5117 12023 5151
rect 12817 5117 12851 5151
rect 4077 5049 4111 5083
rect 5273 5049 5307 5083
rect 14197 5049 14231 5083
rect 3433 4981 3467 5015
rect 4169 4981 4203 5015
rect 6469 4981 6503 5015
rect 7113 4981 7147 5015
rect 10149 4981 10183 5015
rect 10701 4981 10735 5015
rect 1961 4777 1995 4811
rect 5549 4777 5583 4811
rect 6745 4777 6779 4811
rect 6837 4777 6871 4811
rect 7481 4777 7515 4811
rect 8033 4777 8067 4811
rect 8769 4777 8803 4811
rect 9045 4777 9079 4811
rect 9689 4777 9723 4811
rect 10057 4777 10091 4811
rect 11345 4777 11379 4811
rect 14197 4777 14231 4811
rect 2789 4709 2823 4743
rect 3249 4709 3283 4743
rect 4997 4709 5031 4743
rect 5273 4709 5307 4743
rect 5825 4709 5859 4743
rect 7113 4709 7147 4743
rect 10885 4709 10919 4743
rect 13829 4709 13863 4743
rect 2145 4641 2179 4675
rect 2329 4641 2363 4675
rect 3065 4641 3099 4675
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 9505 4641 9539 4675
rect 1777 4573 1811 4607
rect 2881 4573 2915 4607
rect 3893 4573 3927 4607
rect 4721 4573 4755 4607
rect 5181 4573 5215 4607
rect 5457 4573 5491 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 7665 4573 7699 4607
rect 8125 4573 8159 4607
rect 8401 4573 8435 4607
rect 8585 4573 8619 4607
rect 9229 4573 9263 4607
rect 9597 4573 9631 4607
rect 9881 4569 9915 4603
rect 10333 4573 10367 4607
rect 10609 4573 10643 4607
rect 11069 4573 11103 4607
rect 11161 4573 11195 4607
rect 11805 4573 11839 4607
rect 12449 4573 12483 4607
rect 14289 4573 14323 4607
rect 1685 4505 1719 4539
rect 4813 4505 4847 4539
rect 11621 4505 11655 4539
rect 12357 4505 12391 4539
rect 12694 4505 12728 4539
rect 4445 4437 4479 4471
rect 8217 4437 8251 4471
rect 10241 4437 10275 4471
rect 10425 4437 10459 4471
rect 3985 4233 4019 4267
rect 5917 4233 5951 4267
rect 7205 4233 7239 4267
rect 13001 4233 13035 4267
rect 4537 4165 4571 4199
rect 10701 4165 10735 4199
rect 11069 4165 11103 4199
rect 1685 4097 1719 4131
rect 2513 4097 2547 4131
rect 2697 4097 2731 4131
rect 3249 4097 3283 4131
rect 4169 4097 4203 4131
rect 5089 4097 5123 4131
rect 5641 4097 5675 4131
rect 6101 4097 6135 4131
rect 6469 4097 6503 4131
rect 6561 4097 6595 4131
rect 6745 4097 6779 4131
rect 7297 4097 7331 4131
rect 7573 4097 7607 4131
rect 8585 4097 8619 4131
rect 10149 4097 10183 4131
rect 10977 4097 11011 4131
rect 12642 4097 12676 4131
rect 12909 4097 12943 4131
rect 14114 4097 14148 4131
rect 14381 4097 14415 4131
rect 1409 4029 1443 4063
rect 3433 4029 3467 4063
rect 4445 4029 4479 4063
rect 5825 4029 5859 4063
rect 6837 4029 6871 4063
rect 7665 4029 7699 4063
rect 7849 4029 7883 4063
rect 8677 4029 8711 4063
rect 8861 4029 8895 4063
rect 9965 4029 9999 4063
rect 10793 4029 10827 4063
rect 3157 3961 3191 3995
rect 3617 3961 3651 3995
rect 8401 3961 8435 3995
rect 9321 3961 9355 3995
rect 5181 3893 5215 3927
rect 7389 3893 7423 3927
rect 8125 3893 8159 3927
rect 9413 3893 9447 3927
rect 11529 3893 11563 3927
rect 1869 3689 1903 3723
rect 7941 3689 7975 3723
rect 8769 3689 8803 3723
rect 12909 3689 12943 3723
rect 13921 3689 13955 3723
rect 14381 3689 14415 3723
rect 1593 3621 1627 3655
rect 2145 3621 2179 3655
rect 3617 3621 3651 3655
rect 3985 3621 4019 3655
rect 5825 3621 5859 3655
rect 7665 3621 7699 3655
rect 10517 3621 10551 3655
rect 12081 3621 12115 3655
rect 13001 3621 13035 3655
rect 6285 3553 6319 3587
rect 8125 3553 8159 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 4445 3485 4479 3519
rect 6009 3485 6043 3519
rect 8033 3485 8067 3519
rect 8309 3485 8343 3519
rect 9137 3485 9171 3519
rect 10701 3485 10735 3519
rect 12265 3485 12299 3519
rect 13185 3485 13219 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 2504 3417 2538 3451
rect 4712 3417 4746 3451
rect 6530 3417 6564 3451
rect 9404 3417 9438 3451
rect 10968 3417 11002 3451
rect 4261 3349 4295 3383
rect 6101 3349 6135 3383
rect 2789 3145 2823 3179
rect 3249 3145 3283 3179
rect 6377 3145 6411 3179
rect 9873 3145 9907 3179
rect 11529 3145 11563 3179
rect 3065 3077 3099 3111
rect 4362 3077 4396 3111
rect 5273 3077 5307 3111
rect 7573 3077 7607 3111
rect 9413 3077 9447 3111
rect 13185 3077 13219 3111
rect 1685 3009 1719 3043
rect 2421 3009 2455 3043
rect 2881 3009 2915 3043
rect 3157 3009 3191 3043
rect 4629 3009 4663 3043
rect 4813 3009 4847 3043
rect 4997 3009 5031 3043
rect 6009 3009 6043 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 8870 3009 8904 3043
rect 9137 3009 9171 3043
rect 10986 3009 11020 3043
rect 11253 3009 11287 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 14197 3009 14231 3043
rect 14473 3009 14507 3043
rect 1409 2941 1443 2975
rect 5181 2941 5215 2975
rect 5457 2941 5491 2975
rect 6929 2941 6963 2975
rect 12081 2941 12115 2975
rect 12817 2873 12851 2907
rect 2605 2805 2639 2839
rect 6193 2805 6227 2839
rect 7297 2805 7331 2839
rect 7757 2805 7791 2839
rect 9505 2805 9539 2839
rect 12449 2805 12483 2839
rect 13461 2805 13495 2839
rect 4721 2601 4755 2635
rect 7757 2601 7791 2635
rect 8493 2601 8527 2635
rect 8769 2601 8803 2635
rect 10977 2601 11011 2635
rect 13829 2601 13863 2635
rect 2053 2533 2087 2567
rect 2421 2533 2455 2567
rect 4629 2533 4663 2567
rect 5825 2533 5859 2567
rect 6377 2533 6411 2567
rect 9597 2533 9631 2567
rect 3157 2465 3191 2499
rect 3985 2465 4019 2499
rect 6837 2465 6871 2499
rect 7297 2465 7331 2499
rect 7849 2465 7883 2499
rect 10149 2465 10183 2499
rect 10425 2465 10459 2499
rect 3433 2397 3467 2431
rect 4169 2397 4203 2431
rect 5273 2397 5307 2431
rect 6009 2397 6043 2431
rect 6193 2397 6227 2431
rect 7021 2397 7055 2431
rect 7113 2397 7147 2431
rect 8585 2397 8619 2431
rect 9045 2397 9079 2431
rect 11345 2397 11379 2431
rect 12173 2397 12207 2431
rect 13277 2397 13311 2431
rect 13921 2397 13955 2431
rect 14105 2397 14139 2431
rect 1501 2329 1535 2363
rect 1685 2329 1719 2363
rect 1869 2329 1903 2363
rect 2237 2329 2271 2363
rect 10057 2329 10091 2363
rect 11621 2329 11655 2363
rect 12725 2329 12759 2363
rect 9137 2261 9171 2295
rect 11161 2261 11195 2295
rect 11713 2261 11747 2295
rect 12265 2261 12299 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 14197 2261 14231 2295
<< metal1 >>
rect 9858 22108 9864 22160
rect 9916 22148 9922 22160
rect 11422 22148 11428 22160
rect 9916 22120 11428 22148
rect 9916 22108 9922 22120
rect 11422 22108 11428 22120
rect 11480 22108 11486 22160
rect 3786 21972 3792 22024
rect 3844 22012 3850 22024
rect 5258 22012 5264 22024
rect 3844 21984 5264 22012
rect 3844 21972 3850 21984
rect 5258 21972 5264 21984
rect 5316 21972 5322 22024
rect 3970 21904 3976 21956
rect 4028 21944 4034 21956
rect 9214 21944 9220 21956
rect 4028 21916 9220 21944
rect 4028 21904 4034 21916
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 8570 21876 8576 21888
rect 3108 21848 8576 21876
rect 3108 21836 3114 21848
rect 8570 21836 8576 21848
rect 8628 21836 8634 21888
rect 1104 21786 14971 21808
rect 1104 21734 4376 21786
rect 4428 21734 4440 21786
rect 4492 21734 4504 21786
rect 4556 21734 4568 21786
rect 4620 21734 4632 21786
rect 4684 21734 7803 21786
rect 7855 21734 7867 21786
rect 7919 21734 7931 21786
rect 7983 21734 7995 21786
rect 8047 21734 8059 21786
rect 8111 21734 11230 21786
rect 11282 21734 11294 21786
rect 11346 21734 11358 21786
rect 11410 21734 11422 21786
rect 11474 21734 11486 21786
rect 11538 21734 14657 21786
rect 14709 21734 14721 21786
rect 14773 21734 14785 21786
rect 14837 21734 14849 21786
rect 14901 21734 14913 21786
rect 14965 21734 14971 21786
rect 1104 21712 14971 21734
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2774 21672 2780 21684
rect 2455 21644 2780 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 2774 21632 2780 21644
rect 2832 21632 2838 21684
rect 3050 21632 3056 21684
rect 3108 21632 3114 21684
rect 3329 21675 3387 21681
rect 3329 21641 3341 21675
rect 3375 21672 3387 21675
rect 4985 21675 5043 21681
rect 3375 21644 4936 21672
rect 3375 21641 3387 21644
rect 3329 21635 3387 21641
rect 2038 21564 2044 21616
rect 2096 21604 2102 21616
rect 2685 21607 2743 21613
rect 2685 21604 2697 21607
rect 2096 21576 2697 21604
rect 2096 21564 2102 21576
rect 2685 21573 2697 21576
rect 2731 21573 2743 21607
rect 4062 21604 4068 21616
rect 2685 21567 2743 21573
rect 3160 21576 4068 21604
rect 1394 21496 1400 21548
rect 1452 21536 1458 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1452 21508 1685 21536
rect 1452 21496 1458 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1780 21468 1808 21499
rect 2130 21496 2136 21548
rect 2188 21496 2194 21548
rect 3160 21545 3188 21576
rect 4062 21564 4068 21576
rect 4120 21564 4126 21616
rect 4908 21604 4936 21644
rect 4985 21641 4997 21675
rect 5031 21672 5043 21675
rect 5534 21672 5540 21684
rect 5031 21644 5540 21672
rect 5031 21641 5043 21644
rect 4985 21635 5043 21641
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 5810 21672 5816 21684
rect 5644 21644 5816 21672
rect 5258 21604 5264 21616
rect 4908 21576 5264 21604
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21505 2927 21539
rect 2869 21499 2927 21505
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 992 21440 1808 21468
rect 2884 21468 2912 21499
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 3786 21496 3792 21548
rect 3844 21496 3850 21548
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4798 21536 4804 21548
rect 4663 21508 4804 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 2884 21440 3464 21468
rect 992 21428 998 21440
rect 3436 21344 3464 21440
rect 4246 21428 4252 21480
rect 4304 21428 4310 21480
rect 4356 21468 4384 21499
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 4908 21545 4936 21576
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 5166 21496 5172 21548
rect 5224 21496 5230 21548
rect 5644 21545 5672 21644
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 7561 21675 7619 21681
rect 5951 21644 7144 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 6822 21604 6828 21616
rect 5736 21576 6828 21604
rect 5736 21545 5764 21576
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 6914 21564 6920 21616
rect 6972 21564 6978 21616
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21536 6055 21539
rect 6365 21539 6423 21545
rect 6043 21508 6224 21536
rect 6043 21505 6055 21508
rect 5997 21499 6055 21505
rect 6086 21468 6092 21480
rect 4356 21440 6092 21468
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 3513 21403 3571 21409
rect 3513 21369 3525 21403
rect 3559 21400 3571 21403
rect 4525 21403 4583 21409
rect 3559 21372 4476 21400
rect 3559 21369 3571 21372
rect 3513 21363 3571 21369
rect 1578 21292 1584 21344
rect 1636 21292 1642 21344
rect 3418 21292 3424 21344
rect 3476 21292 3482 21344
rect 3970 21292 3976 21344
rect 4028 21292 4034 21344
rect 4448 21332 4476 21372
rect 4525 21369 4537 21403
rect 4571 21400 4583 21403
rect 6196 21400 6224 21508
rect 6365 21505 6377 21539
rect 6411 21536 6423 21539
rect 6932 21536 6960 21564
rect 6411 21508 6960 21536
rect 6411 21505 6423 21508
rect 6365 21499 6423 21505
rect 7006 21496 7012 21548
rect 7064 21496 7070 21548
rect 7116 21545 7144 21644
rect 7561 21641 7573 21675
rect 7607 21641 7619 21675
rect 7561 21635 7619 21641
rect 7576 21604 7604 21635
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 7837 21675 7895 21681
rect 7837 21672 7849 21675
rect 7708 21644 7849 21672
rect 7708 21632 7714 21644
rect 7837 21641 7849 21644
rect 7883 21641 7895 21675
rect 7837 21635 7895 21641
rect 8478 21632 8484 21684
rect 8536 21632 8542 21684
rect 8570 21632 8576 21684
rect 8628 21632 8634 21684
rect 9030 21632 9036 21684
rect 9088 21672 9094 21684
rect 9309 21675 9367 21681
rect 9309 21672 9321 21675
rect 9088 21644 9321 21672
rect 9088 21632 9094 21644
rect 9309 21641 9321 21644
rect 9355 21641 9367 21675
rect 9309 21635 9367 21641
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 9824 21644 10057 21672
rect 9824 21632 9830 21644
rect 10045 21641 10057 21644
rect 10091 21641 10103 21675
rect 10045 21635 10103 21641
rect 10778 21632 10784 21684
rect 10836 21632 10842 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11204 21644 11713 21672
rect 11204 21632 11210 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 14093 21675 14151 21681
rect 14093 21672 14105 21675
rect 13412 21644 14105 21672
rect 13412 21632 13418 21644
rect 14093 21641 14105 21644
rect 14139 21641 14151 21675
rect 14093 21635 14151 21641
rect 8389 21607 8447 21613
rect 8389 21604 8401 21607
rect 7576 21576 8401 21604
rect 8389 21573 8401 21576
rect 8435 21573 8447 21607
rect 8588 21604 8616 21632
rect 11609 21607 11667 21613
rect 11609 21604 11621 21607
rect 8588 21576 11621 21604
rect 8389 21567 8447 21573
rect 11609 21573 11621 21576
rect 11655 21573 11667 21607
rect 11609 21567 11667 21573
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 7340 21508 7389 21536
rect 7340 21496 7346 21508
rect 7377 21505 7389 21508
rect 7423 21505 7435 21539
rect 7377 21499 7435 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 6917 21471 6975 21477
rect 6917 21437 6929 21471
rect 6963 21468 6975 21471
rect 7760 21468 7788 21499
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 8536 21508 9229 21536
rect 8536 21496 8542 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 11333 21539 11391 21545
rect 11333 21505 11345 21539
rect 11379 21536 11391 21539
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 11379 21508 12081 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 14458 21536 14464 21548
rect 14323 21508 14464 21536
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 6963 21440 7788 21468
rect 6963 21437 6975 21440
rect 6917 21431 6975 21437
rect 10134 21428 10140 21480
rect 10192 21468 10198 21480
rect 11348 21468 11376 21499
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 10192 21440 11376 21468
rect 12437 21471 12495 21477
rect 10192 21428 10198 21440
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 4571 21372 6224 21400
rect 6549 21403 6607 21409
rect 4571 21369 4583 21372
rect 4525 21363 4583 21369
rect 6549 21369 6561 21403
rect 6595 21400 6607 21403
rect 7374 21400 7380 21412
rect 6595 21372 7380 21400
rect 6595 21369 6607 21372
rect 6549 21363 6607 21369
rect 7374 21360 7380 21372
rect 7432 21360 7438 21412
rect 7926 21360 7932 21412
rect 7984 21400 7990 21412
rect 12452 21400 12480 21431
rect 12618 21428 12624 21480
rect 12676 21428 12682 21480
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 13173 21471 13231 21477
rect 13173 21468 13185 21471
rect 12860 21440 13185 21468
rect 12860 21428 12866 21440
rect 13173 21437 13185 21440
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 7984 21372 12480 21400
rect 13081 21403 13139 21409
rect 7984 21360 7990 21372
rect 13081 21369 13093 21403
rect 13127 21400 13139 21403
rect 13127 21372 14044 21400
rect 13127 21369 13139 21372
rect 13081 21363 13139 21369
rect 14016 21344 14044 21372
rect 4706 21332 4712 21344
rect 4448 21304 4712 21332
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 4982 21332 4988 21344
rect 4847 21304 4988 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 4982 21292 4988 21304
rect 5040 21292 5046 21344
rect 5350 21292 5356 21344
rect 5408 21292 5414 21344
rect 5442 21292 5448 21344
rect 5500 21292 5506 21344
rect 6089 21335 6147 21341
rect 6089 21301 6101 21335
rect 6135 21332 6147 21335
rect 7098 21332 7104 21344
rect 6135 21304 7104 21332
rect 6135 21301 6147 21304
rect 6089 21295 6147 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 7190 21292 7196 21344
rect 7248 21292 7254 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11241 21335 11299 21341
rect 11241 21332 11253 21335
rect 11112 21304 11253 21332
rect 11112 21292 11118 21304
rect 11241 21301 11253 21304
rect 11287 21301 11299 21335
rect 11241 21295 11299 21301
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 13817 21335 13875 21341
rect 13817 21332 13829 21335
rect 13596 21304 13829 21332
rect 13596 21292 13602 21304
rect 13817 21301 13829 21304
rect 13863 21301 13875 21335
rect 13817 21295 13875 21301
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 1104 21242 14812 21264
rect 1104 21190 2663 21242
rect 2715 21190 2727 21242
rect 2779 21190 2791 21242
rect 2843 21190 2855 21242
rect 2907 21190 2919 21242
rect 2971 21190 6090 21242
rect 6142 21190 6154 21242
rect 6206 21190 6218 21242
rect 6270 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 9517 21242
rect 9569 21190 9581 21242
rect 9633 21190 9645 21242
rect 9697 21190 9709 21242
rect 9761 21190 9773 21242
rect 9825 21190 12944 21242
rect 12996 21190 13008 21242
rect 13060 21190 13072 21242
rect 13124 21190 13136 21242
rect 13188 21190 13200 21242
rect 13252 21190 14812 21242
rect 1104 21168 14812 21190
rect 1486 21088 1492 21140
rect 1544 21088 1550 21140
rect 4246 21088 4252 21140
rect 4304 21088 4310 21140
rect 4985 21131 5043 21137
rect 4985 21097 4997 21131
rect 5031 21128 5043 21131
rect 5902 21128 5908 21140
rect 5031 21100 5908 21128
rect 5031 21097 5043 21100
rect 4985 21091 5043 21097
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 7193 21131 7251 21137
rect 7193 21097 7205 21131
rect 7239 21128 7251 21131
rect 7926 21128 7932 21140
rect 7239 21100 7932 21128
rect 7239 21097 7251 21100
rect 7193 21091 7251 21097
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8478 21088 8484 21140
rect 8536 21088 8542 21140
rect 8757 21131 8815 21137
rect 8757 21097 8769 21131
rect 8803 21128 8815 21131
rect 9950 21128 9956 21140
rect 8803 21100 9956 21128
rect 8803 21097 8815 21100
rect 8757 21091 8815 21097
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 10870 21088 10876 21140
rect 10928 21128 10934 21140
rect 12158 21128 12164 21140
rect 10928 21100 12164 21128
rect 10928 21088 10934 21100
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 15010 21128 15016 21140
rect 12406 21100 15016 21128
rect 3881 21063 3939 21069
rect 3881 21060 3893 21063
rect 2746 21032 3893 21060
rect 2746 20992 2774 21032
rect 3881 21029 3893 21032
rect 3927 21029 3939 21063
rect 4264 21060 4292 21088
rect 11606 21060 11612 21072
rect 4264 21032 6684 21060
rect 3881 21023 3939 21029
rect 2700 20964 2774 20992
rect 2222 20884 2228 20936
rect 2280 20924 2286 20936
rect 2700 20933 2728 20964
rect 3510 20952 3516 21004
rect 3568 20952 3574 21004
rect 3602 20952 3608 21004
rect 3660 20952 3666 21004
rect 5258 20992 5264 21004
rect 5092 20964 5264 20992
rect 2501 20927 2559 20933
rect 2501 20924 2513 20927
rect 2280 20896 2513 20924
rect 2280 20884 2286 20896
rect 2501 20893 2513 20896
rect 2547 20893 2559 20927
rect 2501 20887 2559 20893
rect 2685 20927 2743 20933
rect 2685 20893 2697 20927
rect 2731 20893 2743 20927
rect 2685 20887 2743 20893
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2924 20896 2973 20924
rect 2924 20884 2930 20896
rect 2961 20893 2973 20896
rect 3007 20893 3019 20927
rect 3620 20924 3648 20952
rect 3970 20924 3976 20936
rect 3620 20896 3976 20924
rect 2961 20887 3019 20893
rect 3970 20884 3976 20896
rect 4028 20924 4034 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 4028 20896 4077 20924
rect 4028 20884 4034 20896
rect 4065 20893 4077 20896
rect 4111 20924 4123 20927
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 4111 20896 4169 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 4893 20927 4951 20933
rect 4893 20893 4905 20927
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 1762 20816 1768 20868
rect 1820 20816 1826 20868
rect 1854 20748 1860 20800
rect 1912 20788 1918 20800
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 1912 20760 2053 20788
rect 1912 20748 1918 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 2041 20751 2099 20757
rect 2314 20748 2320 20800
rect 2372 20748 2378 20800
rect 2869 20791 2927 20797
rect 2869 20757 2881 20791
rect 2915 20788 2927 20791
rect 3326 20788 3332 20800
rect 2915 20760 3332 20788
rect 2915 20757 2927 20760
rect 2869 20751 2927 20757
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 4798 20748 4804 20800
rect 4856 20748 4862 20800
rect 4908 20788 4936 20887
rect 5092 20856 5120 20964
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5442 20952 5448 21004
rect 5500 20952 5506 21004
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 5460 20924 5488 20952
rect 5215 20896 5488 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6178 20884 6184 20936
rect 6236 20924 6242 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 6236 20896 6561 20924
rect 6236 20884 6242 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 5537 20859 5595 20865
rect 5537 20856 5549 20859
rect 5092 20828 5549 20856
rect 5537 20825 5549 20828
rect 5583 20825 5595 20859
rect 5537 20819 5595 20825
rect 5718 20816 5724 20868
rect 5776 20816 5782 20868
rect 6656 20856 6684 21032
rect 9968 21032 11612 21060
rect 6733 20995 6791 21001
rect 6733 20961 6745 20995
rect 6779 20992 6791 20995
rect 8113 20995 8171 21001
rect 8113 20992 8125 20995
rect 6779 20964 8125 20992
rect 6779 20961 6791 20964
rect 6733 20955 6791 20961
rect 8113 20961 8125 20964
rect 8159 20961 8171 20995
rect 8113 20955 8171 20961
rect 9968 20936 9996 21032
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 11885 20995 11943 21001
rect 10060 20964 11836 20992
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 7156 20896 7297 20924
rect 7156 20884 7162 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7374 20884 7380 20936
rect 7432 20924 7438 20936
rect 7469 20927 7527 20933
rect 7469 20924 7481 20927
rect 7432 20896 7481 20924
rect 7432 20884 7438 20896
rect 7469 20893 7481 20896
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 8202 20884 8208 20936
rect 8260 20884 8266 20936
rect 8294 20884 8300 20936
rect 8352 20884 8358 20936
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 8846 20924 8852 20936
rect 8619 20896 8852 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 8846 20884 8852 20896
rect 8904 20884 8910 20936
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9950 20924 9956 20936
rect 8987 20896 9956 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 6656 20828 8616 20856
rect 5258 20788 5264 20800
rect 4908 20760 5264 20788
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 5353 20791 5411 20797
rect 5353 20757 5365 20791
rect 5399 20788 5411 20791
rect 5442 20788 5448 20800
rect 5399 20760 5448 20788
rect 5399 20757 5411 20760
rect 5353 20751 5411 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 6454 20748 6460 20800
rect 6512 20748 6518 20800
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 7650 20788 7656 20800
rect 7064 20760 7656 20788
rect 7064 20748 7070 20760
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 8588 20788 8616 20828
rect 8662 20816 8668 20868
rect 8720 20856 8726 20868
rect 9186 20859 9244 20865
rect 9186 20856 9198 20859
rect 8720 20828 9198 20856
rect 8720 20816 8726 20828
rect 9186 20825 9198 20828
rect 9232 20825 9244 20859
rect 9186 20819 9244 20825
rect 10060 20788 10088 20964
rect 10594 20884 10600 20936
rect 10652 20884 10658 20936
rect 10962 20884 10968 20936
rect 11020 20924 11026 20936
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 11020 20896 11253 20924
rect 11020 20884 11026 20896
rect 11241 20893 11253 20896
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 11701 20927 11759 20933
rect 11701 20893 11713 20927
rect 11747 20893 11759 20927
rect 11808 20924 11836 20964
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 12406 20992 12434 21100
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 13817 21063 13875 21069
rect 13817 21029 13829 21063
rect 13863 21060 13875 21063
rect 13863 21032 14136 21060
rect 13863 21029 13875 21032
rect 13817 21023 13875 21029
rect 11931 20964 12434 20992
rect 13265 20995 13323 21001
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 13311 20964 14044 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11808 20896 11989 20924
rect 11701 20887 11759 20893
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 11716 20856 11744 20887
rect 12158 20884 12164 20936
rect 12216 20884 12222 20936
rect 12250 20884 12256 20936
rect 12308 20924 12314 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 12308 20896 12909 20924
rect 12308 20884 12314 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 14016 20868 14044 20964
rect 14108 20936 14136 21032
rect 14090 20884 14096 20936
rect 14148 20884 14154 20936
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 11716 20828 12020 20856
rect 8588 20760 10088 20788
rect 10318 20748 10324 20800
rect 10376 20748 10382 20800
rect 11146 20748 11152 20800
rect 11204 20748 11210 20800
rect 11992 20788 12020 20828
rect 12176 20828 12756 20856
rect 12176 20788 12204 20828
rect 11992 20760 12204 20788
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 12728 20797 12756 20828
rect 12802 20816 12808 20868
rect 12860 20856 12866 20868
rect 13357 20859 13415 20865
rect 13357 20856 13369 20859
rect 12860 20828 13369 20856
rect 12860 20816 12866 20828
rect 13357 20825 13369 20828
rect 13403 20825 13415 20859
rect 13357 20819 13415 20825
rect 13998 20816 14004 20868
rect 14056 20816 14062 20868
rect 12621 20791 12679 20797
rect 12621 20788 12633 20791
rect 12584 20760 12633 20788
rect 12584 20748 12590 20760
rect 12621 20757 12633 20760
rect 12667 20757 12679 20791
rect 12621 20751 12679 20757
rect 12713 20791 12771 20797
rect 12713 20757 12725 20791
rect 12759 20757 12771 20791
rect 12713 20751 12771 20757
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14093 20791 14151 20797
rect 14093 20788 14105 20791
rect 13872 20760 14105 20788
rect 13872 20748 13878 20760
rect 14093 20757 14105 20760
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 1104 20698 14971 20720
rect 1104 20646 4376 20698
rect 4428 20646 4440 20698
rect 4492 20646 4504 20698
rect 4556 20646 4568 20698
rect 4620 20646 4632 20698
rect 4684 20646 7803 20698
rect 7855 20646 7867 20698
rect 7919 20646 7931 20698
rect 7983 20646 7995 20698
rect 8047 20646 8059 20698
rect 8111 20646 11230 20698
rect 11282 20646 11294 20698
rect 11346 20646 11358 20698
rect 11410 20646 11422 20698
rect 11474 20646 11486 20698
rect 11538 20646 14657 20698
rect 14709 20646 14721 20698
rect 14773 20646 14785 20698
rect 14837 20646 14849 20698
rect 14901 20646 14913 20698
rect 14965 20646 14971 20698
rect 1104 20624 14971 20646
rect 2222 20544 2228 20596
rect 2280 20544 2286 20596
rect 2317 20587 2375 20593
rect 2317 20553 2329 20587
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 1765 20519 1823 20525
rect 1765 20485 1777 20519
rect 1811 20516 1823 20519
rect 2332 20516 2360 20547
rect 2406 20544 2412 20596
rect 2464 20584 2470 20596
rect 3418 20584 3424 20596
rect 2464 20556 3424 20584
rect 2464 20544 2470 20556
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 3970 20544 3976 20596
rect 4028 20544 4034 20596
rect 5534 20544 5540 20596
rect 5592 20544 5598 20596
rect 6178 20544 6184 20596
rect 6236 20544 6242 20596
rect 9030 20544 9036 20596
rect 9088 20584 9094 20596
rect 10318 20584 10324 20596
rect 9088 20556 10324 20584
rect 9088 20544 9094 20556
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 10505 20587 10563 20593
rect 10505 20553 10517 20587
rect 10551 20584 10563 20587
rect 10962 20584 10968 20596
rect 10551 20556 10968 20584
rect 10551 20553 10563 20556
rect 10505 20547 10563 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 14182 20584 14188 20596
rect 11256 20556 14188 20584
rect 4332 20519 4390 20525
rect 1811 20488 2360 20516
rect 2608 20488 4108 20516
rect 1811 20485 1823 20488
rect 1765 20479 1823 20485
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20448 2099 20451
rect 2222 20448 2228 20460
rect 2087 20420 2228 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2498 20408 2504 20460
rect 2556 20408 2562 20460
rect 2608 20457 2636 20488
rect 2866 20457 2872 20460
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20417 2651 20451
rect 2860 20448 2872 20457
rect 2827 20420 2872 20448
rect 2593 20411 2651 20417
rect 2860 20411 2872 20420
rect 2866 20408 2872 20411
rect 2924 20408 2930 20460
rect 4080 20392 4108 20488
rect 4332 20485 4344 20519
rect 4378 20516 4390 20519
rect 4798 20516 4804 20528
rect 4378 20488 4804 20516
rect 4378 20485 4390 20488
rect 4332 20479 4390 20485
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 5552 20448 5580 20544
rect 6454 20476 6460 20528
rect 6512 20516 6518 20528
rect 6610 20519 6668 20525
rect 6610 20516 6622 20519
rect 6512 20488 6622 20516
rect 6512 20476 6518 20488
rect 6610 20485 6622 20488
rect 6656 20485 6668 20519
rect 6610 20479 6668 20485
rect 7944 20488 9904 20516
rect 5721 20451 5779 20457
rect 5721 20448 5733 20451
rect 5552 20420 5733 20448
rect 5721 20417 5733 20420
rect 5767 20417 5779 20451
rect 5721 20411 5779 20417
rect 7190 20408 7196 20460
rect 7248 20448 7254 20460
rect 7944 20457 7972 20488
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7248 20420 7941 20448
rect 7248 20408 7254 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8849 20451 8907 20457
rect 8849 20417 8861 20451
rect 8895 20448 8907 20451
rect 9030 20448 9036 20460
rect 8895 20420 9036 20448
rect 8895 20417 8907 20420
rect 8849 20411 8907 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9876 20457 9904 20488
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10594 20408 10600 20460
rect 10652 20408 10658 20460
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 11146 20408 11152 20460
rect 11204 20408 11210 20460
rect 11256 20457 11284 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 11606 20516 11612 20528
rect 11532 20488 11612 20516
rect 11532 20457 11560 20488
rect 11606 20476 11612 20488
rect 11664 20516 11670 20528
rect 13348 20519 13406 20525
rect 11664 20488 13124 20516
rect 11664 20476 11670 20488
rect 13096 20457 13124 20488
rect 13348 20485 13360 20519
rect 13394 20516 13406 20519
rect 13538 20516 13544 20528
rect 13394 20488 13544 20516
rect 13394 20485 13406 20488
rect 13348 20479 13406 20485
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 11241 20451 11299 20457
rect 11241 20417 11253 20451
rect 11287 20417 11299 20451
rect 11241 20411 11299 20417
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11773 20451 11831 20457
rect 11773 20448 11785 20451
rect 11517 20411 11575 20417
rect 11624 20420 11785 20448
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20380 5595 20383
rect 5626 20380 5632 20392
rect 5583 20352 5632 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 6365 20383 6423 20389
rect 6365 20349 6377 20383
rect 6411 20349 6423 20383
rect 6365 20343 6423 20349
rect 934 20204 940 20256
rect 992 20244 998 20256
rect 1489 20247 1547 20253
rect 1489 20244 1501 20247
rect 992 20216 1501 20244
rect 992 20204 998 20216
rect 1489 20213 1501 20216
rect 1535 20213 1547 20247
rect 1489 20207 1547 20213
rect 5445 20247 5503 20253
rect 5445 20213 5457 20247
rect 5491 20244 5503 20247
rect 5718 20244 5724 20256
rect 5491 20216 5724 20244
rect 5491 20213 5503 20216
rect 5445 20207 5503 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 6380 20244 6408 20343
rect 8110 20340 8116 20392
rect 8168 20340 8174 20392
rect 8941 20383 8999 20389
rect 8941 20349 8953 20383
rect 8987 20380 8999 20383
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 8987 20352 9597 20380
rect 8987 20349 8999 20352
rect 8941 20343 8999 20349
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20349 9827 20383
rect 9769 20343 9827 20349
rect 10045 20383 10103 20389
rect 10045 20349 10057 20383
rect 10091 20380 10103 20383
rect 11072 20380 11100 20408
rect 10091 20352 11100 20380
rect 11164 20380 11192 20408
rect 11624 20380 11652 20420
rect 11773 20417 11785 20420
rect 11819 20417 11831 20451
rect 11773 20411 11831 20417
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20417 13139 20451
rect 13081 20411 13139 20417
rect 11164 20352 11652 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 7466 20272 7472 20324
rect 7524 20312 7530 20324
rect 9674 20312 9680 20324
rect 7524 20284 9680 20312
rect 7524 20272 7530 20284
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 6546 20244 6552 20256
rect 6380 20216 6552 20244
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7745 20247 7803 20253
rect 7745 20244 7757 20247
rect 7432 20216 7757 20244
rect 7432 20204 7438 20216
rect 7745 20213 7757 20216
rect 7791 20244 7803 20247
rect 8202 20244 8208 20256
rect 7791 20216 8208 20244
rect 7791 20213 7803 20216
rect 7745 20207 7803 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8573 20247 8631 20253
rect 8573 20213 8585 20247
rect 8619 20244 8631 20247
rect 8754 20244 8760 20256
rect 8619 20216 8760 20244
rect 8619 20213 8631 20216
rect 8573 20207 8631 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 9122 20204 9128 20256
rect 9180 20204 9186 20256
rect 9784 20244 9812 20343
rect 12820 20284 13032 20312
rect 9858 20244 9864 20256
rect 9784 20216 9864 20244
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11149 20247 11207 20253
rect 11149 20213 11161 20247
rect 11195 20244 11207 20247
rect 12820 20244 12848 20284
rect 11195 20216 12848 20244
rect 11195 20213 11207 20216
rect 11149 20207 11207 20213
rect 12894 20204 12900 20256
rect 12952 20204 12958 20256
rect 13004 20244 13032 20284
rect 13446 20244 13452 20256
rect 13004 20216 13452 20244
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 14461 20247 14519 20253
rect 14461 20244 14473 20247
rect 13780 20216 14473 20244
rect 13780 20204 13786 20216
rect 14461 20213 14473 20216
rect 14507 20213 14519 20247
rect 14461 20207 14519 20213
rect 1104 20154 14812 20176
rect 1104 20102 2663 20154
rect 2715 20102 2727 20154
rect 2779 20102 2791 20154
rect 2843 20102 2855 20154
rect 2907 20102 2919 20154
rect 2971 20102 6090 20154
rect 6142 20102 6154 20154
rect 6206 20102 6218 20154
rect 6270 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 9517 20154
rect 9569 20102 9581 20154
rect 9633 20102 9645 20154
rect 9697 20102 9709 20154
rect 9761 20102 9773 20154
rect 9825 20102 12944 20154
rect 12996 20102 13008 20154
rect 13060 20102 13072 20154
rect 13124 20102 13136 20154
rect 13188 20102 13200 20154
rect 13252 20102 14812 20154
rect 1104 20080 14812 20102
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 3936 20012 4844 20040
rect 3936 20000 3942 20012
rect 1765 19975 1823 19981
rect 1765 19941 1777 19975
rect 1811 19941 1823 19975
rect 1765 19935 1823 19941
rect 3513 19975 3571 19981
rect 3513 19941 3525 19975
rect 3559 19972 3571 19975
rect 4706 19972 4712 19984
rect 3559 19944 4712 19972
rect 3559 19941 3571 19944
rect 3513 19935 3571 19941
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1780 19836 1808 19935
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 4816 19972 4844 20012
rect 5994 20000 6000 20052
rect 6052 20040 6058 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 6052 20012 6285 20040
rect 6052 20000 6058 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 6638 20000 6644 20052
rect 6696 20000 6702 20052
rect 8110 20000 8116 20052
rect 8168 20040 8174 20052
rect 8297 20043 8355 20049
rect 8297 20040 8309 20043
rect 8168 20012 8309 20040
rect 8168 20000 8174 20012
rect 8297 20009 8309 20012
rect 8343 20009 8355 20043
rect 9766 20040 9772 20052
rect 8297 20003 8355 20009
rect 8404 20012 9772 20040
rect 6656 19972 6684 20000
rect 4816 19944 6684 19972
rect 8202 19932 8208 19984
rect 8260 19972 8266 19984
rect 8404 19972 8432 20012
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 9858 20000 9864 20052
rect 9916 20040 9922 20052
rect 9953 20043 10011 20049
rect 9953 20040 9965 20043
rect 9916 20012 9965 20040
rect 9916 20000 9922 20012
rect 9953 20009 9965 20012
rect 9999 20009 10011 20043
rect 9953 20003 10011 20009
rect 10505 20043 10563 20049
rect 10505 20009 10517 20043
rect 10551 20040 10563 20043
rect 10686 20040 10692 20052
rect 10551 20012 10692 20040
rect 10551 20009 10563 20012
rect 10505 20003 10563 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 10870 20000 10876 20052
rect 10928 20000 10934 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 11974 20040 11980 20052
rect 11379 20012 11980 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 8260 19944 8432 19972
rect 8665 19975 8723 19981
rect 8260 19932 8266 19944
rect 8665 19941 8677 19975
rect 8711 19972 8723 19975
rect 8711 19944 9168 19972
rect 8711 19941 8723 19944
rect 8665 19935 8723 19941
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 3234 19904 3240 19916
rect 3191 19876 3240 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 3234 19864 3240 19876
rect 3292 19904 3298 19916
rect 4062 19904 4068 19916
rect 3292 19876 4068 19904
rect 3292 19864 3298 19876
rect 4062 19864 4068 19876
rect 4120 19904 4126 19916
rect 6546 19904 6552 19916
rect 4120 19876 6552 19904
rect 4120 19864 4126 19876
rect 6546 19864 6552 19876
rect 6604 19904 6610 19916
rect 9140 19913 9168 19944
rect 9306 19932 9312 19984
rect 9364 19972 9370 19984
rect 10410 19972 10416 19984
rect 9364 19944 10416 19972
rect 9364 19932 9370 19944
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 13722 19972 13728 19984
rect 10520 19944 13728 19972
rect 6641 19907 6699 19913
rect 6641 19904 6653 19907
rect 6604 19876 6653 19904
rect 6604 19864 6610 19876
rect 6641 19873 6653 19876
rect 6687 19873 6699 19907
rect 6641 19867 6699 19873
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 10520 19848 10548 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 10778 19904 10784 19916
rect 10704 19876 10784 19904
rect 3421 19839 3479 19845
rect 3421 19836 3433 19839
rect 1780 19808 3433 19836
rect 1673 19799 1731 19805
rect 1688 19768 1716 19799
rect 2792 19780 2820 19808
rect 3421 19805 3433 19808
rect 3467 19836 3479 19839
rect 3510 19836 3516 19848
rect 3467 19808 3516 19836
rect 3467 19805 3479 19808
rect 3421 19799 3479 19805
rect 3510 19796 3516 19808
rect 3568 19836 3574 19848
rect 3878 19836 3884 19848
rect 3568 19808 3884 19836
rect 3568 19796 3574 19808
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19836 4031 19839
rect 4154 19836 4160 19848
rect 4019 19808 4160 19836
rect 4019 19805 4031 19808
rect 3973 19799 4031 19805
rect 4154 19796 4160 19808
rect 4212 19796 4218 19848
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19805 5779 19839
rect 5721 19799 5779 19805
rect 2222 19768 2228 19780
rect 1688 19740 2228 19768
rect 2222 19728 2228 19740
rect 2280 19728 2286 19780
rect 2774 19728 2780 19780
rect 2832 19728 2838 19780
rect 2900 19771 2958 19777
rect 2900 19737 2912 19771
rect 2946 19768 2958 19771
rect 4062 19768 4068 19780
rect 2946 19740 4068 19768
rect 2946 19737 2958 19740
rect 2900 19731 2958 19737
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 4246 19728 4252 19780
rect 4304 19728 4310 19780
rect 4798 19728 4804 19780
rect 4856 19728 4862 19780
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 5077 19771 5135 19777
rect 5077 19768 5089 19771
rect 4948 19740 5089 19768
rect 4948 19728 4954 19740
rect 5077 19737 5089 19740
rect 5123 19737 5135 19771
rect 5077 19731 5135 19737
rect 1578 19660 1584 19712
rect 1636 19660 1642 19712
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 3050 19700 3056 19712
rect 2004 19672 3056 19700
rect 2004 19660 2010 19672
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 4157 19703 4215 19709
rect 4157 19669 4169 19703
rect 4203 19700 4215 19703
rect 5552 19700 5580 19799
rect 4203 19672 5580 19700
rect 5736 19700 5764 19799
rect 5902 19796 5908 19848
rect 5960 19796 5966 19848
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8754 19796 8760 19848
rect 8812 19836 8818 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8812 19808 8953 19836
rect 8812 19796 8818 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 10045 19839 10103 19845
rect 10045 19805 10057 19839
rect 10091 19805 10103 19839
rect 10045 19799 10103 19805
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 10502 19836 10508 19848
rect 10367 19808 10508 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 5920 19768 5948 19796
rect 6454 19768 6460 19780
rect 5920 19740 6460 19768
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 6908 19771 6966 19777
rect 6908 19737 6920 19771
rect 6954 19768 6966 19771
rect 7006 19768 7012 19780
rect 6954 19740 7012 19768
rect 6954 19737 6966 19740
rect 6908 19731 6966 19737
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 7650 19728 7656 19780
rect 7708 19768 7714 19780
rect 8662 19768 8668 19780
rect 7708 19740 8668 19768
rect 7708 19728 7714 19740
rect 8662 19728 8668 19740
rect 8720 19728 8726 19780
rect 10060 19768 10088 19799
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 10594 19796 10600 19848
rect 10652 19796 10658 19848
rect 10704 19845 10732 19876
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 11517 19907 11575 19913
rect 11517 19873 11529 19907
rect 11563 19904 11575 19907
rect 11790 19904 11796 19916
rect 11563 19876 11796 19904
rect 11563 19873 11575 19876
rect 11517 19867 11575 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 12621 19907 12679 19913
rect 12621 19873 12633 19907
rect 12667 19904 12679 19907
rect 13354 19904 13360 19916
rect 12667 19876 13360 19904
rect 12667 19873 12679 19876
rect 12621 19867 12679 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 11698 19796 11704 19848
rect 11756 19796 11762 19848
rect 12161 19839 12219 19845
rect 12161 19805 12173 19839
rect 12207 19836 12219 19839
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 12207 19808 12449 19836
rect 12207 19805 12219 19808
rect 12161 19799 12219 19805
rect 12437 19805 12449 19808
rect 12483 19836 12495 19839
rect 12526 19836 12532 19848
rect 12483 19808 12532 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 15286 19836 15292 19848
rect 14139 19808 15292 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 10778 19768 10784 19780
rect 10060 19740 10784 19768
rect 10778 19728 10784 19740
rect 10836 19728 10842 19780
rect 11057 19771 11115 19777
rect 11057 19737 11069 19771
rect 11103 19768 11115 19771
rect 11146 19768 11152 19780
rect 11103 19740 11152 19768
rect 11103 19737 11115 19740
rect 11057 19731 11115 19737
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 13081 19771 13139 19777
rect 13081 19737 13093 19771
rect 13127 19768 13139 19771
rect 13262 19768 13268 19780
rect 13127 19740 13268 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 13262 19728 13268 19740
rect 13320 19728 13326 19780
rect 13357 19771 13415 19777
rect 13357 19737 13369 19771
rect 13403 19737 13415 19771
rect 13357 19731 13415 19737
rect 13909 19771 13967 19777
rect 13909 19737 13921 19771
rect 13955 19768 13967 19771
rect 13955 19740 14136 19768
rect 13955 19737 13967 19740
rect 13909 19731 13967 19737
rect 6730 19700 6736 19712
rect 5736 19672 6736 19700
rect 4203 19669 4215 19672
rect 4157 19663 4215 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 8021 19703 8079 19709
rect 8021 19700 8033 19703
rect 7616 19672 8033 19700
rect 7616 19660 7622 19672
rect 8021 19669 8033 19672
rect 8067 19669 8079 19703
rect 8021 19663 8079 19669
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 9585 19703 9643 19709
rect 9585 19700 9597 19703
rect 8352 19672 9597 19700
rect 8352 19660 8358 19672
rect 9585 19669 9597 19672
rect 9631 19669 9643 19703
rect 9585 19663 9643 19669
rect 10137 19703 10195 19709
rect 10137 19669 10149 19703
rect 10183 19700 10195 19703
rect 10226 19700 10232 19712
rect 10183 19672 10232 19700
rect 10183 19669 10195 19672
rect 10137 19663 10195 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 13372 19700 13400 19731
rect 14108 19712 14136 19740
rect 10468 19672 13400 19700
rect 10468 19660 10474 19672
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 14277 19703 14335 19709
rect 14277 19669 14289 19703
rect 14323 19700 14335 19703
rect 14366 19700 14372 19712
rect 14323 19672 14372 19700
rect 14323 19669 14335 19672
rect 14277 19663 14335 19669
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 1104 19610 14971 19632
rect 1104 19558 4376 19610
rect 4428 19558 4440 19610
rect 4492 19558 4504 19610
rect 4556 19558 4568 19610
rect 4620 19558 4632 19610
rect 4684 19558 7803 19610
rect 7855 19558 7867 19610
rect 7919 19558 7931 19610
rect 7983 19558 7995 19610
rect 8047 19558 8059 19610
rect 8111 19558 11230 19610
rect 11282 19558 11294 19610
rect 11346 19558 11358 19610
rect 11410 19558 11422 19610
rect 11474 19558 11486 19610
rect 11538 19558 14657 19610
rect 14709 19558 14721 19610
rect 14773 19558 14785 19610
rect 14837 19558 14849 19610
rect 14901 19558 14913 19610
rect 14965 19558 14971 19610
rect 1104 19536 14971 19558
rect 2501 19499 2559 19505
rect 2501 19465 2513 19499
rect 2547 19496 2559 19499
rect 3970 19496 3976 19508
rect 2547 19468 3976 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4062 19456 4068 19508
rect 4120 19456 4126 19508
rect 4525 19499 4583 19505
rect 4525 19465 4537 19499
rect 4571 19496 4583 19499
rect 4890 19496 4896 19508
rect 4571 19468 4896 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 6086 19456 6092 19508
rect 6144 19456 6150 19508
rect 6914 19456 6920 19508
rect 6972 19456 6978 19508
rect 7006 19456 7012 19508
rect 7064 19456 7070 19508
rect 7193 19499 7251 19505
rect 7193 19465 7205 19499
rect 7239 19465 7251 19499
rect 7193 19459 7251 19465
rect 2774 19428 2780 19440
rect 2608 19400 2780 19428
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 2608 19369 2636 19400
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 3326 19388 3332 19440
rect 3384 19428 3390 19440
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 3384 19400 3801 19428
rect 3384 19388 3390 19400
rect 3789 19397 3801 19400
rect 3835 19397 3847 19431
rect 4080 19428 4108 19456
rect 5261 19431 5319 19437
rect 5261 19428 5273 19431
rect 4080 19400 5273 19428
rect 3789 19391 3847 19397
rect 5261 19397 5273 19400
rect 5307 19397 5319 19431
rect 6932 19428 6960 19456
rect 7208 19428 7236 19459
rect 7650 19456 7656 19508
rect 7708 19456 7714 19508
rect 7929 19499 7987 19505
rect 7929 19465 7941 19499
rect 7975 19496 7987 19499
rect 8478 19496 8484 19508
rect 7975 19468 8484 19496
rect 7975 19465 7987 19468
rect 7929 19459 7987 19465
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 9398 19456 9404 19508
rect 9456 19456 9462 19508
rect 9674 19456 9680 19508
rect 9732 19456 9738 19508
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10686 19496 10692 19508
rect 9824 19468 10692 19496
rect 9824 19456 9830 19468
rect 10686 19456 10692 19468
rect 10744 19496 10750 19508
rect 11514 19496 11520 19508
rect 10744 19468 11520 19496
rect 10744 19456 10750 19468
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 12345 19499 12403 19505
rect 12345 19496 12357 19499
rect 11756 19468 12357 19496
rect 11756 19456 11762 19468
rect 12345 19465 12357 19468
rect 12391 19465 12403 19499
rect 12345 19459 12403 19465
rect 12618 19456 12624 19508
rect 12676 19456 12682 19508
rect 13262 19456 13268 19508
rect 13320 19456 13326 19508
rect 13998 19456 14004 19508
rect 14056 19456 14062 19508
rect 14182 19456 14188 19508
rect 14240 19456 14246 19508
rect 14550 19456 14556 19508
rect 14608 19456 14614 19508
rect 8294 19428 8300 19440
rect 5261 19391 5319 19397
rect 5644 19400 6868 19428
rect 6932 19400 7236 19428
rect 7300 19400 8300 19428
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 2593 19363 2651 19369
rect 2593 19360 2605 19363
rect 2363 19332 2605 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 2593 19329 2605 19332
rect 2639 19329 2651 19363
rect 2593 19323 2651 19329
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 3053 19363 3111 19369
rect 3053 19360 3065 19363
rect 2731 19332 3065 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 3053 19329 3065 19332
rect 3099 19329 3111 19363
rect 3053 19323 3111 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5169 19363 5227 19369
rect 4764 19332 5028 19360
rect 4764 19320 4770 19332
rect 2406 19252 2412 19304
rect 2464 19292 2470 19304
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2464 19264 2881 19292
rect 2464 19252 2470 19264
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 3697 19295 3755 19301
rect 3697 19292 3709 19295
rect 3568 19264 3709 19292
rect 3568 19252 3574 19264
rect 3697 19261 3709 19264
rect 3743 19261 3755 19295
rect 3697 19255 3755 19261
rect 4338 19252 4344 19304
rect 4396 19292 4402 19304
rect 4890 19292 4896 19304
rect 4396 19264 4896 19292
rect 4396 19252 4402 19264
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5000 19301 5028 19332
rect 5169 19329 5181 19363
rect 5215 19360 5227 19363
rect 5644 19360 5672 19400
rect 5215 19332 5672 19360
rect 5215 19329 5227 19332
rect 5169 19323 5227 19329
rect 5718 19320 5724 19372
rect 5776 19360 5782 19372
rect 5997 19363 6055 19369
rect 5997 19360 6009 19363
rect 5776 19332 6009 19360
rect 5776 19320 5782 19332
rect 5997 19329 6009 19332
rect 6043 19329 6055 19363
rect 6840 19360 6868 19400
rect 7300 19360 7328 19400
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 9858 19428 9864 19440
rect 8628 19400 8892 19428
rect 8628 19388 8634 19400
rect 5997 19323 6055 19329
rect 6288 19332 6500 19360
rect 6840 19332 7328 19360
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19261 5043 19295
rect 5905 19295 5963 19301
rect 5905 19292 5917 19295
rect 4985 19255 5043 19261
rect 5092 19264 5917 19292
rect 2222 19184 2228 19236
rect 2280 19224 2286 19236
rect 3602 19224 3608 19236
rect 2280 19196 3608 19224
rect 2280 19184 2286 19196
rect 3602 19184 3608 19196
rect 3660 19224 3666 19236
rect 5092 19224 5120 19264
rect 5905 19261 5917 19264
rect 5951 19292 5963 19295
rect 6288 19292 6316 19332
rect 5951 19264 6316 19292
rect 6365 19295 6423 19301
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 6365 19261 6377 19295
rect 6411 19261 6423 19295
rect 6472 19292 6500 19332
rect 7374 19320 7380 19372
rect 7432 19320 7438 19372
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19360 7803 19363
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 7791 19332 8033 19360
rect 7791 19329 7803 19332
rect 7745 19323 7803 19329
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8159 19332 8800 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 6546 19292 6552 19304
rect 6472 19264 6552 19292
rect 6365 19255 6423 19261
rect 6380 19224 6408 19255
rect 6546 19252 6552 19264
rect 6604 19292 6610 19304
rect 7558 19292 7564 19304
rect 6604 19264 7564 19292
rect 6604 19252 6610 19264
rect 7558 19252 7564 19264
rect 7616 19292 7622 19304
rect 7760 19292 7788 19323
rect 8772 19301 8800 19332
rect 7616 19264 7788 19292
rect 8757 19295 8815 19301
rect 7616 19252 7622 19264
rect 8757 19261 8769 19295
rect 8803 19261 8815 19295
rect 8864 19292 8892 19400
rect 8956 19400 9864 19428
rect 8956 19369 8984 19400
rect 9858 19388 9864 19400
rect 9916 19388 9922 19440
rect 10134 19388 10140 19440
rect 10192 19428 10198 19440
rect 10505 19431 10563 19437
rect 10192 19400 10364 19428
rect 10192 19388 10198 19400
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 9214 19320 9220 19372
rect 9272 19320 9278 19372
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 10336 19360 10364 19400
rect 10505 19397 10517 19431
rect 10551 19428 10563 19431
rect 11606 19428 11612 19440
rect 10551 19400 11612 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 12636 19428 12664 19456
rect 14568 19428 14596 19456
rect 12124 19400 12664 19428
rect 14016 19400 14596 19428
rect 12124 19388 12130 19400
rect 14016 19372 14044 19400
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 9493 19323 9551 19329
rect 9876 19332 10180 19360
rect 10336 19332 10609 19360
rect 9508 19292 9536 19323
rect 9876 19301 9904 19332
rect 10152 19304 10180 19332
rect 10597 19329 10609 19332
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 8864 19264 9536 19292
rect 9861 19295 9919 19301
rect 8757 19255 8815 19261
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 10042 19252 10048 19304
rect 10100 19252 10106 19304
rect 10134 19252 10140 19304
rect 10192 19252 10198 19304
rect 10410 19252 10416 19304
rect 10468 19292 10474 19304
rect 10612 19292 10640 19323
rect 10468 19264 10640 19292
rect 10980 19292 11008 19323
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11112 19332 11529 19360
rect 11112 19320 11118 19332
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 12250 19360 12256 19372
rect 11517 19323 11575 19329
rect 11624 19332 12256 19360
rect 11624 19292 11652 19332
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12400 19332 12449 19360
rect 12400 19320 12406 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 13354 19320 13360 19372
rect 13412 19320 13418 19372
rect 13998 19320 14004 19372
rect 14056 19320 14062 19372
rect 14093 19363 14151 19369
rect 14093 19329 14105 19363
rect 14139 19360 14151 19363
rect 14550 19360 14556 19372
rect 14139 19332 14556 19360
rect 14139 19329 14151 19332
rect 14093 19323 14151 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 10980 19264 11652 19292
rect 11701 19295 11759 19301
rect 10468 19252 10474 19264
rect 11701 19261 11713 19295
rect 11747 19261 11759 19295
rect 11701 19255 11759 19261
rect 7834 19224 7840 19236
rect 3660 19196 5120 19224
rect 5920 19196 7840 19224
rect 3660 19184 3666 19196
rect 5920 19168 5948 19196
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 11149 19227 11207 19233
rect 7984 19196 10824 19224
rect 7984 19184 7990 19196
rect 934 19116 940 19168
rect 992 19156 998 19168
rect 1489 19159 1547 19165
rect 1489 19156 1501 19159
rect 992 19128 1501 19156
rect 992 19116 998 19128
rect 1489 19125 1501 19128
rect 1535 19125 1547 19159
rect 1489 19119 1547 19125
rect 2130 19116 2136 19168
rect 2188 19116 2194 19168
rect 5902 19116 5908 19168
rect 5960 19116 5966 19168
rect 7852 19156 7880 19184
rect 8294 19156 8300 19168
rect 7852 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 8938 19156 8944 19168
rect 8444 19128 8944 19156
rect 8444 19116 8450 19128
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 10686 19116 10692 19168
rect 10744 19116 10750 19168
rect 10796 19156 10824 19196
rect 11149 19193 11161 19227
rect 11195 19224 11207 19227
rect 11716 19224 11744 19255
rect 11882 19252 11888 19304
rect 11940 19292 11946 19304
rect 12805 19295 12863 19301
rect 11940 19264 12572 19292
rect 11940 19252 11946 19264
rect 12544 19224 12572 19264
rect 12805 19261 12817 19295
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 12820 19224 12848 19255
rect 11195 19196 11744 19224
rect 11808 19196 12434 19224
rect 12544 19196 12848 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 11808 19156 11836 19196
rect 10796 19128 11836 19156
rect 12158 19116 12164 19168
rect 12216 19116 12222 19168
rect 12406 19156 12434 19196
rect 13556 19156 13584 19255
rect 12406 19128 13584 19156
rect 1104 19066 14812 19088
rect 1104 19014 2663 19066
rect 2715 19014 2727 19066
rect 2779 19014 2791 19066
rect 2843 19014 2855 19066
rect 2907 19014 2919 19066
rect 2971 19014 6090 19066
rect 6142 19014 6154 19066
rect 6206 19014 6218 19066
rect 6270 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 9517 19066
rect 9569 19014 9581 19066
rect 9633 19014 9645 19066
rect 9697 19014 9709 19066
rect 9761 19014 9773 19066
rect 9825 19014 12944 19066
rect 12996 19014 13008 19066
rect 13060 19014 13072 19066
rect 13124 19014 13136 19066
rect 13188 19014 13200 19066
rect 13252 19014 14812 19066
rect 1104 18992 14812 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 1946 18952 1952 18964
rect 1627 18924 1952 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 2038 18912 2044 18964
rect 2096 18912 2102 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3510 18952 3516 18964
rect 3467 18924 3516 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 4154 18912 4160 18964
rect 4212 18912 4218 18964
rect 4430 18912 4436 18964
rect 4488 18912 4494 18964
rect 8386 18952 8392 18964
rect 4724 18924 8392 18952
rect 2056 18884 2084 18912
rect 4617 18887 4675 18893
rect 4617 18884 4629 18887
rect 2056 18856 4629 18884
rect 4617 18853 4629 18856
rect 4663 18853 4675 18887
rect 4617 18847 4675 18853
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18816 2099 18819
rect 2314 18816 2320 18828
rect 2087 18788 2320 18816
rect 2087 18785 2099 18788
rect 2041 18779 2099 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 3418 18776 3424 18828
rect 3476 18816 3482 18828
rect 3476 18788 4292 18816
rect 3476 18776 3482 18788
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1412 18680 1440 18711
rect 1854 18708 1860 18760
rect 1912 18708 1918 18760
rect 2222 18708 2228 18760
rect 2280 18708 2286 18760
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3786 18748 3792 18760
rect 3007 18720 3792 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 2240 18680 2268 18708
rect 1412 18652 2268 18680
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2501 18615 2559 18621
rect 2501 18612 2513 18615
rect 2372 18584 2513 18612
rect 2372 18572 2378 18584
rect 2501 18581 2513 18584
rect 2547 18612 2559 18615
rect 2792 18612 2820 18711
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4264 18757 4292 18788
rect 4724 18757 4752 18924
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9677 18955 9735 18961
rect 8496 18924 8892 18952
rect 4985 18887 5043 18893
rect 4985 18853 4997 18887
rect 5031 18853 5043 18887
rect 4985 18847 5043 18853
rect 5261 18887 5319 18893
rect 5261 18853 5273 18887
rect 5307 18884 5319 18887
rect 7561 18887 7619 18893
rect 5307 18856 5580 18884
rect 5307 18853 5319 18856
rect 5261 18847 5319 18853
rect 3973 18751 4031 18757
rect 3973 18748 3985 18751
rect 3936 18720 3985 18748
rect 3936 18708 3942 18720
rect 3973 18717 3985 18720
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18717 4307 18751
rect 4249 18711 4307 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18717 4859 18751
rect 5000 18748 5028 18847
rect 5552 18825 5580 18856
rect 7561 18853 7573 18887
rect 7607 18853 7619 18887
rect 7561 18847 7619 18853
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18785 5595 18819
rect 5537 18779 5595 18785
rect 5626 18776 5632 18828
rect 5684 18816 5690 18828
rect 6181 18819 6239 18825
rect 6181 18816 6193 18819
rect 5684 18788 6193 18816
rect 5684 18776 5690 18788
rect 6181 18785 6193 18788
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 7576 18816 7604 18847
rect 7926 18844 7932 18896
rect 7984 18844 7990 18896
rect 8496 18893 8524 18924
rect 8205 18887 8263 18893
rect 8205 18853 8217 18887
rect 8251 18884 8263 18887
rect 8481 18887 8539 18893
rect 8251 18856 8432 18884
rect 8251 18853 8263 18856
rect 8205 18847 8263 18853
rect 8110 18816 8116 18828
rect 6696 18788 6960 18816
rect 7576 18788 8116 18816
rect 6696 18776 6702 18788
rect 5077 18751 5135 18757
rect 5077 18748 5089 18751
rect 5000 18720 5089 18748
rect 4801 18711 4859 18717
rect 5077 18717 5089 18720
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5644 18748 5672 18776
rect 6932 18757 6960 18788
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 5399 18720 5672 18748
rect 6917 18751 6975 18757
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 6917 18717 6929 18751
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 7239 18720 7481 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7469 18717 7481 18720
rect 7515 18748 7527 18751
rect 7558 18748 7564 18760
rect 7515 18720 7564 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 4816 18680 4844 18711
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7650 18708 7656 18760
rect 7708 18748 7714 18760
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 7708 18720 7757 18748
rect 7708 18708 7714 18720
rect 7745 18717 7757 18720
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 7834 18708 7840 18760
rect 7892 18748 7898 18760
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7892 18720 8033 18748
rect 7892 18708 7898 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18750 8355 18751
rect 8404 18750 8432 18856
rect 8481 18853 8493 18887
rect 8527 18853 8539 18887
rect 8481 18847 8539 18853
rect 8570 18844 8576 18896
rect 8628 18844 8634 18896
rect 8580 18757 8608 18844
rect 8864 18816 8892 18924
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 9858 18952 9864 18964
rect 9723 18924 9864 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 9858 18912 9864 18924
rect 9916 18952 9922 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 9916 18924 10517 18952
rect 9916 18912 9922 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 11606 18912 11612 18964
rect 11664 18912 11670 18964
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12342 18952 12348 18964
rect 12216 18924 12348 18952
rect 12216 18912 12222 18924
rect 12342 18912 12348 18924
rect 12400 18952 12406 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 12400 18924 12449 18952
rect 12400 18912 12406 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 12437 18915 12495 18921
rect 12710 18912 12716 18964
rect 12768 18952 12774 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12768 18924 13001 18952
rect 12768 18912 12774 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 13817 18955 13875 18961
rect 13817 18921 13829 18955
rect 13863 18952 13875 18955
rect 13906 18952 13912 18964
rect 13863 18924 13912 18952
rect 13863 18921 13875 18924
rect 13817 18915 13875 18921
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 8938 18844 8944 18896
rect 8996 18884 9002 18896
rect 8996 18856 11560 18884
rect 8996 18844 9002 18856
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 8864 18788 9229 18816
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 10134 18816 10140 18828
rect 9217 18779 9275 18785
rect 9692 18788 10140 18816
rect 9692 18760 9720 18788
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 10318 18776 10324 18828
rect 10376 18776 10382 18828
rect 10686 18776 10692 18828
rect 10744 18816 10750 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 10744 18788 11437 18816
rect 10744 18776 10750 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 8343 18722 8432 18750
rect 8573 18751 8631 18757
rect 8343 18717 8355 18722
rect 8297 18711 8355 18717
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18748 8723 18751
rect 8938 18748 8944 18760
rect 8711 18720 8944 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9033 18751 9091 18757
rect 9033 18717 9045 18751
rect 9079 18748 9091 18751
rect 9674 18748 9680 18760
rect 9079 18720 9680 18748
rect 9079 18717 9091 18720
rect 9033 18711 9091 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 10336 18748 10364 18776
rect 9907 18720 10364 18748
rect 10413 18751 10471 18757
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 10594 18748 10600 18760
rect 10459 18720 10600 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10962 18708 10968 18760
rect 11020 18708 11026 18760
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 11112 18720 11161 18748
rect 11112 18708 11118 18720
rect 11149 18717 11161 18720
rect 11195 18748 11207 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 11195 18720 11253 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11532 18748 11560 18856
rect 11624 18816 11652 18912
rect 14090 18884 14096 18896
rect 12084 18856 14096 18884
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11624 18788 11989 18816
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12084 18748 12112 18856
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 11532 18720 12112 18748
rect 11241 18711 11299 18717
rect 12158 18708 12164 18760
rect 12216 18708 12222 18760
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 13722 18748 13728 18760
rect 13587 18720 13728 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18748 14151 18751
rect 15194 18748 15200 18760
rect 14139 18720 15200 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 5534 18680 5540 18692
rect 4816 18652 5540 18680
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 6270 18640 6276 18692
rect 6328 18640 6334 18692
rect 6825 18683 6883 18689
rect 6825 18649 6837 18683
rect 6871 18680 6883 18683
rect 7282 18680 7288 18692
rect 6871 18652 7288 18680
rect 6871 18649 6883 18652
rect 6825 18643 6883 18649
rect 7282 18640 7288 18652
rect 7340 18640 7346 18692
rect 7392 18652 8156 18680
rect 2547 18584 2820 18612
rect 2547 18581 2559 18584
rect 2501 18575 2559 18581
rect 5994 18572 6000 18624
rect 6052 18572 6058 18624
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18612 7159 18615
rect 7190 18612 7196 18624
rect 7147 18584 7196 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 7392 18621 7420 18652
rect 7377 18615 7435 18621
rect 7377 18581 7389 18615
rect 7423 18581 7435 18615
rect 8128 18612 8156 18652
rect 8404 18652 12434 18680
rect 8404 18612 8432 18652
rect 8128 18584 8432 18612
rect 7377 18575 7435 18581
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 12066 18612 12072 18624
rect 8536 18584 12072 18612
rect 8536 18572 8542 18584
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12406 18612 12434 18652
rect 12894 18640 12900 18692
rect 12952 18640 12958 18692
rect 13372 18652 14504 18680
rect 13372 18612 13400 18652
rect 14476 18624 14504 18652
rect 12406 18584 13400 18612
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 14277 18615 14335 18621
rect 14277 18612 14289 18615
rect 14240 18584 14289 18612
rect 14240 18572 14246 18584
rect 14277 18581 14289 18584
rect 14323 18581 14335 18615
rect 14277 18575 14335 18581
rect 14458 18572 14464 18624
rect 14516 18572 14522 18624
rect 1104 18522 14971 18544
rect 1104 18470 4376 18522
rect 4428 18470 4440 18522
rect 4492 18470 4504 18522
rect 4556 18470 4568 18522
rect 4620 18470 4632 18522
rect 4684 18470 7803 18522
rect 7855 18470 7867 18522
rect 7919 18470 7931 18522
rect 7983 18470 7995 18522
rect 8047 18470 8059 18522
rect 8111 18470 11230 18522
rect 11282 18470 11294 18522
rect 11346 18470 11358 18522
rect 11410 18470 11422 18522
rect 11474 18470 11486 18522
rect 11538 18470 14657 18522
rect 14709 18470 14721 18522
rect 14773 18470 14785 18522
rect 14837 18470 14849 18522
rect 14901 18470 14913 18522
rect 14965 18470 14971 18522
rect 1104 18448 14971 18470
rect 2314 18368 2320 18420
rect 2372 18368 2378 18420
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18377 5135 18411
rect 5077 18371 5135 18377
rect 5353 18411 5411 18417
rect 5353 18377 5365 18411
rect 5399 18408 5411 18411
rect 5399 18380 7420 18408
rect 5399 18377 5411 18380
rect 5353 18371 5411 18377
rect 3620 18340 3648 18368
rect 3344 18312 3648 18340
rect 5092 18340 5120 18371
rect 6270 18340 6276 18352
rect 5092 18312 6276 18340
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1857 18275 1915 18281
rect 1857 18272 1869 18275
rect 1636 18244 1869 18272
rect 1636 18232 1642 18244
rect 1857 18241 1869 18244
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 3344 18281 3372 18312
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 6454 18300 6460 18352
rect 6512 18300 6518 18352
rect 6546 18300 6552 18352
rect 6604 18300 6610 18352
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7248 18312 7328 18340
rect 7248 18300 7254 18312
rect 2593 18275 2651 18281
rect 2593 18272 2605 18275
rect 2188 18244 2605 18272
rect 2188 18232 2194 18244
rect 2593 18241 2605 18244
rect 2639 18241 2651 18275
rect 2593 18235 2651 18241
rect 3329 18275 3387 18281
rect 3329 18241 3341 18275
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 3510 18232 3516 18284
rect 3568 18272 3574 18284
rect 3677 18275 3735 18281
rect 3677 18272 3689 18275
rect 3568 18244 3689 18272
rect 3568 18232 3574 18244
rect 3677 18241 3689 18244
rect 3723 18241 3735 18275
rect 3677 18235 3735 18241
rect 4890 18232 4896 18284
rect 4948 18232 4954 18284
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18272 5319 18275
rect 5534 18272 5540 18284
rect 5307 18244 5540 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 5534 18232 5540 18244
rect 5592 18272 5598 18284
rect 6089 18275 6147 18281
rect 6089 18272 6101 18275
rect 5592 18244 6101 18272
rect 5592 18232 5598 18244
rect 6089 18241 6101 18244
rect 6135 18241 6147 18275
rect 6089 18235 6147 18241
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 2222 18204 2228 18216
rect 1719 18176 2228 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2455 18176 2774 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2746 18136 2774 18176
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3292 18176 3433 18204
rect 3292 18164 3298 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 2746 18108 3372 18136
rect 3344 18080 3372 18108
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 2406 18028 2412 18080
rect 2464 18068 2470 18080
rect 2777 18071 2835 18077
rect 2777 18068 2789 18071
rect 2464 18040 2789 18068
rect 2464 18028 2470 18040
rect 2777 18037 2789 18040
rect 2823 18037 2835 18071
rect 2777 18031 2835 18037
rect 3234 18028 3240 18080
rect 3292 18028 3298 18080
rect 3326 18028 3332 18080
rect 3384 18028 3390 18080
rect 3436 18068 3464 18167
rect 5994 18164 6000 18216
rect 6052 18164 6058 18216
rect 6454 18164 6460 18216
rect 6512 18204 6518 18216
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6512 18176 7205 18204
rect 6512 18164 6518 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7300 18204 7328 18312
rect 7392 18281 7420 18380
rect 8294 18368 8300 18420
rect 8352 18368 8358 18420
rect 8757 18411 8815 18417
rect 8757 18377 8769 18411
rect 8803 18408 8815 18411
rect 10962 18408 10968 18420
rect 8803 18380 10968 18408
rect 8803 18377 8815 18380
rect 8757 18371 8815 18377
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 12158 18408 12164 18420
rect 11655 18380 12164 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 12268 18380 14136 18408
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8312 18272 8340 18368
rect 8938 18300 8944 18352
rect 8996 18340 9002 18352
rect 11054 18340 11060 18352
rect 8996 18312 11060 18340
rect 8996 18300 9002 18312
rect 8389 18275 8447 18281
rect 8389 18272 8401 18275
rect 8159 18244 8248 18272
rect 8312 18244 8401 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 7300 18176 8156 18204
rect 7193 18167 7251 18173
rect 4801 18139 4859 18145
rect 4801 18105 4813 18139
rect 4847 18136 4859 18139
rect 5902 18136 5908 18148
rect 4847 18108 5908 18136
rect 4847 18105 4859 18108
rect 4801 18099 4859 18105
rect 5902 18096 5908 18108
rect 5960 18096 5966 18148
rect 4062 18068 4068 18080
rect 3436 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 5534 18028 5540 18080
rect 5592 18028 5598 18080
rect 6012 18068 6040 18164
rect 8128 18148 8156 18176
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 7282 18136 7288 18148
rect 7055 18108 7288 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 7282 18096 7288 18108
rect 7340 18096 7346 18148
rect 8110 18096 8116 18148
rect 8168 18096 8174 18148
rect 8220 18145 8248 18244
rect 8389 18241 8401 18244
rect 8435 18272 8447 18275
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8435 18244 8677 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18272 9183 18275
rect 9214 18272 9220 18284
rect 9171 18244 9220 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9214 18232 9220 18244
rect 9272 18232 9278 18284
rect 9968 18281 9996 18312
rect 11054 18300 11060 18312
rect 11112 18300 11118 18352
rect 12268 18340 12296 18380
rect 11164 18312 12296 18340
rect 12360 18312 12480 18340
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9416 18244 9597 18272
rect 9416 18216 9444 18244
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 10410 18272 10416 18284
rect 9953 18235 10011 18241
rect 10060 18244 10416 18272
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 10060 18204 10088 18244
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 9456 18176 10088 18204
rect 9456 18164 9462 18176
rect 10134 18164 10140 18216
rect 10192 18164 10198 18216
rect 10318 18164 10324 18216
rect 10376 18204 10382 18216
rect 10612 18204 10640 18232
rect 10376 18176 10640 18204
rect 10689 18207 10747 18213
rect 10376 18164 10382 18176
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18105 8263 18139
rect 8205 18099 8263 18105
rect 9217 18139 9275 18145
rect 9217 18105 9229 18139
rect 9263 18136 9275 18139
rect 9674 18136 9680 18148
rect 9263 18108 9680 18136
rect 9263 18105 9275 18108
rect 9217 18099 9275 18105
rect 9674 18096 9680 18108
rect 9732 18136 9738 18148
rect 10704 18136 10732 18167
rect 10870 18164 10876 18216
rect 10928 18164 10934 18216
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11164 18204 11192 18312
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11563 18244 11652 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11624 18216 11652 18244
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 12158 18272 12164 18284
rect 11756 18244 12164 18272
rect 11756 18232 11762 18244
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12360 18272 12388 18312
rect 12452 18281 12480 18312
rect 13906 18300 13912 18352
rect 13964 18300 13970 18352
rect 14108 18349 14136 18380
rect 14093 18343 14151 18349
rect 14093 18309 14105 18343
rect 14139 18309 14151 18343
rect 14093 18303 14151 18309
rect 12268 18244 12388 18272
rect 12437 18275 12495 18281
rect 11112 18176 11192 18204
rect 11112 18164 11118 18176
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 12268 18204 12296 18244
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 12584 18244 13553 18272
rect 12584 18232 12590 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 11664 18176 12296 18204
rect 11664 18164 11670 18176
rect 12342 18164 12348 18216
rect 12400 18204 12406 18216
rect 12713 18207 12771 18213
rect 12713 18204 12725 18207
rect 12400 18176 12725 18204
rect 12400 18164 12406 18176
rect 12713 18173 12725 18176
rect 12759 18173 12771 18207
rect 12713 18167 12771 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13446 18204 13452 18216
rect 12943 18176 13452 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 9732 18108 10732 18136
rect 9732 18096 9738 18108
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 11882 18136 11888 18148
rect 11020 18108 11888 18136
rect 11020 18096 11026 18108
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 12250 18096 12256 18148
rect 12308 18096 12314 18148
rect 6822 18068 6828 18080
rect 6012 18040 6828 18068
rect 6822 18028 6828 18040
rect 6880 18068 6886 18080
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 6880 18040 7573 18068
rect 6880 18028 6886 18040
rect 7561 18037 7573 18040
rect 7607 18037 7619 18071
rect 7561 18031 7619 18037
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 8018 18068 8024 18080
rect 7975 18040 8024 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 9858 18068 9864 18080
rect 9815 18040 9864 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 10643 18040 11345 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 11333 18037 11345 18040
rect 11379 18068 11391 18071
rect 11698 18068 11704 18080
rect 11379 18040 11704 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12066 18028 12072 18080
rect 12124 18028 12130 18080
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 14458 18068 14464 18080
rect 14415 18040 14464 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 1104 17978 14812 18000
rect 1104 17926 2663 17978
rect 2715 17926 2727 17978
rect 2779 17926 2791 17978
rect 2843 17926 2855 17978
rect 2907 17926 2919 17978
rect 2971 17926 6090 17978
rect 6142 17926 6154 17978
rect 6206 17926 6218 17978
rect 6270 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 9517 17978
rect 9569 17926 9581 17978
rect 9633 17926 9645 17978
rect 9697 17926 9709 17978
rect 9761 17926 9773 17978
rect 9825 17926 12944 17978
rect 12996 17926 13008 17978
rect 13060 17926 13072 17978
rect 13124 17926 13136 17978
rect 13188 17926 13200 17978
rect 13252 17926 14812 17978
rect 1104 17904 14812 17926
rect 2406 17824 2412 17876
rect 2464 17824 2470 17876
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 3878 17864 3884 17876
rect 3384 17836 3884 17864
rect 3384 17824 3390 17836
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 7650 17824 7656 17876
rect 7708 17824 7714 17876
rect 8570 17824 8576 17876
rect 8628 17824 8634 17876
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 9401 17867 9459 17873
rect 9401 17864 9413 17867
rect 9364 17836 9413 17864
rect 9364 17824 9370 17836
rect 9401 17833 9413 17836
rect 9447 17833 9459 17867
rect 9401 17827 9459 17833
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10042 17864 10048 17876
rect 9999 17836 10048 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10192 17836 10701 17864
rect 10192 17824 10198 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 10870 17824 10876 17876
rect 10928 17824 10934 17876
rect 12529 17867 12587 17873
rect 11348 17836 12434 17864
rect 7101 17799 7159 17805
rect 7101 17765 7113 17799
rect 7147 17765 7159 17799
rect 7668 17796 7696 17824
rect 9493 17799 9551 17805
rect 9493 17796 9505 17799
rect 7668 17768 9505 17796
rect 7101 17759 7159 17765
rect 9493 17765 9505 17768
rect 9539 17765 9551 17799
rect 10226 17796 10232 17808
rect 9493 17759 9551 17765
rect 9600 17768 10232 17796
rect 2593 17731 2651 17737
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 3234 17728 3240 17740
rect 2639 17700 3240 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 4172 17700 5181 17728
rect 4172 17672 4200 17700
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 7116 17728 7144 17759
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7116 17700 7389 17728
rect 5169 17691 5227 17697
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 8294 17728 8300 17740
rect 7975 17700 8300 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 992 17632 1409 17660
rect 992 17620 998 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 2866 17660 2872 17672
rect 2823 17632 2872 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3881 17663 3939 17669
rect 3881 17660 3893 17663
rect 3620 17632 3893 17660
rect 1762 17552 1768 17604
rect 1820 17552 1826 17604
rect 3620 17536 3648 17632
rect 3881 17629 3893 17632
rect 3927 17629 3939 17663
rect 3881 17623 3939 17629
rect 4154 17620 4160 17672
rect 4212 17620 4218 17672
rect 4798 17620 4804 17672
rect 4856 17620 4862 17672
rect 6914 17620 6920 17672
rect 6972 17620 6978 17672
rect 7098 17620 7104 17672
rect 7156 17660 7162 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 7156 17632 7205 17660
rect 7156 17620 7162 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 8018 17620 8024 17672
rect 8076 17660 8082 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 8076 17632 8125 17660
rect 8076 17620 8082 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 8113 17623 8171 17629
rect 8680 17632 8953 17660
rect 5436 17595 5494 17601
rect 5436 17561 5448 17595
rect 5482 17592 5494 17595
rect 5534 17592 5540 17604
rect 5482 17564 5540 17592
rect 5482 17561 5494 17564
rect 5436 17555 5494 17561
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 8680 17536 8708 17632
rect 8941 17629 8953 17632
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17660 9275 17663
rect 9600 17660 9628 17768
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 11348 17805 11376 17836
rect 10505 17799 10563 17805
rect 10505 17765 10517 17799
rect 10551 17765 10563 17799
rect 10505 17759 10563 17765
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17765 11391 17799
rect 11333 17759 11391 17765
rect 11425 17799 11483 17805
rect 11425 17765 11437 17799
rect 11471 17765 11483 17799
rect 11425 17759 11483 17765
rect 10520 17728 10548 17759
rect 10520 17700 11100 17728
rect 9263 17632 9628 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 9674 17620 9680 17672
rect 9732 17620 9738 17672
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10042 17620 10048 17672
rect 10100 17620 10106 17672
rect 11072 17669 11100 17700
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 10367 17656 10456 17660
rect 10612 17656 10793 17660
rect 10367 17632 10793 17656
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 10428 17628 10640 17632
rect 10134 17592 10140 17604
rect 9140 17564 10140 17592
rect 2869 17527 2927 17533
rect 2869 17493 2881 17527
rect 2915 17524 2927 17527
rect 2958 17524 2964 17536
rect 2915 17496 2964 17524
rect 2915 17493 2927 17496
rect 2869 17487 2927 17493
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 3602 17484 3608 17536
rect 3660 17484 3666 17536
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 3973 17527 4031 17533
rect 3973 17524 3985 17527
rect 3936 17496 3985 17524
rect 3936 17484 3942 17496
rect 3973 17493 3985 17496
rect 4019 17493 4031 17527
rect 3973 17487 4031 17493
rect 4246 17484 4252 17536
rect 4304 17484 4310 17536
rect 6549 17527 6607 17533
rect 6549 17493 6561 17527
rect 6595 17524 6607 17527
rect 7006 17524 7012 17536
rect 6595 17496 7012 17524
rect 6595 17493 6607 17496
rect 6549 17487 6607 17493
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7248 17496 7849 17524
rect 7248 17484 7254 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 8662 17484 8668 17536
rect 8720 17484 8726 17536
rect 9140 17533 9168 17564
rect 10134 17552 10140 17564
rect 10192 17552 10198 17604
rect 10704 17536 10732 17632
rect 10781 17629 10793 17632
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 11440 17660 11468 17759
rect 11624 17700 12020 17728
rect 11624 17669 11652 17700
rect 11195 17632 11468 17660
rect 11609 17663 11667 17669
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 11609 17629 11621 17663
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 11882 17620 11888 17672
rect 11940 17620 11946 17672
rect 11992 17660 12020 17700
rect 12066 17688 12072 17740
rect 12124 17688 12130 17740
rect 12406 17728 12434 17836
rect 12529 17833 12541 17867
rect 12575 17864 12587 17867
rect 12618 17864 12624 17876
rect 12575 17836 12624 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 12618 17824 12624 17836
rect 12676 17864 12682 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12676 17836 13001 17864
rect 12676 17824 12682 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 13446 17824 13452 17876
rect 13504 17824 13510 17876
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 12406 17700 12817 17728
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 11992 17632 12112 17660
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 11974 17592 11980 17604
rect 10928 17564 11980 17592
rect 10928 17552 10934 17564
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12084 17592 12112 17632
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12400 17632 12633 17660
rect 12400 17620 12406 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 12621 17623 12679 17629
rect 13464 17632 13553 17660
rect 12158 17592 12164 17604
rect 12084 17564 12164 17592
rect 12158 17552 12164 17564
rect 12216 17592 12222 17604
rect 12216 17564 12434 17592
rect 12216 17552 12222 17564
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17493 9183 17527
rect 9125 17487 9183 17493
rect 10226 17484 10232 17536
rect 10284 17484 10290 17536
rect 10686 17484 10692 17536
rect 10744 17484 10750 17536
rect 12406 17524 12434 17564
rect 13464 17536 13492 17632
rect 13541 17629 13553 17632
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 13630 17620 13636 17672
rect 13688 17620 13694 17672
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14056 17632 14289 17660
rect 14056 17620 14062 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 12710 17524 12716 17536
rect 12406 17496 12716 17524
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 13722 17484 13728 17536
rect 13780 17484 13786 17536
rect 14090 17484 14096 17536
rect 14148 17484 14154 17536
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1452 17292 1961 17320
rect 1452 17280 1458 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 3418 17320 3424 17332
rect 1949 17283 2007 17289
rect 2424 17292 3424 17320
rect 2424 17196 2452 17292
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4246 17280 4252 17332
rect 4304 17280 4310 17332
rect 4890 17280 4896 17332
rect 4948 17320 4954 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 4948 17292 5733 17320
rect 4948 17280 4954 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 5721 17283 5779 17289
rect 6089 17323 6147 17329
rect 6089 17289 6101 17323
rect 6135 17320 6147 17323
rect 6546 17320 6552 17332
rect 6135 17292 6552 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7561 17323 7619 17329
rect 7561 17320 7573 17323
rect 6972 17292 7573 17320
rect 6972 17280 6978 17292
rect 7561 17289 7573 17292
rect 7607 17289 7619 17323
rect 7561 17283 7619 17289
rect 8849 17323 8907 17329
rect 8849 17289 8861 17323
rect 8895 17320 8907 17323
rect 9122 17320 9128 17332
rect 8895 17292 9128 17320
rect 8895 17289 8907 17292
rect 8849 17283 8907 17289
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9968 17292 11928 17320
rect 4264 17252 4292 17280
rect 4402 17255 4460 17261
rect 4402 17252 4414 17255
rect 2700 17224 4200 17252
rect 4264 17224 4414 17252
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 2130 17144 2136 17196
rect 2188 17144 2194 17196
rect 2406 17144 2412 17196
rect 2464 17144 2470 17196
rect 2700 17193 2728 17224
rect 2958 17193 2964 17196
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17153 2743 17187
rect 2952 17184 2964 17193
rect 2919 17156 2964 17184
rect 2685 17147 2743 17153
rect 2952 17147 2964 17156
rect 2958 17144 2964 17147
rect 3016 17144 3022 17196
rect 4172 17128 4200 17224
rect 4402 17221 4414 17224
rect 4448 17221 4460 17255
rect 4402 17215 4460 17221
rect 7098 17212 7104 17264
rect 7156 17252 7162 17264
rect 9861 17255 9919 17261
rect 9861 17252 9873 17255
rect 7156 17224 9873 17252
rect 7156 17212 7162 17224
rect 9861 17221 9873 17224
rect 9907 17221 9919 17255
rect 9861 17215 9919 17221
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 9968 17193 9996 17292
rect 10410 17212 10416 17264
rect 10468 17212 10474 17264
rect 10502 17212 10508 17264
rect 10560 17212 10566 17264
rect 10962 17212 10968 17264
rect 11020 17212 11026 17264
rect 11422 17252 11428 17264
rect 11072 17224 11428 17252
rect 5905 17187 5963 17193
rect 5905 17184 5917 17187
rect 5868 17156 5917 17184
rect 5868 17144 5874 17156
rect 5905 17153 5917 17156
rect 5951 17184 5963 17187
rect 5997 17187 6055 17193
rect 5997 17184 6009 17187
rect 5951 17156 6009 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 5997 17153 6009 17156
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17184 6699 17187
rect 7009 17187 7067 17193
rect 7009 17184 7021 17187
rect 6687 17156 7021 17184
rect 6687 17153 6699 17156
rect 6641 17147 6699 17153
rect 7009 17153 7021 17156
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 7745 17147 7803 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 7929 17147 7987 17153
rect 8128 17156 9137 17184
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 5537 17051 5595 17057
rect 5537 17017 5549 17051
rect 5583 17048 5595 17051
rect 5626 17048 5632 17060
rect 5583 17020 5632 17048
rect 5583 17017 5595 17020
rect 5537 17011 5595 17017
rect 5626 17008 5632 17020
rect 5684 17008 5690 17060
rect 6564 17048 6592 17147
rect 6822 17076 6828 17128
rect 6880 17076 6886 17128
rect 7760 17116 7788 17147
rect 6932 17088 7788 17116
rect 7944 17116 7972 17147
rect 8018 17116 8024 17128
rect 7944 17088 8024 17116
rect 6932 17048 6960 17088
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8128 17057 8156 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9953 17187 10011 17193
rect 9539 17156 9904 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8294 17116 8300 17128
rect 8251 17088 8300 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8435 17088 8984 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8956 17057 8984 17088
rect 6564 17020 6960 17048
rect 6932 16992 6960 17020
rect 8113 17051 8171 17057
rect 8113 17017 8125 17051
rect 8159 17017 8171 17051
rect 8113 17011 8171 17017
rect 8941 17051 8999 17057
rect 8941 17017 8953 17051
rect 8987 17017 8999 17051
rect 8941 17011 8999 17017
rect 934 16940 940 16992
rect 992 16980 998 16992
rect 1489 16983 1547 16989
rect 1489 16980 1501 16983
rect 992 16952 1501 16980
rect 992 16940 998 16952
rect 1489 16949 1501 16952
rect 1535 16949 1547 16983
rect 1489 16943 1547 16949
rect 2222 16940 2228 16992
rect 2280 16940 2286 16992
rect 4065 16983 4123 16989
rect 4065 16949 4077 16983
rect 4111 16980 4123 16983
rect 4798 16980 4804 16992
rect 4111 16952 4804 16980
rect 4111 16949 4123 16952
rect 4065 16943 4123 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 6914 16940 6920 16992
rect 6972 16940 6978 16992
rect 7190 16940 7196 16992
rect 7248 16940 7254 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 9508 16980 9536 17147
rect 9876 17128 9904 17156
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10520 17184 10548 17212
rect 10367 17156 10548 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 9858 17076 9864 17128
rect 9916 17076 9922 17128
rect 10060 17116 10088 17147
rect 10594 17144 10600 17196
rect 10652 17144 10658 17196
rect 10980 17184 11008 17212
rect 11072 17193 11100 17224
rect 11422 17212 11428 17224
rect 11480 17212 11486 17264
rect 11900 17252 11928 17292
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12434 17320 12440 17332
rect 12032 17292 12440 17320
rect 12032 17280 12038 17292
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13354 17280 13360 17332
rect 13412 17280 13418 17332
rect 13262 17252 13268 17264
rect 11900 17224 13268 17252
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 10704 17156 11008 17184
rect 11057 17187 11115 17193
rect 10502 17116 10508 17128
rect 10060 17088 10508 17116
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 9585 17051 9643 17057
rect 9585 17017 9597 17051
rect 9631 17048 9643 17051
rect 10704 17048 10732 17156
rect 11057 17153 11069 17187
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17153 11207 17187
rect 11514 17184 11520 17196
rect 11572 17193 11578 17196
rect 11483 17156 11520 17184
rect 11149 17147 11207 17153
rect 11164 17116 11192 17147
rect 11514 17144 11520 17156
rect 11572 17147 11583 17193
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17184 14243 17187
rect 14366 17184 14372 17196
rect 14231 17156 14372 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 11572 17144 11578 17147
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 10796 17088 11192 17116
rect 10796 17057 10824 17088
rect 11882 17076 11888 17128
rect 11940 17076 11946 17128
rect 12069 17119 12127 17125
rect 12069 17085 12081 17119
rect 12115 17116 12127 17119
rect 12158 17116 12164 17128
rect 12115 17088 12164 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12400 17088 12633 17116
rect 12400 17076 12406 17088
rect 9631 17020 10732 17048
rect 10781 17051 10839 17057
rect 9631 17017 9643 17020
rect 9585 17011 9643 17017
rect 10781 17017 10793 17051
rect 10827 17017 10839 17051
rect 10781 17011 10839 17017
rect 10870 17008 10876 17060
rect 10928 17008 10934 17060
rect 11054 17008 11060 17060
rect 11112 17008 11118 17060
rect 11974 17048 11980 17060
rect 11256 17020 11980 17048
rect 7616 16952 9536 16980
rect 10229 16983 10287 16989
rect 7616 16940 7622 16952
rect 10229 16949 10241 16983
rect 10275 16980 10287 16983
rect 11072 16980 11100 17008
rect 11256 16989 11284 17020
rect 11974 17008 11980 17020
rect 12032 17008 12038 17060
rect 12452 16992 12480 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12802 17076 12808 17128
rect 12860 17076 12866 17128
rect 13814 17076 13820 17128
rect 13872 17076 13878 17128
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 12529 17051 12587 17057
rect 12529 17017 12541 17051
rect 12575 17048 12587 17051
rect 12989 17051 13047 17057
rect 12989 17048 13001 17051
rect 12575 17020 13001 17048
rect 12575 17017 12587 17020
rect 12529 17011 12587 17017
rect 12989 17017 13001 17020
rect 13035 17048 13047 17051
rect 14016 17048 14044 17079
rect 13035 17020 14044 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 10275 16952 11100 16980
rect 11241 16983 11299 16989
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 11241 16949 11253 16983
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 11701 16983 11759 16989
rect 11701 16949 11713 16983
rect 11747 16980 11759 16983
rect 12342 16980 12348 16992
rect 11747 16952 12348 16980
rect 11747 16949 11759 16952
rect 11701 16943 11759 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12434 16940 12440 16992
rect 12492 16940 12498 16992
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 3878 16776 3884 16788
rect 3752 16748 3884 16776
rect 3752 16736 3758 16748
rect 3878 16736 3884 16748
rect 3936 16776 3942 16788
rect 7374 16776 7380 16788
rect 3936 16748 4476 16776
rect 3936 16736 3942 16748
rect 3142 16668 3148 16720
rect 3200 16708 3206 16720
rect 4062 16708 4068 16720
rect 3200 16680 4068 16708
rect 3200 16668 3206 16680
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 4154 16668 4160 16720
rect 4212 16668 4218 16720
rect 1578 16600 1584 16652
rect 1636 16600 1642 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 4172 16640 4200 16668
rect 2823 16612 4200 16640
rect 4341 16643 4399 16649
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 4341 16609 4353 16643
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 1596 16572 1624 16600
rect 2869 16575 2927 16581
rect 1596 16544 2820 16572
rect 2498 16464 2504 16516
rect 2556 16513 2562 16516
rect 2556 16467 2568 16513
rect 2792 16504 2820 16544
rect 2869 16541 2881 16575
rect 2915 16572 2927 16575
rect 2958 16572 2964 16584
rect 2915 16544 2964 16572
rect 2915 16541 2927 16544
rect 2869 16535 2927 16541
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3694 16572 3700 16584
rect 3053 16535 3111 16541
rect 3160 16544 3700 16572
rect 3068 16504 3096 16535
rect 2792 16476 3096 16504
rect 2556 16464 2562 16467
rect 1394 16396 1400 16448
rect 1452 16396 1458 16448
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3160 16436 3188 16544
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 3878 16532 3884 16584
rect 3936 16532 3942 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 3988 16544 4169 16572
rect 3513 16507 3571 16513
rect 3513 16473 3525 16507
rect 3559 16504 3571 16507
rect 3988 16504 4016 16544
rect 4157 16541 4169 16544
rect 4203 16572 4215 16575
rect 4246 16572 4252 16584
rect 4203 16544 4252 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 4356 16504 4384 16603
rect 3559 16476 4016 16504
rect 4080 16476 4384 16504
rect 4448 16504 4476 16748
rect 5644 16748 7380 16776
rect 5644 16652 5672 16748
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 9122 16736 9128 16788
rect 9180 16736 9186 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 12713 16779 12771 16785
rect 10284 16748 12434 16776
rect 10284 16736 10290 16748
rect 5721 16711 5779 16717
rect 5721 16677 5733 16711
rect 5767 16708 5779 16711
rect 9140 16708 9168 16736
rect 11241 16711 11299 16717
rect 5767 16680 6592 16708
rect 9140 16680 9260 16708
rect 5767 16677 5779 16680
rect 5721 16671 5779 16677
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 6564 16649 6592 16680
rect 6549 16643 6607 16649
rect 6288 16612 6500 16640
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4856 16544 4905 16572
rect 4856 16532 4862 16544
rect 4893 16541 4905 16544
rect 4939 16572 4951 16575
rect 5353 16575 5411 16581
rect 5353 16572 5365 16575
rect 4939 16544 5365 16572
rect 4939 16541 4951 16544
rect 4893 16535 4951 16541
rect 5353 16541 5365 16544
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 5644 16572 5672 16600
rect 6288 16581 6316 16612
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 5644 16544 5825 16572
rect 5537 16535 5595 16541
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 5552 16504 5580 16535
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 6472 16504 6500 16612
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 8018 16640 8024 16652
rect 7524 16612 8024 16640
rect 7524 16600 7530 16612
rect 8018 16600 8024 16612
rect 8076 16640 8082 16652
rect 8665 16643 8723 16649
rect 8076 16612 8340 16640
rect 8076 16600 8082 16612
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 7009 16575 7067 16581
rect 7009 16572 7021 16575
rect 6788 16544 7021 16572
rect 6788 16532 6794 16544
rect 7009 16541 7021 16544
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16541 7343 16575
rect 7285 16535 7343 16541
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8312 16572 8340 16612
rect 8665 16609 8677 16643
rect 8711 16640 8723 16643
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8711 16612 9137 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 8389 16575 8447 16581
rect 8389 16572 8401 16575
rect 8159 16544 8248 16572
rect 8312 16544 8401 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 6638 16504 6644 16516
rect 4448 16476 5304 16504
rect 5552 16476 6132 16504
rect 6472 16476 6644 16504
rect 3559 16473 3571 16476
rect 3513 16467 3571 16473
rect 4080 16445 4108 16476
rect 3016 16408 3188 16436
rect 4065 16439 4123 16445
rect 3016 16396 3022 16408
rect 4065 16405 4077 16439
rect 4111 16405 4123 16439
rect 4065 16399 4123 16405
rect 4706 16396 4712 16448
rect 4764 16436 4770 16448
rect 4801 16439 4859 16445
rect 4801 16436 4813 16439
rect 4764 16408 4813 16436
rect 4764 16396 4770 16408
rect 4801 16405 4813 16408
rect 4847 16405 4859 16439
rect 4801 16399 4859 16405
rect 4982 16396 4988 16448
rect 5040 16396 5046 16448
rect 5166 16396 5172 16448
rect 5224 16396 5230 16448
rect 5276 16436 5304 16476
rect 5718 16436 5724 16448
rect 5276 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16436 5963 16439
rect 5994 16436 6000 16448
rect 5951 16408 6000 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 6104 16445 6132 16476
rect 6638 16464 6644 16476
rect 6696 16504 6702 16516
rect 7300 16504 7328 16535
rect 6696 16476 7328 16504
rect 6696 16464 6702 16476
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16405 6147 16439
rect 6089 16399 6147 16405
rect 7374 16396 7380 16448
rect 7432 16396 7438 16448
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 8220 16445 8248 16544
rect 8389 16541 8401 16544
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8754 16572 8760 16584
rect 8619 16544 8760 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8404 16504 8432 16535
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16572 8999 16575
rect 9232 16572 9260 16680
rect 11241 16677 11253 16711
rect 11287 16708 11299 16711
rect 11514 16708 11520 16720
rect 11287 16680 11520 16708
rect 11287 16677 11299 16680
rect 11241 16671 11299 16677
rect 11514 16668 11520 16680
rect 11572 16708 11578 16720
rect 12406 16708 12434 16748
rect 12713 16745 12725 16779
rect 12759 16776 12771 16779
rect 12802 16776 12808 16788
rect 12759 16748 12808 16776
rect 12759 16745 12771 16748
rect 12713 16739 12771 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 13320 16748 13369 16776
rect 13320 16736 13326 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 11572 16680 12112 16708
rect 12406 16680 13124 16708
rect 11572 16668 11578 16680
rect 12084 16652 12112 16680
rect 12066 16640 12072 16652
rect 10888 16612 11928 16640
rect 12027 16612 12072 16640
rect 8987 16544 9260 16572
rect 9861 16575 9919 16581
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 9950 16572 9956 16584
rect 9907 16544 9956 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10888 16572 10916 16612
rect 10060 16544 10916 16572
rect 11900 16572 11928 16612
rect 12066 16600 12072 16612
rect 12124 16640 12130 16652
rect 12124 16612 12848 16640
rect 12124 16600 12130 16612
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11900 16544 12265 16572
rect 9030 16504 9036 16516
rect 8404 16476 9036 16504
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 10060 16504 10088 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 12820 16581 12848 16612
rect 13096 16581 13124 16680
rect 13464 16612 14412 16640
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 12400 16544 12541 16572
rect 12400 16532 12406 16544
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16572 13231 16575
rect 13464 16572 13492 16612
rect 13219 16544 13492 16572
rect 13219 16541 13231 16544
rect 13173 16535 13231 16541
rect 13538 16532 13544 16584
rect 13596 16532 13602 16584
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13679 16544 14105 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 10134 16513 10140 16516
rect 9508 16476 10088 16504
rect 7929 16439 7987 16445
rect 7929 16436 7941 16439
rect 7708 16408 7941 16436
rect 7708 16396 7714 16408
rect 7929 16405 7941 16408
rect 7975 16405 7987 16439
rect 7929 16399 7987 16405
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16405 8263 16439
rect 8205 16399 8263 16405
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 9508 16436 9536 16476
rect 10128 16467 10140 16513
rect 10134 16464 10140 16467
rect 10192 16464 10198 16516
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12897 16507 12955 16513
rect 12897 16504 12909 16507
rect 12216 16476 12909 16504
rect 12216 16464 12222 16476
rect 12897 16473 12909 16476
rect 12943 16473 12955 16507
rect 13446 16504 13452 16516
rect 12897 16467 12955 16473
rect 13280 16476 13452 16504
rect 13280 16448 13308 16476
rect 13446 16464 13452 16476
rect 13504 16504 13510 16516
rect 13648 16504 13676 16535
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 14384 16572 14412 16612
rect 15010 16572 15016 16584
rect 14384 16544 15016 16572
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 13504 16476 13676 16504
rect 13504 16464 13510 16476
rect 8720 16408 9536 16436
rect 8720 16396 8726 16408
rect 9582 16396 9588 16448
rect 9640 16396 9646 16448
rect 11517 16439 11575 16445
rect 11517 16405 11529 16439
rect 11563 16436 11575 16439
rect 11790 16436 11796 16448
rect 11563 16408 11796 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 12342 16396 12348 16448
rect 12400 16396 12406 16448
rect 13262 16396 13268 16448
rect 13320 16396 13326 16448
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 13906 16436 13912 16448
rect 13863 16408 13912 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 14292 16445 14320 16532
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16405 14335 16439
rect 14277 16399 14335 16405
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 1394 16192 1400 16244
rect 1452 16192 1458 16244
rect 2774 16232 2780 16244
rect 2746 16192 2780 16232
rect 2832 16192 2838 16244
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3878 16232 3884 16244
rect 3283 16204 3884 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 4706 16232 4712 16244
rect 4571 16204 4712 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 4706 16192 4712 16204
rect 4764 16232 4770 16244
rect 4764 16204 4936 16232
rect 4764 16192 4770 16204
rect 1412 16164 1440 16192
rect 2746 16164 2774 16192
rect 4338 16164 4344 16176
rect 1412 16136 3096 16164
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 2746 16105 2774 16136
rect 3068 16105 3096 16136
rect 3896 16136 4344 16164
rect 2746 16099 2827 16105
rect 2746 16068 2781 16099
rect 2769 16065 2781 16068
rect 2815 16065 2827 16099
rect 2769 16059 2827 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3329 16099 3387 16105
rect 3329 16096 3341 16099
rect 3099 16068 3341 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3329 16065 3341 16068
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3896 16105 3924 16136
rect 4338 16124 4344 16136
rect 4396 16124 4402 16176
rect 4798 16124 4804 16176
rect 4856 16124 4862 16176
rect 4908 16164 4936 16204
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5040 16204 5672 16232
rect 5040 16192 5046 16204
rect 5644 16173 5672 16204
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7193 16235 7251 16241
rect 7193 16232 7205 16235
rect 6788 16204 7205 16232
rect 6788 16192 6794 16204
rect 7193 16201 7205 16204
rect 7239 16201 7251 16235
rect 7193 16195 7251 16201
rect 7374 16192 7380 16244
rect 7432 16192 7438 16244
rect 8757 16235 8815 16241
rect 8757 16201 8769 16235
rect 8803 16232 8815 16235
rect 9306 16232 9312 16244
rect 8803 16204 9312 16232
rect 8803 16201 8815 16204
rect 8757 16195 8815 16201
rect 9306 16192 9312 16204
rect 9364 16232 9370 16244
rect 9582 16232 9588 16244
rect 9364 16204 9588 16232
rect 9364 16192 9370 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 11241 16235 11299 16241
rect 11241 16201 11253 16235
rect 11287 16232 11299 16235
rect 12526 16232 12532 16244
rect 11287 16204 12532 16232
rect 11287 16201 11299 16204
rect 11241 16195 11299 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13446 16232 13452 16244
rect 12768 16204 13452 16232
rect 12768 16192 12774 16204
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 13906 16192 13912 16244
rect 13964 16192 13970 16244
rect 5537 16167 5595 16173
rect 5537 16164 5549 16167
rect 4908 16136 5549 16164
rect 5537 16133 5549 16136
rect 5583 16133 5595 16167
rect 5537 16127 5595 16133
rect 5629 16167 5687 16173
rect 5629 16133 5641 16167
rect 5675 16133 5687 16167
rect 5629 16127 5687 16133
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 5776 16136 6500 16164
rect 5776 16124 5782 16136
rect 6472 16105 6500 16136
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 3476 16068 3617 16096
rect 3476 16056 3482 16068
rect 3605 16065 3617 16068
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 6457 16099 6515 16105
rect 6457 16065 6469 16099
rect 6503 16065 6515 16099
rect 7392 16096 7420 16192
rect 9950 16124 9956 16176
rect 10008 16164 10014 16176
rect 13814 16164 13820 16176
rect 10008 16136 13820 16164
rect 10008 16124 10014 16136
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7392 16068 7665 16096
rect 6457 16059 6515 16065
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16096 8171 16099
rect 8386 16096 8392 16108
rect 8159 16068 8392 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 10318 16056 10324 16108
rect 10376 16105 10382 16108
rect 10612 16105 10640 16136
rect 10376 16096 10388 16105
rect 10597 16099 10655 16105
rect 10376 16068 10421 16096
rect 10376 16059 10388 16068
rect 10597 16065 10609 16099
rect 10643 16096 10655 16099
rect 10643 16068 10677 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 10376 16056 10382 16059
rect 10870 16056 10876 16108
rect 10928 16056 10934 16108
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 11532 16105 11560 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 11790 16105 11796 16108
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16096 11575 16099
rect 11784 16096 11796 16105
rect 11563 16068 11597 16096
rect 11751 16068 11796 16096
rect 11563 16065 11575 16068
rect 11517 16059 11575 16065
rect 11784 16059 11796 16068
rect 11790 16056 11796 16059
rect 11848 16056 11854 16108
rect 13630 16096 13636 16108
rect 12636 16068 13636 16096
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 15997 2467 16031
rect 2409 15991 2467 15997
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 16028 2651 16031
rect 2958 16028 2964 16040
rect 2639 16000 2964 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 2424 15960 2452 15991
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3436 16000 4077 16028
rect 3142 15960 3148 15972
rect 2424 15932 3148 15960
rect 3142 15920 3148 15932
rect 3200 15920 3206 15972
rect 3436 15969 3464 16000
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 4065 15991 4123 15997
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 15997 4767 16031
rect 4709 15991 4767 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15929 3479 15963
rect 3421 15923 3479 15929
rect 3602 15920 3608 15972
rect 3660 15960 3666 15972
rect 4724 15960 4752 15991
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 7558 15988 7564 16040
rect 7616 16028 7622 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7616 16000 7849 16028
rect 7616 15988 7622 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8294 15988 8300 16040
rect 8352 15988 8358 16040
rect 10781 16031 10839 16037
rect 10781 15997 10793 16031
rect 10827 16028 10839 16031
rect 10962 16028 10968 16040
rect 10827 16000 10968 16028
rect 10827 15997 10839 16000
rect 10781 15991 10839 15997
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 3660 15932 4752 15960
rect 5261 15963 5319 15969
rect 3660 15920 3666 15932
rect 5261 15929 5273 15963
rect 5307 15960 5319 15963
rect 6089 15963 6147 15969
rect 6089 15960 6101 15963
rect 5307 15932 6101 15960
rect 5307 15929 5319 15932
rect 5261 15923 5319 15929
rect 6089 15929 6101 15932
rect 6135 15960 6147 15963
rect 6135 15932 9352 15960
rect 6135 15929 6147 15932
rect 6089 15923 6147 15929
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1489 15895 1547 15901
rect 1489 15892 1501 15895
rect 992 15864 1501 15892
rect 992 15852 998 15864
rect 1489 15861 1501 15864
rect 1535 15861 1547 15895
rect 1489 15855 1547 15861
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 2406 15892 2412 15904
rect 2271 15864 2412 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3050 15892 3056 15904
rect 2915 15864 3056 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 3694 15852 3700 15904
rect 3752 15852 3758 15904
rect 7006 15852 7012 15904
rect 7064 15852 7070 15904
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9214 15892 9220 15904
rect 8812 15864 9220 15892
rect 8812 15852 8818 15864
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9324 15892 9352 15932
rect 10612 15932 10916 15960
rect 10612 15892 10640 15932
rect 9324 15864 10640 15892
rect 10888 15892 10916 15932
rect 12636 15892 12664 16068
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 13924 16105 13952 16192
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13262 16028 13268 16040
rect 13127 16000 13268 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 12710 15920 12716 15972
rect 12768 15960 12774 15972
rect 13725 15963 13783 15969
rect 13725 15960 13737 15963
rect 12768 15932 13737 15960
rect 12768 15920 12774 15932
rect 13725 15929 13737 15932
rect 13771 15929 13783 15963
rect 13725 15923 13783 15929
rect 10888 15864 12664 15892
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13262 15892 13268 15904
rect 12943 15864 13268 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13630 15852 13636 15904
rect 13688 15852 13694 15904
rect 14366 15852 14372 15904
rect 14424 15852 14430 15904
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2593 15691 2651 15697
rect 2593 15688 2605 15691
rect 2556 15660 2605 15688
rect 2556 15648 2562 15660
rect 2593 15657 2605 15660
rect 2639 15657 2651 15691
rect 2593 15651 2651 15657
rect 3142 15648 3148 15700
rect 3200 15688 3206 15700
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 3200 15660 3525 15688
rect 3200 15648 3206 15660
rect 3513 15657 3525 15660
rect 3559 15657 3571 15691
rect 3513 15651 3571 15657
rect 3602 15648 3608 15700
rect 3660 15648 3666 15700
rect 3694 15648 3700 15700
rect 3752 15648 3758 15700
rect 3786 15648 3792 15700
rect 3844 15648 3850 15700
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4246 15688 4252 15700
rect 4111 15660 4252 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 5166 15648 5172 15700
rect 5224 15648 5230 15700
rect 5721 15691 5779 15697
rect 5721 15657 5733 15691
rect 5767 15688 5779 15691
rect 6638 15688 6644 15700
rect 5767 15660 6644 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 7006 15648 7012 15700
rect 7064 15648 7070 15700
rect 7650 15648 7656 15700
rect 7708 15648 7714 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8386 15688 8392 15700
rect 8067 15660 8392 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8570 15648 8576 15700
rect 8628 15648 8634 15700
rect 13354 15648 13360 15700
rect 13412 15648 13418 15700
rect 1857 15623 1915 15629
rect 1857 15589 1869 15623
rect 1903 15620 1915 15623
rect 3329 15623 3387 15629
rect 1903 15592 2774 15620
rect 1903 15589 1915 15592
rect 1857 15583 1915 15589
rect 2222 15552 2228 15564
rect 1688 15524 2228 15552
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 1688 15493 1716 15524
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 2746 15552 2774 15592
rect 3329 15589 3341 15623
rect 3375 15620 3387 15623
rect 3620 15620 3648 15648
rect 3375 15592 3648 15620
rect 3375 15589 3387 15592
rect 3329 15583 3387 15589
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2746 15524 2881 15552
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 3712 15552 3740 15648
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 3712 15524 4537 15552
rect 2869 15515 2927 15521
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 2056 15416 2084 15447
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 2685 15487 2743 15493
rect 2685 15484 2697 15487
rect 2556 15456 2697 15484
rect 2556 15444 2562 15456
rect 2685 15453 2697 15456
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 3651 15456 3685 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 2130 15416 2136 15428
rect 2056 15388 2136 15416
rect 2130 15376 2136 15388
rect 2188 15416 2194 15428
rect 3418 15416 3424 15428
rect 2188 15388 3424 15416
rect 2188 15376 2194 15388
rect 3418 15376 3424 15388
rect 3476 15416 3482 15428
rect 3620 15416 3648 15447
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5184 15484 5212 15648
rect 5994 15620 6000 15632
rect 5031 15456 5212 15484
rect 5460 15592 6000 15620
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 3786 15416 3792 15428
rect 3476 15388 3792 15416
rect 3476 15376 3482 15388
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 4724 15416 4752 15447
rect 5460 15416 5488 15592
rect 5994 15580 6000 15592
rect 6052 15620 6058 15632
rect 6052 15592 6664 15620
rect 6052 15580 6058 15592
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5951 15524 6561 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 6043 15456 6285 15484
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 6273 15453 6285 15456
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6365 15487 6423 15493
rect 6365 15453 6377 15487
rect 6411 15484 6423 15487
rect 6636 15484 6664 15592
rect 7024 15552 7052 15648
rect 7561 15555 7619 15561
rect 7024 15524 7512 15552
rect 6411 15456 6664 15484
rect 6411 15453 6423 15456
rect 6365 15447 6423 15453
rect 4724 15388 5488 15416
rect 5552 15416 5580 15447
rect 6288 15416 6316 15447
rect 7374 15444 7380 15496
rect 7432 15444 7438 15496
rect 7484 15484 7512 15524
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 7668 15552 7696 15648
rect 8588 15620 8616 15648
rect 10778 15620 10784 15632
rect 8588 15592 10784 15620
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 12342 15620 12348 15632
rect 11204 15592 12348 15620
rect 11204 15580 11210 15592
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 12802 15580 12808 15632
rect 12860 15580 12866 15632
rect 9953 15555 10011 15561
rect 7607 15524 7696 15552
rect 8220 15524 9168 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 8113 15487 8171 15493
rect 8113 15484 8125 15487
rect 7484 15456 8125 15484
rect 8113 15453 8125 15456
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 8220 15416 8248 15524
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 9030 15484 9036 15496
rect 8343 15456 9036 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9140 15493 9168 15524
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10226 15552 10232 15564
rect 9999 15524 10232 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9214 15484 9220 15496
rect 9171 15456 9220 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9214 15444 9220 15456
rect 9272 15484 9278 15496
rect 9968 15484 9996 15515
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 10468 15524 11192 15552
rect 10468 15512 10474 15524
rect 9272 15456 9996 15484
rect 9272 15444 9278 15456
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 11164 15493 11192 15524
rect 11606 15512 11612 15564
rect 11664 15552 11670 15564
rect 11882 15552 11888 15564
rect 11664 15524 11888 15552
rect 11664 15512 11670 15524
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12299 15524 12633 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 13372 15552 13400 15648
rect 13311 15524 13400 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 5552 15388 6132 15416
rect 6288 15388 8248 15416
rect 8757 15419 8815 15425
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 6104 15357 6132 15388
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 9674 15416 9680 15428
rect 8803 15388 9680 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 9674 15376 9680 15388
rect 9732 15416 9738 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 9732 15388 10241 15416
rect 9732 15376 9738 15388
rect 10229 15385 10241 15388
rect 10275 15385 10287 15419
rect 10229 15379 10287 15385
rect 10321 15419 10379 15425
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 10980 15416 11008 15444
rect 10367 15388 11008 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11256 15416 11284 15447
rect 11112 15388 11284 15416
rect 12360 15416 12388 15447
rect 12434 15444 12440 15496
rect 12492 15444 12498 15496
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 13262 15416 13268 15428
rect 12360 15388 13268 15416
rect 11112 15376 11118 15388
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 13357 15419 13415 15425
rect 13357 15385 13369 15419
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 6089 15351 6147 15357
rect 6089 15317 6101 15351
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 8938 15308 8944 15360
rect 8996 15308 9002 15360
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9180 15320 9321 15348
rect 9180 15308 9186 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 9309 15311 9367 15317
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 10100 15320 10977 15348
rect 10100 15308 10106 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 11425 15351 11483 15357
rect 11425 15317 11437 15351
rect 11471 15348 11483 15351
rect 11606 15348 11612 15360
rect 11471 15320 11612 15348
rect 11471 15317 11483 15320
rect 11425 15311 11483 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 13372 15348 13400 15379
rect 13906 15376 13912 15428
rect 13964 15376 13970 15428
rect 14185 15351 14243 15357
rect 14185 15348 14197 15351
rect 13372 15320 14197 15348
rect 14185 15317 14197 15320
rect 14231 15317 14243 15351
rect 14185 15311 14243 15317
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2038 15144 2044 15156
rect 1627 15116 2044 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3421 15147 3479 15153
rect 2148 15116 3372 15144
rect 2148 15076 2176 15116
rect 1688 15048 2176 15076
rect 1578 14968 1584 15020
rect 1636 14968 1642 15020
rect 1688 15017 1716 15048
rect 2222 15036 2228 15088
rect 2280 15076 2286 15088
rect 2406 15076 2412 15088
rect 2280 15048 2412 15076
rect 2280 15036 2286 15048
rect 2406 15036 2412 15048
rect 2464 15076 2470 15088
rect 3344 15076 3372 15116
rect 3421 15113 3433 15147
rect 3467 15144 3479 15147
rect 3602 15144 3608 15156
rect 3467 15116 3608 15144
rect 3467 15113 3479 15116
rect 3421 15107 3479 15113
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4890 15144 4896 15156
rect 3712 15116 4896 15144
rect 3712 15076 3740 15116
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8386 15144 8392 15156
rect 8343 15116 8392 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9732 15116 9965 15144
rect 9732 15104 9738 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 11698 15104 11704 15156
rect 11756 15104 11762 15156
rect 12161 15147 12219 15153
rect 12161 15113 12173 15147
rect 12207 15144 12219 15147
rect 12434 15144 12440 15156
rect 12207 15116 12440 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12434 15104 12440 15116
rect 12492 15104 12498 15156
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 13780 15116 14228 15144
rect 13780 15104 13786 15116
rect 5258 15076 5264 15088
rect 2464 15048 2820 15076
rect 3344 15048 3740 15076
rect 3804 15048 4108 15076
rect 2464 15036 2470 15048
rect 2792 15017 2820 15048
rect 3804 15020 3832 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 1811 14980 2513 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3050 15008 3056 15020
rect 3007 14980 3056 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3234 14968 3240 15020
rect 3292 15008 3298 15020
rect 3513 15011 3571 15017
rect 3513 15008 3525 15011
rect 3292 14980 3525 15008
rect 3292 14968 3298 14980
rect 3513 14977 3525 14980
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 3786 14968 3792 15020
rect 3844 14968 3850 15020
rect 4080 15017 4108 15048
rect 4448 15048 5264 15076
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 14977 4123 15011
rect 4065 14971 4123 14977
rect 1596 14940 1624 14968
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1596 14912 1961 14940
rect 1949 14909 1961 14912
rect 1995 14909 2007 14943
rect 3988 14940 4016 14971
rect 4448 14940 4476 15048
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 9217 15079 9275 15085
rect 9217 15045 9229 15079
rect 9263 15076 9275 15079
rect 10152 15076 10180 15104
rect 9263 15048 10180 15076
rect 10597 15079 10655 15085
rect 9263 15045 9275 15048
rect 9217 15039 9275 15045
rect 10597 15045 10609 15079
rect 10643 15076 10655 15079
rect 10778 15076 10784 15088
rect 10643 15048 10784 15076
rect 10643 15045 10655 15048
rect 10597 15039 10655 15045
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 11146 15036 11152 15088
rect 11204 15036 11210 15088
rect 4522 14968 4528 15020
rect 4580 14968 4586 15020
rect 7558 14968 7564 15020
rect 7616 15008 7622 15020
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7616 14980 7665 15008
rect 7616 14968 7622 14980
rect 7653 14977 7665 14980
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 11716 15008 11744 15104
rect 13630 15036 13636 15088
rect 13688 15085 13694 15088
rect 13688 15076 13700 15085
rect 13688 15048 13733 15076
rect 13688 15039 13700 15048
rect 13688 15036 13694 15039
rect 11563 14980 11744 15008
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12124 14980 12449 15008
rect 12124 14968 12130 14980
rect 12437 14977 12449 14980
rect 12483 15008 12495 15011
rect 12526 15008 12532 15020
rect 12483 14980 12532 15008
rect 12483 14977 12495 14980
rect 12437 14971 12495 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14200 15017 14228 15116
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13872 14980 13921 15008
rect 13872 14968 13878 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 1949 14903 2007 14909
rect 2056 14912 4016 14940
rect 4080 14912 4476 14940
rect 1118 14832 1124 14884
rect 1176 14872 1182 14884
rect 2056 14872 2084 14912
rect 1176 14844 2084 14872
rect 1176 14832 1182 14844
rect 3234 14832 3240 14884
rect 3292 14872 3298 14884
rect 3789 14875 3847 14881
rect 3789 14872 3801 14875
rect 3292 14844 3801 14872
rect 3292 14832 3298 14844
rect 3789 14841 3801 14844
rect 3835 14841 3847 14875
rect 3789 14835 3847 14841
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 2498 14804 2504 14816
rect 2455 14776 2504 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 4080 14804 4108 14912
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6972 14912 7205 14940
rect 6972 14900 6978 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9398 14940 9404 14952
rect 8628 14912 9404 14940
rect 8628 14900 8634 14912
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 9858 14940 9864 14952
rect 9539 14912 9864 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 11020 14912 11253 14940
rect 11020 14900 11026 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 11747 14912 12357 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 14274 14832 14280 14884
rect 14332 14832 14338 14884
rect 3743 14776 4108 14804
rect 4157 14807 4215 14813
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4246 14804 4252 14816
rect 4203 14776 4252 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4706 14764 4712 14816
rect 4764 14764 4770 14816
rect 6638 14764 6644 14816
rect 6696 14764 6702 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 12529 14807 12587 14813
rect 12529 14804 12541 14807
rect 11756 14776 12541 14804
rect 11756 14764 11762 14776
rect 12529 14773 12541 14776
rect 12575 14804 12587 14807
rect 14292 14804 14320 14832
rect 12575 14776 14320 14804
rect 12575 14773 12587 14776
rect 12529 14767 12587 14773
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 1544 14572 2697 14600
rect 1544 14560 1550 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 4246 14560 4252 14612
rect 4304 14560 4310 14612
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14600 4491 14603
rect 4890 14600 4896 14612
rect 4479 14572 4896 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 7466 14560 7472 14612
rect 7524 14560 7530 14612
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7892 14572 8033 14600
rect 7892 14560 7898 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 9030 14560 9036 14612
rect 9088 14560 9094 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9916 14572 10149 14600
rect 9916 14560 9922 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 11698 14560 11704 14612
rect 11756 14560 11762 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12434 14600 12440 14612
rect 12207 14572 12440 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12802 14560 12808 14612
rect 12860 14560 12866 14612
rect 3326 14464 3332 14476
rect 2884 14436 3332 14464
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 2406 14396 2412 14408
rect 2363 14368 2412 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2590 14356 2596 14408
rect 2648 14356 2654 14408
rect 2884 14405 2912 14436
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 4264 14473 4292 14560
rect 7484 14532 7512 14560
rect 7484 14504 8156 14532
rect 4249 14467 4307 14473
rect 3436 14436 4200 14464
rect 3436 14405 3464 14436
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14396 3203 14399
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 3191 14368 3433 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3786 14356 3792 14408
rect 3844 14356 3850 14408
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4172 14396 4200 14436
rect 4249 14433 4261 14467
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7616 14436 7665 14464
rect 7616 14424 7622 14436
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 7653 14427 7711 14433
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 4172 14368 5457 14396
rect 4065 14359 4123 14365
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 1765 14331 1823 14337
rect 1765 14297 1777 14331
rect 1811 14328 1823 14331
rect 2225 14331 2283 14337
rect 2225 14328 2237 14331
rect 1811 14300 2237 14328
rect 1811 14297 1823 14300
rect 1765 14291 1823 14297
rect 2225 14297 2237 14300
rect 2271 14297 2283 14331
rect 3804 14328 3832 14356
rect 2225 14291 2283 14297
rect 2884 14300 3832 14328
rect 4080 14328 4108 14359
rect 4246 14328 4252 14340
rect 4080 14300 4252 14328
rect 2884 14272 2912 14300
rect 4246 14288 4252 14300
rect 4304 14288 4310 14340
rect 4522 14288 4528 14340
rect 4580 14288 4586 14340
rect 5460 14328 5488 14359
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 5592 14368 6929 14396
rect 5592 14356 5598 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7466 14356 7472 14408
rect 7524 14356 7530 14408
rect 8128 14405 8156 14504
rect 10042 14492 10048 14544
rect 10100 14492 10106 14544
rect 11716 14532 11744 14560
rect 10980 14504 11744 14532
rect 10060 14464 10088 14492
rect 9232 14436 10088 14464
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8938 14396 8944 14408
rect 8619 14368 8944 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 9232 14405 9260 14436
rect 10410 14424 10416 14476
rect 10468 14424 10474 14476
rect 10870 14424 10876 14476
rect 10928 14424 10934 14476
rect 10980 14473 11008 14504
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 11664 14436 11713 14464
rect 11664 14424 11670 14436
rect 11701 14433 11713 14436
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 12710 14464 12716 14476
rect 12667 14436 12716 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12820 14464 12848 14560
rect 13817 14535 13875 14541
rect 13817 14501 13829 14535
rect 13863 14532 13875 14535
rect 13906 14532 13912 14544
rect 13863 14504 13912 14532
rect 13863 14501 13875 14504
rect 13817 14495 13875 14501
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 12820 14436 13277 14464
rect 13265 14433 13277 14436
rect 13311 14433 13323 14467
rect 13265 14427 13323 14433
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 10042 14396 10048 14408
rect 9999 14368 10048 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 10042 14356 10048 14368
rect 10100 14396 10106 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 10100 14368 10241 14396
rect 10100 14356 10106 14368
rect 10229 14365 10241 14368
rect 10275 14396 10287 14399
rect 10428 14396 10456 14424
rect 10275 14368 10456 14396
rect 10888 14396 10916 14424
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 10888 14368 11069 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 12158 14396 12164 14408
rect 11563 14368 12164 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12434 14356 12440 14408
rect 12492 14356 12498 14408
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 6672 14331 6730 14337
rect 5460 14300 5580 14328
rect 2406 14220 2412 14272
rect 2464 14220 2470 14272
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 3326 14220 3332 14272
rect 3384 14220 3390 14272
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 3602 14260 3608 14272
rect 3559 14232 3608 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14260 4031 14263
rect 4540 14260 4568 14288
rect 4019 14232 4568 14260
rect 4019 14229 4031 14232
rect 3973 14223 4031 14229
rect 4798 14220 4804 14272
rect 4856 14220 4862 14272
rect 5552 14269 5580 14300
rect 6672 14297 6684 14331
rect 6718 14328 6730 14331
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 6718 14300 10333 14328
rect 6718 14297 6730 14300
rect 6672 14291 6730 14297
rect 10321 14297 10333 14300
rect 10367 14297 10379 14331
rect 10321 14291 10379 14297
rect 13354 14288 13360 14340
rect 13412 14288 13418 14340
rect 5537 14263 5595 14269
rect 5537 14229 5549 14263
rect 5583 14260 5595 14263
rect 5718 14260 5724 14272
rect 5583 14232 5724 14260
rect 5583 14229 5595 14232
rect 5537 14223 5595 14229
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 7098 14260 7104 14272
rect 7055 14232 7104 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 9306 14220 9312 14272
rect 9364 14220 9370 14272
rect 11241 14263 11299 14269
rect 11241 14229 11253 14263
rect 11287 14260 11299 14263
rect 11606 14260 11612 14272
rect 11287 14232 11612 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 13722 14260 13728 14272
rect 12032 14232 13728 14260
rect 12032 14220 12038 14232
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 14090 14220 14096 14272
rect 14148 14220 14154 14272
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1452 14028 1593 14056
rect 1452 14016 1458 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 2498 14016 2504 14068
rect 2556 14016 2562 14068
rect 2866 14056 2872 14068
rect 2746 14028 2872 14056
rect 2746 13988 2774 14028
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 4798 14056 4804 14068
rect 4080 14028 4804 14056
rect 1780 13960 2774 13988
rect 3993 13991 4051 13997
rect 1780 13929 1808 13960
rect 3993 13957 4005 13991
rect 4039 13988 4051 13991
rect 4080 13988 4108 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5534 14056 5540 14068
rect 4908 14028 5540 14056
rect 4039 13960 4108 13988
rect 4039 13957 4051 13960
rect 3993 13951 4051 13957
rect 4154 13948 4160 14000
rect 4212 13988 4218 14000
rect 4908 13988 4936 14028
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 7285 14059 7343 14065
rect 7285 14025 7297 14059
rect 7331 14056 7343 14059
rect 7466 14056 7472 14068
rect 7331 14028 7472 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7558 14016 7564 14068
rect 7616 14016 7622 14068
rect 8754 14056 8760 14068
rect 7668 14028 8760 14056
rect 4212 13960 4936 13988
rect 5368 13960 5764 13988
rect 4212 13948 4218 13960
rect 4264 13929 4292 13960
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1596 13892 1777 13920
rect 1596 13864 1624 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 1578 13812 1584 13864
rect 1636 13812 1642 13864
rect 1854 13812 1860 13864
rect 1912 13812 1918 13864
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 4540 13784 4568 13883
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4764 13892 5273 13920
rect 4764 13880 4770 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5368 13852 5396 13960
rect 5736 13929 5764 13960
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 4663 13824 5396 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 4540 13756 4844 13784
rect 4816 13716 4844 13756
rect 4890 13744 4896 13796
rect 4948 13744 4954 13796
rect 5460 13784 5488 13883
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7668 13929 7696 14028
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 10042 14056 10048 14068
rect 9171 14028 10048 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10318 14016 10324 14068
rect 10376 14016 10382 14068
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 10870 14056 10876 14068
rect 10643 14028 10876 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 11020 14028 11345 14056
rect 11020 14016 11026 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 7760 13960 9996 13988
rect 7760 13932 7788 13960
rect 9232 13932 9260 13960
rect 9968 13932 9996 13960
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6512 13892 7113 13920
rect 6512 13880 6518 13892
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 7742 13880 7748 13932
rect 7800 13880 7806 13932
rect 8012 13923 8070 13929
rect 8012 13889 8024 13923
rect 8058 13920 8070 13923
rect 9122 13920 9128 13932
rect 8058 13892 9128 13920
rect 8058 13889 8070 13892
rect 8012 13883 8070 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 9214 13880 9220 13932
rect 9272 13880 9278 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9473 13923 9531 13929
rect 9473 13920 9485 13923
rect 9364 13892 9485 13920
rect 9364 13880 9370 13892
rect 9473 13889 9485 13892
rect 9519 13889 9531 13923
rect 9473 13883 9531 13889
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10336 13920 10364 14016
rect 10888 13988 10916 14016
rect 10888 13960 11100 13988
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10336 13892 10885 13920
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 11072 13920 11100 13960
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 11532 13988 11560 14019
rect 11606 14016 11612 14068
rect 11664 14016 11670 14068
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12492 14028 12633 14056
rect 12492 14016 12498 14028
rect 12621 14025 12633 14028
rect 12667 14056 12679 14059
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12667 14028 12725 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 13412 14028 13737 14056
rect 13412 14016 13418 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 11204 13960 11560 13988
rect 11204 13948 11210 13960
rect 11238 13920 11244 13932
rect 11072 13892 11244 13920
rect 10873 13883 10931 13889
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 11624 13920 11652 14016
rect 14108 13988 14136 14016
rect 13924 13960 14136 13988
rect 13924 13929 13952 13960
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11624 13892 11713 13920
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13889 13967 13923
rect 13909 13883 13967 13889
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 6730 13852 6736 13864
rect 5583 13824 6736 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 6822 13812 6828 13864
rect 6880 13812 6886 13864
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 7374 13852 7380 13864
rect 7248 13824 7380 13852
rect 7248 13812 7254 13824
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10778 13852 10784 13864
rect 10735 13824 10784 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11882 13852 11888 13864
rect 11204 13824 11888 13852
rect 11204 13812 11210 13824
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 11974 13812 11980 13864
rect 12032 13812 12038 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12618 13852 12624 13864
rect 12207 13824 12624 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13262 13852 13268 13864
rect 13219 13824 13268 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 5905 13787 5963 13793
rect 5905 13784 5917 13787
rect 5460 13756 5917 13784
rect 5905 13753 5917 13756
rect 5951 13784 5963 13787
rect 6365 13787 6423 13793
rect 6365 13784 6377 13787
rect 5951 13756 6377 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 6365 13753 6377 13756
rect 6411 13753 6423 13787
rect 6365 13747 6423 13753
rect 5718 13716 5724 13728
rect 4816 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 14369 13719 14427 13725
rect 14369 13685 14381 13719
rect 14415 13716 14427 13719
rect 14458 13716 14464 13728
rect 14415 13688 14464 13716
rect 14415 13685 14427 13688
rect 14369 13679 14427 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 2038 13512 2044 13524
rect 1719 13484 2044 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2280 13484 2421 13512
rect 2280 13472 2286 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 3568 13484 3617 13512
rect 3568 13472 3574 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 3605 13475 3663 13481
rect 4246 13472 4252 13524
rect 4304 13472 4310 13524
rect 6638 13512 6644 13524
rect 4356 13484 6644 13512
rect 1946 13404 1952 13456
rect 2004 13444 2010 13456
rect 2004 13416 3556 13444
rect 2004 13404 2010 13416
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 2406 13376 2412 13388
rect 2271 13348 2412 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 3528 13320 3556 13416
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 4356 13444 4384 13484
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 6788 13484 7205 13512
rect 6788 13472 6794 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7742 13512 7748 13524
rect 7193 13475 7251 13481
rect 7392 13484 7748 13512
rect 4120 13416 4384 13444
rect 4120 13404 4126 13416
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 6748 13444 6776 13472
rect 5040 13416 6776 13444
rect 5040 13404 5046 13416
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7064 13416 7328 13444
rect 7064 13404 7070 13416
rect 7300 13388 7328 13416
rect 4540 13348 7144 13376
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1596 13280 1777 13308
rect 1596 13252 1624 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 1946 13268 1952 13320
rect 2004 13308 2010 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 2004 13280 2053 13308
rect 2004 13268 2010 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3568 13280 3801 13308
rect 3568 13268 3574 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 4540 13317 4568 13348
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4856 13280 4997 13308
rect 4856 13268 4862 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 7006 13268 7012 13320
rect 7064 13268 7070 13320
rect 7116 13317 7144 13348
rect 7282 13336 7288 13388
rect 7340 13336 7346 13388
rect 7392 13385 7420 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8536 13484 9045 13512
rect 8536 13472 8542 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10134 13512 10140 13524
rect 9999 13484 10140 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10962 13472 10968 13524
rect 11020 13472 11026 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12676 13484 12909 13512
rect 12676 13472 12682 13484
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 13262 13472 13268 13524
rect 13320 13472 13326 13524
rect 10042 13404 10048 13456
rect 10100 13404 10106 13456
rect 10778 13404 10784 13456
rect 10836 13444 10842 13456
rect 12161 13447 12219 13453
rect 12161 13444 12173 13447
rect 10836 13416 12173 13444
rect 10836 13404 10842 13416
rect 12161 13413 12173 13416
rect 12207 13413 12219 13447
rect 12161 13407 12219 13413
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 9306 13376 9312 13388
rect 8812 13348 9312 13376
rect 8812 13336 8818 13348
rect 9306 13336 9312 13348
rect 9364 13376 9370 13388
rect 9364 13348 9444 13376
rect 9364 13336 9370 13348
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 8202 13308 8208 13320
rect 7147 13280 8208 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9416 13317 9444 13348
rect 10060 13317 10088 13404
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10183 13348 10517 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 11238 13336 11244 13388
rect 11296 13336 11302 13388
rect 13354 13336 13360 13388
rect 13412 13336 13418 13388
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9815 13280 10057 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 1578 13200 1584 13252
rect 1636 13200 1642 13252
rect 1670 13200 1676 13252
rect 1728 13240 1734 13252
rect 7466 13240 7472 13252
rect 1728 13212 6960 13240
rect 1728 13200 1734 13212
rect 4706 13132 4712 13184
rect 4764 13132 4770 13184
rect 5077 13175 5135 13181
rect 5077 13141 5089 13175
rect 5123 13172 5135 13175
rect 5258 13172 5264 13184
rect 5123 13144 5264 13172
rect 5123 13141 5135 13144
rect 5077 13135 5135 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5534 13132 5540 13184
rect 5592 13132 5598 13184
rect 6932 13172 6960 13212
rect 7116 13212 7472 13240
rect 7116 13172 7144 13212
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 7650 13249 7656 13252
rect 7644 13203 7656 13249
rect 7650 13200 7656 13203
rect 7708 13200 7714 13252
rect 8956 13184 8984 13271
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13308 11207 13311
rect 11256 13308 11284 13336
rect 11195 13280 11284 13308
rect 11793 13311 11851 13317
rect 11195 13277 11207 13280
rect 11149 13271 11207 13277
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11808 13240 11836 13271
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12526 13308 12532 13320
rect 12124 13280 12532 13308
rect 12124 13268 12130 13280
rect 12526 13268 12532 13280
rect 12584 13308 12590 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12584 13280 12817 13308
rect 12584 13268 12590 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13096 13240 13124 13271
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13320 13280 14289 13308
rect 13320 13268 13326 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 11808 13212 12020 13240
rect 11992 13184 12020 13212
rect 12728 13212 13124 13240
rect 6932 13144 7144 13172
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8628 13144 8769 13172
rect 8628 13132 8634 13144
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 9180 13144 9229 13172
rect 9180 13132 9186 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9217 13135 9275 13141
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 11698 13132 11704 13184
rect 11756 13132 11762 13184
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 12728 13181 12756 13212
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 13998 13240 14004 13252
rect 13596 13212 14004 13240
rect 13596 13200 13602 13212
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 12713 13175 12771 13181
rect 12713 13141 12725 13175
rect 12759 13141 12771 13175
rect 12713 13135 12771 13141
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 13872 13144 14105 13172
rect 13872 13132 13878 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 1949 12971 2007 12977
rect 1949 12968 1961 12971
rect 1912 12940 1961 12968
rect 1912 12928 1918 12940
rect 1949 12937 1961 12940
rect 1995 12937 2007 12971
rect 1949 12931 2007 12937
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2314 12968 2320 12980
rect 2271 12940 2320 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 3234 12928 3240 12980
rect 3292 12928 3298 12980
rect 3326 12928 3332 12980
rect 3384 12928 3390 12980
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 3970 12968 3976 12980
rect 3467 12940 3976 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4246 12968 4252 12980
rect 4203 12940 4252 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12937 5687 12971
rect 5629 12931 5687 12937
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6181 12971 6239 12977
rect 5951 12940 6040 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 2406 12900 2412 12912
rect 1872 12872 2412 12900
rect 1578 12792 1584 12844
rect 1636 12792 1642 12844
rect 1872 12841 1900 12872
rect 2406 12860 2412 12872
rect 2464 12900 2470 12912
rect 3252 12900 3280 12928
rect 2464 12872 2636 12900
rect 2464 12860 2470 12872
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2130 12792 2136 12844
rect 2188 12792 2194 12844
rect 2498 12724 2504 12776
rect 2556 12724 2562 12776
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 2516 12696 2544 12724
rect 1811 12668 2544 12696
rect 2608 12696 2636 12872
rect 3160 12872 3280 12900
rect 3160 12841 3188 12872
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2731 12804 3157 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3344 12832 3372 12928
rect 5644 12900 5672 12931
rect 5644 12872 5948 12900
rect 3283 12804 3372 12832
rect 3513 12835 3571 12841
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 4249 12835 4307 12841
rect 4249 12832 4261 12835
rect 3559 12804 4261 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 4249 12801 4261 12804
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3528 12764 3556 12795
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 4580 12804 5365 12832
rect 4580 12792 4586 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5626 12832 5632 12844
rect 5491 12804 5632 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 3108 12736 3556 12764
rect 3108 12724 3114 12736
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3660 12736 3709 12764
rect 3660 12724 3666 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 4430 12724 4436 12776
rect 4488 12724 4494 12776
rect 5920 12764 5948 12872
rect 6012 12841 6040 12940
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6822 12968 6828 12980
rect 6227 12940 6828 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7098 12968 7104 12980
rect 7024 12940 7104 12968
rect 7024 12909 7052 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7282 12928 7288 12980
rect 7340 12928 7346 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 7524 12940 7573 12968
rect 7524 12928 7530 12940
rect 7561 12937 7573 12940
rect 7607 12937 7619 12971
rect 7561 12931 7619 12937
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9272 12940 9321 12968
rect 9272 12928 9278 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9674 12928 9680 12980
rect 9732 12928 9738 12980
rect 10778 12928 10784 12980
rect 10836 12928 10842 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11112 12940 11529 12968
rect 11112 12928 11118 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11882 12968 11888 12980
rect 11517 12931 11575 12937
rect 11624 12940 11888 12968
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 6288 12872 6929 12900
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6288 12764 6316 12872
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 6917 12863 6975 12869
rect 7009 12903 7067 12909
rect 7009 12869 7021 12903
rect 7055 12869 7067 12903
rect 7300 12900 7328 12928
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 7300 12872 7849 12900
rect 7009 12863 7067 12869
rect 7837 12869 7849 12872
rect 7883 12900 7895 12903
rect 8294 12900 8300 12912
rect 7883 12872 8300 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 9692 12900 9720 12928
rect 10965 12903 11023 12909
rect 9692 12872 10180 12900
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 8938 12832 8944 12844
rect 7791 12804 8944 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 10152 12841 10180 12872
rect 10965 12869 10977 12903
rect 11011 12900 11023 12903
rect 11624 12900 11652 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13817 12971 13875 12977
rect 12406 12940 13768 12968
rect 12066 12900 12072 12912
rect 11011 12872 11652 12900
rect 11716 12872 12072 12900
rect 11011 12869 11023 12872
rect 10965 12863 11023 12869
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 5920 12736 6316 12764
rect 6730 12724 6736 12776
rect 6788 12724 6794 12776
rect 9692 12764 9720 12795
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 11716 12841 11744 12872
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 10284 12804 10885 12832
rect 10284 12792 10290 12804
rect 10873 12801 10885 12804
rect 10919 12832 10931 12835
rect 11701 12835 11759 12841
rect 10919 12804 11008 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 10244 12764 10272 12792
rect 10980 12776 11008 12804
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12832 11851 12835
rect 12406 12832 12434 12940
rect 11839 12804 12434 12832
rect 11839 12801 11851 12804
rect 11793 12795 11851 12801
rect 9692 12736 10272 12764
rect 10318 12724 10324 12776
rect 10376 12724 10382 12776
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 11808 12764 11836 12795
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13740 12832 13768 12940
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 13863 12940 14136 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 14108 12909 14136 12940
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 15194 12832 15200 12844
rect 13740 12804 15200 12832
rect 13633 12795 13691 12801
rect 11882 12764 11888 12776
rect 11808 12736 11888 12764
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 13648 12764 13676 12795
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 12492 12736 13676 12764
rect 12492 12724 12498 12736
rect 15286 12696 15292 12708
rect 2608 12668 15292 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 2869 12631 2927 12637
rect 2869 12597 2881 12631
rect 2915 12628 2927 12631
rect 4062 12628 4068 12640
rect 2915 12600 4068 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4614 12588 4620 12640
rect 4672 12588 4678 12640
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 9858 12588 9864 12640
rect 9916 12588 9922 12640
rect 11885 12631 11943 12637
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 11974 12628 11980 12640
rect 11931 12600 11980 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12710 12588 12716 12640
rect 12768 12588 12774 12640
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12860 12600 13461 12628
rect 12860 12588 12866 12600
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 14369 12631 14427 12637
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 14918 12628 14924 12640
rect 14415 12600 14924 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2130 12424 2136 12436
rect 1627 12396 2136 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 12434 12424 12440 12436
rect 2746 12396 12440 12424
rect 2746 12356 2774 12396
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 14090 12384 14096 12436
rect 14148 12384 14154 12436
rect 1780 12328 2774 12356
rect 4157 12359 4215 12365
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1780 12229 1808 12328
rect 4157 12325 4169 12359
rect 4203 12356 4215 12359
rect 4430 12356 4436 12368
rect 4203 12328 4436 12356
rect 4203 12325 4215 12328
rect 4157 12319 4215 12325
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 5350 12356 5356 12368
rect 4672 12328 5356 12356
rect 4672 12316 4678 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5626 12316 5632 12368
rect 5684 12356 5690 12368
rect 5997 12359 6055 12365
rect 5997 12356 6009 12359
rect 5684 12328 6009 12356
rect 5684 12316 5690 12328
rect 5997 12325 6009 12328
rect 6043 12325 6055 12359
rect 5997 12319 6055 12325
rect 7834 12316 7840 12368
rect 7892 12316 7898 12368
rect 10045 12359 10103 12365
rect 10045 12325 10057 12359
rect 10091 12356 10103 12359
rect 10318 12356 10324 12368
rect 10091 12328 10324 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 10318 12316 10324 12328
rect 10376 12316 10382 12368
rect 10410 12316 10416 12368
rect 10468 12316 10474 12368
rect 12342 12316 12348 12368
rect 12400 12316 12406 12368
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 1912 12260 2053 12288
rect 1912 12248 1918 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2958 12248 2964 12300
rect 3016 12248 3022 12300
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5166 12288 5172 12300
rect 4847 12260 5172 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6086 12288 6092 12300
rect 5592 12260 6092 12288
rect 5592 12248 5598 12260
rect 6086 12248 6092 12260
rect 6144 12288 6150 12300
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6144 12260 6377 12288
rect 6144 12248 6150 12260
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7432 12260 8309 12288
rect 7432 12248 7438 12260
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8628 12260 9045 12288
rect 8628 12248 8634 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 9272 12260 10977 12288
rect 9272 12248 9278 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 992 12192 1409 12220
rect 992 12180 998 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1765 12223 1823 12229
rect 1765 12220 1777 12223
rect 1397 12183 1455 12189
rect 1504 12192 1777 12220
rect 1504 12096 1532 12192
rect 1765 12189 1777 12192
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 1946 12180 1952 12232
rect 2004 12180 2010 12232
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 1857 12155 1915 12161
rect 1857 12121 1869 12155
rect 1903 12152 1915 12155
rect 1964 12152 1992 12180
rect 1903 12124 1992 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 2240 12152 2268 12183
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3835 12192 4077 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 4065 12189 4077 12192
rect 4111 12220 4123 12223
rect 4111 12192 4660 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4522 12152 4528 12164
rect 2096 12124 2268 12152
rect 3988 12124 4528 12152
rect 2096 12112 2102 12124
rect 1486 12044 1492 12096
rect 1544 12044 1550 12096
rect 2498 12044 2504 12096
rect 2556 12084 2562 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2556 12056 2697 12084
rect 2556 12044 2562 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2685 12047 2743 12053
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 3694 12084 3700 12096
rect 3651 12056 3700 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3988 12093 4016 12124
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12053 4031 12087
rect 4632 12084 4660 12192
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5960 12192 6193 12220
rect 5960 12180 5966 12192
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6621 12223 6679 12229
rect 6621 12220 6633 12223
rect 6512 12192 6633 12220
rect 6512 12180 6518 12192
rect 6621 12189 6633 12192
rect 6667 12189 6679 12223
rect 6621 12183 6679 12189
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12220 8815 12223
rect 8803 12192 8892 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 5169 12155 5227 12161
rect 5169 12121 5181 12155
rect 5215 12121 5227 12155
rect 5169 12115 5227 12121
rect 5074 12084 5080 12096
rect 4632 12056 5080 12084
rect 3973 12047 4031 12053
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 5184 12084 5212 12115
rect 5258 12112 5264 12164
rect 5316 12112 5322 12164
rect 5350 12112 5356 12164
rect 5408 12112 5414 12164
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12152 5871 12155
rect 5994 12152 6000 12164
rect 5859 12124 6000 12152
rect 5859 12121 5871 12124
rect 5813 12115 5871 12121
rect 5994 12112 6000 12124
rect 6052 12152 6058 12164
rect 6730 12152 6736 12164
rect 6052 12124 6736 12152
rect 6052 12112 6058 12124
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 8864 12152 8892 12192
rect 9858 12180 9864 12232
rect 9916 12180 9922 12232
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11054 12220 11060 12232
rect 10919 12192 11060 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 8496 12124 8892 12152
rect 5368 12084 5396 12112
rect 5184 12056 5396 12084
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 8496 12084 8524 12124
rect 8864 12096 8892 12124
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12152 9183 12155
rect 9214 12152 9220 12164
rect 9171 12124 9220 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 9677 12155 9735 12161
rect 9677 12121 9689 12155
rect 9723 12121 9735 12155
rect 10704 12152 10732 12183
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11232 12223 11290 12229
rect 11232 12189 11244 12223
rect 11278 12220 11290 12223
rect 11698 12220 11704 12232
rect 11278 12192 11704 12220
rect 11278 12189 11290 12192
rect 11232 12183 11290 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12360 12220 12388 12316
rect 12526 12288 12532 12300
rect 12452 12260 12532 12288
rect 12452 12229 12480 12260
rect 12526 12248 12532 12260
rect 12584 12288 12590 12300
rect 13446 12288 13452 12300
rect 12584 12260 13452 12288
rect 12584 12248 12590 12260
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 11992 12192 12388 12220
rect 12437 12223 12495 12229
rect 11882 12152 11888 12164
rect 10704 12124 11888 12152
rect 9677 12115 9735 12121
rect 7791 12056 8524 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 8846 12044 8852 12096
rect 8904 12044 8910 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9692 12084 9720 12115
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 11992 12084 12020 12192
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 15010 12220 15016 12232
rect 14323 12192 15016 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 12636 12152 12664 12180
rect 13354 12152 13360 12164
rect 12636 12124 13360 12152
rect 13354 12112 13360 12124
rect 13412 12152 13418 12164
rect 13449 12155 13507 12161
rect 13449 12152 13461 12155
rect 13412 12124 13461 12152
rect 13412 12112 13418 12124
rect 13449 12121 13461 12124
rect 13495 12121 13507 12155
rect 13449 12115 13507 12121
rect 9456 12056 12020 12084
rect 12345 12087 12403 12093
rect 9456 12044 9462 12056
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12434 12084 12440 12096
rect 12391 12056 12440 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12434 12044 12440 12056
rect 12492 12084 12498 12096
rect 13556 12084 13584 12183
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 12492 12056 13584 12084
rect 12492 12044 12498 12056
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 2958 11840 2964 11892
rect 3016 11840 3022 11892
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 4157 11883 4215 11889
rect 4157 11880 4169 11883
rect 3200 11852 4169 11880
rect 3200 11840 3206 11852
rect 4157 11849 4169 11852
rect 4203 11849 4215 11883
rect 4157 11843 4215 11849
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 7282 11880 7288 11892
rect 5132 11852 7288 11880
rect 5132 11840 5138 11852
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1535 11716 1777 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1765 11713 1777 11716
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 1780 11608 1808 11707
rect 1854 11704 1860 11756
rect 1912 11744 1918 11756
rect 2041 11747 2099 11753
rect 2041 11744 2053 11747
rect 1912 11716 2053 11744
rect 1912 11704 1918 11716
rect 2041 11713 2053 11716
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2222 11636 2228 11688
rect 2280 11636 2286 11688
rect 2792 11676 2820 11707
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 3016 11716 3065 11744
rect 3016 11704 3022 11716
rect 3053 11713 3065 11716
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3326 11704 3332 11756
rect 3384 11704 3390 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3436 11716 4261 11744
rect 3436 11676 3464 11716
rect 4249 11713 4261 11716
rect 4295 11744 4307 11747
rect 5833 11747 5891 11753
rect 4295 11716 5120 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 2792 11648 3464 11676
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3237 11611 3295 11617
rect 1780 11580 2535 11608
rect 1670 11500 1676 11552
rect 1728 11500 1734 11552
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 2406 11500 2412 11552
rect 2464 11500 2470 11552
rect 2507 11540 2535 11580
rect 3237 11577 3249 11611
rect 3283 11608 3295 11611
rect 3528 11608 3556 11639
rect 5092 11620 5120 11716
rect 5833 11713 5845 11747
rect 5879 11744 5891 11747
rect 5879 11716 6040 11744
rect 5879 11713 5891 11716
rect 5833 11707 5891 11713
rect 6012 11676 6040 11716
rect 6086 11704 6092 11756
rect 6144 11704 6150 11756
rect 6270 11704 6276 11756
rect 6328 11704 6334 11756
rect 6380 11753 6408 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7650 11840 7656 11892
rect 7708 11840 7714 11892
rect 10962 11840 10968 11892
rect 11020 11840 11026 11892
rect 11241 11883 11299 11889
rect 11241 11849 11253 11883
rect 11287 11849 11299 11883
rect 11241 11843 11299 11849
rect 6638 11772 6644 11824
rect 6696 11812 6702 11824
rect 7745 11815 7803 11821
rect 7745 11812 7757 11815
rect 6696 11784 7757 11812
rect 6696 11772 6702 11784
rect 7745 11781 7757 11784
rect 7791 11781 7803 11815
rect 7745 11775 7803 11781
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 8754 11744 8760 11756
rect 6963 11716 8760 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 8754 11704 8760 11716
rect 8812 11744 8818 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 8812 11716 9597 11744
rect 8812 11704 8818 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 10980 11744 11008 11840
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10980 11716 11069 11744
rect 9585 11707 9643 11713
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11256 11744 11284 11843
rect 11882 11840 11888 11892
rect 11940 11840 11946 11892
rect 12526 11840 12532 11892
rect 12584 11840 12590 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12986 11880 12992 11892
rect 12667 11852 12992 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13412 11852 13553 11880
rect 13412 11840 13418 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 13630 11840 13636 11892
rect 13688 11840 13694 11892
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11256 11716 11713 11744
rect 11057 11707 11115 11713
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12434 11744 12440 11756
rect 12299 11716 12440 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 6012 11648 6224 11676
rect 3283 11580 3556 11608
rect 3620 11580 4752 11608
rect 3283 11577 3295 11580
rect 3237 11571 3295 11577
rect 3620 11540 3648 11580
rect 4724 11552 4752 11580
rect 5074 11568 5080 11620
rect 5132 11568 5138 11620
rect 2507 11512 3648 11540
rect 3694 11500 3700 11552
rect 3752 11500 3758 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 5902 11540 5908 11552
rect 4764 11512 5908 11540
rect 4764 11500 4770 11512
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6196 11540 6224 11648
rect 6288 11608 6316 11704
rect 7006 11636 7012 11688
rect 7064 11636 7070 11688
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 8904 11648 10885 11676
rect 8904 11636 8910 11648
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 11072 11676 11100 11707
rect 11808 11676 11836 11707
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 12544 11753 12572 11840
rect 13648 11812 13676 11840
rect 13648 11784 13952 11812
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12768 11716 13093 11744
rect 12768 11704 12774 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13722 11704 13728 11756
rect 13780 11704 13786 11756
rect 13924 11753 13952 11784
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 11072 11648 11836 11676
rect 10873 11639 10931 11645
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12676 11648 12909 11676
rect 12676 11636 12682 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13262 11636 13268 11688
rect 13320 11636 13326 11688
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 6288 11580 6561 11608
rect 6549 11577 6561 11580
rect 6595 11577 6607 11611
rect 7190 11608 7196 11620
rect 6549 11571 6607 11577
rect 6748 11580 7196 11608
rect 6748 11540 6776 11580
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 9033 11611 9091 11617
rect 9033 11608 9045 11611
rect 8352 11580 9045 11608
rect 8352 11568 8358 11580
rect 9033 11577 9045 11580
rect 9079 11577 9091 11611
rect 9033 11571 9091 11577
rect 9214 11568 9220 11620
rect 9272 11568 9278 11620
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 12176 11608 12204 11636
rect 11112 11580 12204 11608
rect 12437 11611 12495 11617
rect 11112 11568 11118 11580
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 13280 11608 13308 11636
rect 12483 11580 13308 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 6196 11512 6776 11540
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 9232 11540 9260 11568
rect 6871 11512 9260 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 10226 11500 10232 11552
rect 10284 11500 10290 11552
rect 10318 11500 10324 11552
rect 10376 11500 10382 11552
rect 11514 11500 11520 11552
rect 11572 11500 11578 11552
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 14056 11512 14105 11540
rect 14056 11500 14062 11512
rect 14093 11509 14105 11512
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 1854 11296 1860 11348
rect 1912 11296 1918 11348
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2222 11336 2228 11348
rect 1995 11308 2228 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 8754 11296 8760 11348
rect 8812 11296 8818 11348
rect 10318 11336 10324 11348
rect 8956 11308 10324 11336
rect 1688 11200 1716 11296
rect 1872 11200 1900 11296
rect 4617 11271 4675 11277
rect 4617 11237 4629 11271
rect 4663 11268 4675 11271
rect 4798 11268 4804 11280
rect 4663 11240 4804 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 6825 11271 6883 11277
rect 6825 11237 6837 11271
rect 6871 11268 6883 11271
rect 7006 11268 7012 11280
rect 6871 11240 7012 11268
rect 6871 11237 6883 11240
rect 6825 11231 6883 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 1688 11172 1808 11200
rect 1872 11172 2329 11200
rect 1780 11141 1808 11172
rect 2317 11169 2329 11172
rect 2363 11169 2375 11203
rect 2317 11163 2375 11169
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2556 11172 2973 11200
rect 2556 11160 2562 11172
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 4982 11160 4988 11212
rect 5040 11160 5046 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 6472 11172 7389 11200
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 1688 11064 1716 11095
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 2004 11104 2145 11132
rect 2004 11092 2010 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 4847 11104 5181 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5169 11101 5181 11104
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5534 11132 5540 11144
rect 5491 11104 5540 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 1854 11064 1860 11076
rect 1688 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2222 11024 2228 11076
rect 2280 11064 2286 11076
rect 2406 11064 2412 11076
rect 2280 11036 2412 11064
rect 2280 11024 2286 11036
rect 2406 11024 2412 11036
rect 2464 11064 2470 11076
rect 2777 11067 2835 11073
rect 2777 11064 2789 11067
rect 2464 11036 2789 11064
rect 2464 11024 2470 11036
rect 2777 11033 2789 11036
rect 2823 11033 2835 11067
rect 2777 11027 2835 11033
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5276 11064 5304 11095
rect 5534 11092 5540 11104
rect 5592 11132 5598 11144
rect 6472 11132 6500 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 7377 11163 7435 11169
rect 5592 11104 6500 11132
rect 5592 11092 5598 11104
rect 7006 11092 7012 11144
rect 7064 11132 7070 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 7064 11104 7113 11132
rect 7064 11092 7070 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7644 11135 7702 11141
rect 7644 11101 7656 11135
rect 7690 11132 7702 11135
rect 8956 11132 8984 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 11514 11296 11520 11348
rect 11572 11296 11578 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11940 11308 11989 11336
rect 11940 11296 11946 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 11532 11268 11560 11296
rect 10888 11240 11560 11268
rect 11793 11271 11851 11277
rect 10888 11209 10916 11240
rect 11793 11237 11805 11271
rect 11839 11268 11851 11271
rect 11839 11240 14320 11268
rect 11839 11237 11851 11240
rect 11793 11231 11851 11237
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11169 10931 11203
rect 10873 11163 10931 11169
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11379 11172 12265 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12492 11172 12572 11200
rect 12492 11160 12498 11172
rect 7690 11104 8984 11132
rect 10065 11135 10123 11141
rect 7690 11101 7702 11104
rect 7644 11095 7702 11101
rect 10065 11101 10077 11135
rect 10111 11132 10123 11135
rect 10226 11132 10232 11144
rect 10111 11104 10232 11132
rect 10111 11101 10123 11104
rect 10065 11095 10123 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 11057 11135 11115 11141
rect 10367 11104 11008 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 5718 11073 5724 11076
rect 5132 11036 5304 11064
rect 5132 11024 5138 11036
rect 5712 11027 5724 11073
rect 5718 11024 5724 11027
rect 5776 11024 5782 11076
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10996 1639 10999
rect 2130 10996 2136 11008
rect 1627 10968 2136 10996
rect 1627 10965 1639 10968
rect 1581 10959 1639 10965
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 3970 10996 3976 11008
rect 3651 10968 3976 10996
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 6914 10956 6920 11008
rect 6972 10956 6978 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 8202 10996 8208 11008
rect 7340 10968 8208 10996
rect 7340 10956 7346 10968
rect 8202 10956 8208 10968
rect 8260 10996 8266 11008
rect 8941 10999 8999 11005
rect 8941 10996 8953 10999
rect 8260 10968 8953 10996
rect 8260 10956 8266 10968
rect 8941 10965 8953 10968
rect 8987 10965 8999 10999
rect 10980 10996 11008 11104
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11072 11064 11100 11095
rect 11422 11092 11428 11144
rect 11480 11132 11486 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11480 11104 11897 11132
rect 11480 11092 11486 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12544 11141 12572 11172
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 13262 11200 13268 11212
rect 12860 11172 13268 11200
rect 12860 11160 12866 11172
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11132 12403 11135
rect 12529 11135 12587 11141
rect 12391 11104 12480 11132
rect 12391 11101 12403 11104
rect 12345 11095 12403 11101
rect 12084 11064 12112 11092
rect 11072 11036 12112 11064
rect 12452 11064 12480 11104
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 13449 11135 13507 11141
rect 12575 11104 12940 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11064 12624 11076
rect 12452 11036 12624 11064
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 12912 11064 12940 11104
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 14090 11132 14096 11144
rect 13495 11104 14096 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14182 11092 14188 11144
rect 14240 11092 14246 11144
rect 13722 11064 13728 11076
rect 12912 11036 13728 11064
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 13909 11067 13967 11073
rect 13909 11033 13921 11067
rect 13955 11064 13967 11067
rect 14292 11064 14320 11240
rect 14384 11212 14412 11299
rect 14366 11160 14372 11212
rect 14424 11160 14430 11212
rect 14458 11064 14464 11076
rect 13955 11036 14464 11064
rect 13955 11033 13967 11036
rect 13909 11027 13967 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 11606 10996 11612 11008
rect 10980 10968 11612 10996
rect 8941 10959 8999 10965
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 13173 10999 13231 11005
rect 13173 10965 13185 10999
rect 13219 10996 13231 10999
rect 13354 10996 13360 11008
rect 13219 10968 13360 10996
rect 13219 10965 13231 10968
rect 13173 10959 13231 10965
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2038 10792 2044 10804
rect 1811 10764 2044 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2498 10752 2504 10804
rect 2556 10792 2562 10804
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2556 10764 2697 10792
rect 2556 10752 2562 10764
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3200 10764 3525 10792
rect 3200 10752 3206 10764
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 5718 10792 5724 10804
rect 5399 10764 5724 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10761 6699 10795
rect 6641 10755 6699 10761
rect 6656 10724 6684 10755
rect 8754 10752 8760 10804
rect 8812 10752 8818 10804
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 6917 10727 6975 10733
rect 6917 10724 6929 10727
rect 3620 10696 4844 10724
rect 3620 10668 3648 10696
rect 1578 10616 1584 10668
rect 1636 10616 1642 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 1688 10628 3249 10656
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1688 10588 1716 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3602 10616 3608 10668
rect 3660 10616 3666 10668
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4338 10656 4344 10668
rect 4203 10628 4344 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 1360 10560 1716 10588
rect 1360 10548 1366 10560
rect 1946 10548 1952 10600
rect 2004 10588 2010 10600
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 2004 10560 2053 10588
rect 2004 10548 2010 10560
rect 2041 10557 2053 10560
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2188 10560 2237 10588
rect 2188 10548 2194 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 3050 10588 3056 10600
rect 2823 10560 3056 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3896 10520 3924 10619
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4522 10656 4528 10668
rect 4479 10628 4528 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 4816 10665 4844 10696
rect 6012 10696 6592 10724
rect 6656 10696 6929 10724
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 4847 10628 5641 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 5629 10625 5641 10628
rect 5675 10656 5687 10659
rect 5902 10656 5908 10668
rect 5675 10628 5908 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 6012 10588 6040 10696
rect 6457 10659 6515 10665
rect 6457 10625 6469 10659
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 4028 10560 6040 10588
rect 4028 10548 4034 10560
rect 5350 10520 5356 10532
rect 3896 10492 5356 10520
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 6472 10520 6500 10619
rect 6564 10588 6592 10696
rect 6917 10693 6929 10696
rect 6963 10693 6975 10727
rect 6917 10687 6975 10693
rect 7466 10684 7472 10736
rect 7524 10724 7530 10736
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 7524 10696 7757 10724
rect 7524 10684 7530 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 7745 10687 7803 10693
rect 8570 10616 8576 10668
rect 8628 10616 8634 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8772 10656 8800 10752
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 10428 10724 10456 10755
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 14056 10764 14105 10792
rect 14056 10752 14062 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 14550 10724 14556 10736
rect 9171 10696 10456 10724
rect 10704 10696 14556 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 8711 10628 8800 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 9950 10616 9956 10668
rect 10008 10616 10014 10668
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6564 10560 6837 10588
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7650 10548 7656 10600
rect 7708 10548 7714 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8812 10560 9045 10588
rect 8812 10548 8818 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 10612 10588 10640 10619
rect 9508 10560 10640 10588
rect 6932 10520 6960 10548
rect 6472 10492 6960 10520
rect 7377 10523 7435 10529
rect 7377 10489 7389 10523
rect 7423 10520 7435 10523
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 7423 10492 8217 10520
rect 7423 10489 7435 10492
rect 7377 10483 7435 10489
rect 8205 10489 8217 10492
rect 8251 10520 8263 10523
rect 8849 10523 8907 10529
rect 8251 10492 8800 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 1820 10424 3065 10452
rect 1820 10412 1826 10424
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3568 10424 3801 10452
rect 3568 10412 3574 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 4062 10412 4068 10464
rect 4120 10412 4126 10464
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4304 10424 4353 10452
rect 4304 10412 4310 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5258 10452 5264 10464
rect 4580 10424 5264 10452
rect 4580 10412 4586 10424
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5442 10412 5448 10464
rect 5500 10412 5506 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8772 10452 8800 10492
rect 8849 10489 8861 10523
rect 8895 10520 8907 10523
rect 9508 10520 9536 10560
rect 10704 10520 10732 10696
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 11146 10616 11152 10668
rect 11204 10616 11210 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11790 10656 11796 10668
rect 11563 10628 11796 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11480 10560 11713 10588
rect 11480 10548 11486 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 13188 10588 13216 10619
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13320 10628 13461 10656
rect 13320 10616 13326 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10656 13691 10659
rect 13814 10656 13820 10668
rect 13679 10628 13820 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14274 10656 14280 10668
rect 14231 10628 14280 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 13188 10560 13676 10588
rect 12437 10551 12495 10557
rect 8895 10492 9536 10520
rect 9692 10492 10732 10520
rect 11333 10523 11391 10529
rect 8895 10489 8907 10492
rect 8849 10483 8907 10489
rect 9692 10452 9720 10492
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 12452 10520 12480 10551
rect 11379 10492 12480 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 12986 10480 12992 10532
rect 13044 10480 13050 10532
rect 13648 10464 13676 10560
rect 8772 10424 9720 10452
rect 9858 10412 9864 10464
rect 9916 10412 9922 10464
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12802 10452 12808 10464
rect 12207 10424 12808 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13630 10412 13636 10464
rect 13688 10412 13694 10464
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 1673 10251 1731 10257
rect 1673 10248 1685 10251
rect 1636 10220 1685 10248
rect 1636 10208 1642 10220
rect 1673 10217 1685 10220
rect 1719 10217 1731 10251
rect 1673 10211 1731 10217
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3602 10248 3608 10260
rect 3384 10220 3608 10248
rect 3384 10208 3390 10220
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4028 10220 4169 10248
rect 4028 10208 4034 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 5442 10248 5448 10260
rect 4157 10211 4215 10217
rect 5000 10220 5448 10248
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 4525 10183 4583 10189
rect 4525 10180 4537 10183
rect 4120 10152 4537 10180
rect 4120 10140 4126 10152
rect 4525 10149 4537 10152
rect 4571 10149 4583 10183
rect 4525 10143 4583 10149
rect 4632 10084 4936 10112
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 1964 9976 1992 10007
rect 2222 10004 2228 10056
rect 2280 10004 2286 10056
rect 3786 10004 3792 10056
rect 3844 10004 3850 10056
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 2498 9985 2504 9988
rect 1596 9948 1992 9976
rect 1596 9917 1624 9948
rect 2492 9939 2504 9985
rect 2498 9936 2504 9939
rect 2556 9936 2562 9988
rect 4632 9976 4660 10084
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 2746 9948 4660 9976
rect 4908 9976 4936 10084
rect 5000 10053 5028 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5905 10251 5963 10257
rect 5905 10217 5917 10251
rect 5951 10248 5963 10251
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 5951 10220 6285 10248
rect 5951 10217 5963 10220
rect 5905 10211 5963 10217
rect 6273 10217 6285 10220
rect 6319 10248 6331 10251
rect 7650 10248 7656 10260
rect 6319 10220 7656 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8662 10208 8668 10260
rect 8720 10208 8726 10260
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 11146 10208 11152 10260
rect 11204 10208 11210 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 11480 10220 11621 10248
rect 11480 10208 11486 10220
rect 11609 10217 11621 10220
rect 11655 10217 11667 10251
rect 11609 10211 11667 10217
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12526 10248 12532 10260
rect 12207 10220 12532 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12526 10208 12532 10220
rect 12584 10248 12590 10260
rect 12710 10248 12716 10260
rect 12584 10220 12716 10248
rect 12584 10208 12590 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13630 10248 13636 10260
rect 12820 10220 13636 10248
rect 5169 10183 5227 10189
rect 5169 10149 5181 10183
rect 5215 10180 5227 10183
rect 8680 10180 8708 10208
rect 5215 10152 5488 10180
rect 5215 10149 5227 10152
rect 5169 10143 5227 10149
rect 5460 10121 5488 10152
rect 7208 10152 8708 10180
rect 7208 10121 7236 10152
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7374 10072 7380 10124
rect 7432 10072 7438 10124
rect 8478 10112 8484 10124
rect 7944 10084 8484 10112
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5626 10044 5632 10056
rect 5307 10016 5632 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7944 10044 7972 10084
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9876 10112 9904 10208
rect 12820 10112 12848 10220
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14090 10208 14096 10260
rect 14148 10208 14154 10260
rect 9723 10084 9904 10112
rect 10152 10084 11376 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 6779 10016 7972 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8435 10016 8677 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8665 10013 8677 10016
rect 8711 10044 8723 10047
rect 8846 10044 8852 10056
rect 8711 10016 8852 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 4908 9948 7144 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2746 9908 2774 9948
rect 2087 9880 2774 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 5166 9908 5172 9920
rect 4396 9880 5172 9908
rect 4396 9868 4402 9880
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 7116 9908 7144 9948
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 7248 9948 7481 9976
rect 7248 9936 7254 9948
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 7469 9939 7527 9945
rect 7650 9936 7656 9988
rect 7708 9976 7714 9988
rect 8404 9976 8432 10007
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9324 10016 9505 10044
rect 7708 9948 8432 9976
rect 7708 9936 7714 9948
rect 8662 9908 8668 9920
rect 7116 9880 8668 9908
rect 8662 9868 8668 9880
rect 8720 9908 8726 9920
rect 9324 9908 9352 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10152 10044 10180 10084
rect 9916 10016 10180 10044
rect 9916 10004 9922 10016
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 11348 10053 11376 10084
rect 12268 10084 12848 10112
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10044 11391 10047
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11379 10016 11529 10044
rect 11379 10013 11391 10016
rect 11333 10007 11391 10013
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 10428 9976 10456 10007
rect 9416 9948 10456 9976
rect 9416 9917 9444 9948
rect 8720 9880 9352 9908
rect 9401 9911 9459 9917
rect 8720 9868 8726 9880
rect 9401 9877 9413 9911
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10192 9880 10885 9908
rect 10192 9868 10198 9880
rect 10873 9877 10885 9880
rect 10919 9877 10931 9911
rect 11532 9908 11560 10007
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 12268 10053 12296 10084
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 12253 10007 12311 10013
rect 12406 10016 13829 10044
rect 11624 9976 11652 10004
rect 12406 9976 12434 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13964 10016 14289 10044
rect 13964 10004 13970 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 11624 9948 12434 9976
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 13550 9979 13608 9985
rect 13550 9976 13562 9979
rect 13412 9948 13562 9976
rect 13412 9936 13418 9948
rect 13550 9945 13562 9948
rect 13596 9945 13608 9979
rect 13550 9939 13608 9945
rect 12158 9908 12164 9920
rect 11532 9880 12164 9908
rect 10873 9871 10931 9877
rect 12158 9868 12164 9880
rect 12216 9908 12222 9920
rect 12437 9911 12495 9917
rect 12437 9908 12449 9911
rect 12216 9880 12449 9908
rect 12216 9868 12222 9880
rect 12437 9877 12449 9880
rect 12483 9877 12495 9911
rect 12437 9871 12495 9877
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 2961 9707 3019 9713
rect 2961 9673 2973 9707
rect 3007 9704 3019 9707
rect 3234 9704 3240 9716
rect 3007 9676 3240 9704
rect 3007 9673 3019 9676
rect 2961 9667 3019 9673
rect 3234 9664 3240 9676
rect 3292 9704 3298 9716
rect 3786 9704 3792 9716
rect 3292 9676 3792 9704
rect 3292 9664 3298 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 3881 9707 3939 9713
rect 3881 9673 3893 9707
rect 3927 9704 3939 9707
rect 3970 9704 3976 9716
rect 3927 9676 3976 9704
rect 3927 9673 3939 9676
rect 3881 9667 3939 9673
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 5997 9707 6055 9713
rect 4080 9676 5856 9704
rect 4080 9636 4108 9676
rect 5718 9636 5724 9648
rect 1688 9608 4108 9636
rect 4172 9608 5724 9636
rect 1688 9577 1716 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 1912 9540 3249 9568
rect 1912 9528 1918 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 934 9460 940 9512
rect 992 9500 998 9512
rect 1397 9503 1455 9509
rect 1397 9500 1409 9503
rect 992 9472 1409 9500
rect 992 9460 998 9472
rect 1397 9469 1409 9472
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 2188 9472 2329 9500
rect 2188 9460 2194 9472
rect 2317 9469 2329 9472
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2547 9472 3157 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3252 9364 3280 9531
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3436 9432 3464 9531
rect 3384 9404 3464 9432
rect 3605 9435 3663 9441
rect 3384 9392 3390 9404
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 3712 9432 3740 9531
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4172 9577 4200 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 5828 9636 5856 9676
rect 5997 9673 6009 9707
rect 6043 9704 6055 9707
rect 6454 9704 6460 9716
rect 6043 9676 6460 9704
rect 6043 9673 6055 9676
rect 5997 9667 6055 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9673 6975 9707
rect 6917 9667 6975 9673
rect 7101 9707 7159 9713
rect 7101 9673 7113 9707
rect 7147 9704 7159 9707
rect 7466 9704 7472 9716
rect 7147 9676 7472 9704
rect 7147 9673 7159 9676
rect 7101 9667 7159 9673
rect 6932 9636 6960 9667
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 8754 9704 8760 9716
rect 8435 9676 8760 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 9272 9676 9597 9704
rect 9272 9664 9278 9676
rect 9585 9673 9597 9676
rect 9631 9673 9643 9707
rect 9585 9667 9643 9673
rect 10045 9707 10103 9713
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10226 9704 10232 9716
rect 10091 9676 10232 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 12897 9707 12955 9713
rect 12897 9673 12909 9707
rect 12943 9673 12955 9707
rect 12897 9667 12955 9673
rect 5828 9608 6040 9636
rect 6932 9608 9352 9636
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3936 9540 4077 9568
rect 3936 9528 3942 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4341 9531 4399 9537
rect 4540 9540 4629 9568
rect 3651 9404 3740 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 4154 9364 4160 9376
rect 3252 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9364 4218 9376
rect 4356 9364 4384 9531
rect 4540 9441 4568 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5442 9568 5448 9580
rect 4939 9540 5448 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 4908 9500 4936 9531
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 4632 9472 4936 9500
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9401 4583 9435
rect 4525 9395 4583 9401
rect 4632 9364 4660 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 5132 9472 5181 9500
rect 5132 9460 5138 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 4801 9435 4859 9441
rect 4801 9401 4813 9435
rect 4847 9432 4859 9435
rect 5368 9432 5396 9463
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5684 9472 5825 9500
rect 5684 9460 5690 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 4847 9404 5396 9432
rect 6012 9432 6040 9608
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6748 9500 6776 9531
rect 7006 9528 7012 9580
rect 7064 9528 7070 9580
rect 7653 9571 7711 9577
rect 7116 9540 7604 9568
rect 7116 9500 7144 9540
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 6748 9472 7144 9500
rect 7300 9472 7481 9500
rect 6012 9404 7236 9432
rect 4847 9401 4859 9404
rect 4801 9395 4859 9401
rect 7208 9376 7236 9404
rect 7300 9376 7328 9472
rect 7469 9469 7481 9472
rect 7515 9469 7527 9503
rect 7576 9500 7604 9540
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 8386 9568 8392 9580
rect 7699 9540 8392 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 9324 9577 9352 9608
rect 9858 9596 9864 9648
rect 9916 9596 9922 9648
rect 12912 9636 12940 9667
rect 13906 9664 13912 9716
rect 13964 9664 13970 9716
rect 13924 9636 13952 9664
rect 12452 9608 12848 9636
rect 12912 9608 13952 9636
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8588 9540 9045 9568
rect 8113 9503 8171 9509
rect 7576 9472 7696 9500
rect 7469 9463 7527 9469
rect 7668 9444 7696 9472
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 8496 9500 8524 9528
rect 8159 9472 8524 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 7650 9392 7656 9444
rect 7708 9392 7714 9444
rect 8588 9376 8616 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9876 9568 9904 9596
rect 9815 9540 9904 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 10192 9540 10241 9568
rect 10192 9528 10198 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 8864 9432 8892 9463
rect 10410 9460 10416 9512
rect 10468 9460 10474 9512
rect 11716 9500 11744 9531
rect 12158 9528 12164 9580
rect 12216 9528 12222 9580
rect 12452 9577 12480 9608
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12676 9540 12725 9568
rect 12676 9528 12682 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12820 9568 12848 9608
rect 12820 9540 13952 9568
rect 12713 9531 12771 9537
rect 13924 9512 13952 9540
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 14056 9540 14381 9568
rect 14056 9528 14062 9540
rect 14369 9537 14381 9540
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 12526 9500 12532 9512
rect 11716 9472 12532 9500
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13446 9460 13452 9512
rect 13504 9460 13510 9512
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13596 9472 13645 9500
rect 13596 9460 13602 9472
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 9125 9435 9183 9441
rect 9125 9432 9137 9435
rect 8864 9404 9137 9432
rect 9125 9401 9137 9404
rect 9171 9401 9183 9435
rect 9125 9395 9183 9401
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 14200 9432 14228 9463
rect 12299 9404 14228 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 4212 9336 4660 9364
rect 4212 9324 4218 9336
rect 4982 9324 4988 9376
rect 5040 9324 5046 9376
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5810 9364 5816 9376
rect 5316 9336 5816 9364
rect 5316 9324 5322 9336
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6454 9364 6460 9376
rect 6411 9336 6460 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7190 9324 7196 9376
rect 7248 9324 7254 9376
rect 7282 9324 7288 9376
rect 7340 9324 7346 9376
rect 8570 9324 8576 9376
rect 8628 9324 8634 9376
rect 10686 9324 10692 9376
rect 10744 9324 10750 9376
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 12618 9324 12624 9376
rect 12676 9324 12682 9376
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 13725 9367 13783 9373
rect 13725 9364 13737 9367
rect 13320 9336 13737 9364
rect 13320 9324 13326 9336
rect 13725 9333 13737 9336
rect 13771 9333 13783 9367
rect 13725 9327 13783 9333
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 3234 9160 3240 9172
rect 2179 9132 3240 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3418 9120 3424 9172
rect 3476 9120 3482 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4706 9160 4712 9172
rect 3936 9132 4712 9160
rect 3936 9120 3942 9132
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5626 9120 5632 9172
rect 5684 9120 5690 9172
rect 6454 9120 6460 9172
rect 6512 9120 6518 9172
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 8297 9163 8355 9169
rect 7248 9132 7420 9160
rect 7248 9120 7254 9132
rect 3050 9092 3056 9104
rect 2516 9064 3056 9092
rect 2516 9033 2544 9064
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9061 3203 9095
rect 3145 9055 3203 9061
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 8993 2559 9027
rect 3160 9024 3188 9055
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3384 9064 3801 9092
rect 3384 9052 3390 9064
rect 3789 9061 3801 9064
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 4154 9024 4160 9036
rect 2501 8987 2559 8993
rect 2792 8996 3188 9024
rect 3344 8996 4160 9024
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 2792 8965 2820 8996
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2777 8959 2835 8965
rect 2363 8928 2636 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 2130 8820 2136 8832
rect 1719 8792 2136 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 2608 8829 2636 8928
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 2884 8888 2912 8919
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3344 8965 3372 8996
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 5000 9024 5028 9120
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 5316 9064 6316 9092
rect 5316 9052 5322 9064
rect 5353 9027 5411 9033
rect 5353 9024 5365 9027
rect 5000 8996 5365 9024
rect 5353 8993 5365 8996
rect 5399 8993 5411 9027
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 5353 8987 5411 8993
rect 5460 8996 6193 9024
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3292 8928 3341 8956
rect 3292 8916 3298 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3602 8916 3608 8968
rect 3660 8916 3666 8968
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 4706 8956 4712 8968
rect 4663 8928 4712 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 4338 8888 4344 8900
rect 2740 8860 2912 8888
rect 3988 8860 4344 8888
rect 2740 8848 2746 8860
rect 3988 8832 4016 8860
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8820 3019 8823
rect 3510 8820 3516 8832
rect 3007 8792 3516 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 4908 8820 4936 8916
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5460 8888 5488 8996
rect 6181 8993 6193 8996
rect 6227 8993 6239 9027
rect 6181 8987 6239 8993
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6288 8956 6316 9064
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6472 9024 6500 9120
rect 6825 9095 6883 9101
rect 6825 9061 6837 9095
rect 6871 9092 6883 9095
rect 7282 9092 7288 9104
rect 6871 9064 7288 9092
rect 6871 9061 6883 9064
rect 6825 9055 6883 9061
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7392 9092 7420 9132
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8754 9160 8760 9172
rect 8343 9132 8760 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 10505 9163 10563 9169
rect 10505 9160 10517 9163
rect 10468 9132 10517 9160
rect 10468 9120 10474 9132
rect 10505 9129 10517 9132
rect 10551 9129 10563 9163
rect 10505 9123 10563 9129
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 11940 9132 13400 9160
rect 11940 9120 11946 9132
rect 10318 9092 10324 9104
rect 7392 9064 10324 9092
rect 6411 8996 6500 9024
rect 7837 9027 7895 9033
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 7837 8993 7849 9027
rect 7883 9024 7895 9027
rect 8294 9024 8300 9036
rect 7883 8996 8300 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9272 8996 9597 9024
rect 9272 8984 9278 8996
rect 9585 8993 9597 8996
rect 9631 9024 9643 9027
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 9631 8996 9781 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6288 8928 6929 8956
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 5040 8860 5488 8888
rect 5997 8891 6055 8897
rect 5040 8848 5046 8860
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 7116 8888 7144 8919
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 9876 8965 9904 9064
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 11146 9052 11152 9104
rect 11204 9092 11210 9104
rect 11425 9095 11483 9101
rect 11425 9092 11437 9095
rect 11204 9064 11437 9092
rect 11204 9052 11210 9064
rect 11425 9061 11437 9064
rect 11471 9092 11483 9095
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 11471 9064 11713 9092
rect 11471 9061 11483 9064
rect 11425 9055 11483 9061
rect 11701 9061 11713 9064
rect 11747 9061 11759 9095
rect 11701 9055 11759 9061
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12216 8996 12480 9024
rect 12216 8984 12222 8996
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8444 8928 9413 8956
rect 8444 8916 8450 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10244 8928 10333 8956
rect 9122 8888 9128 8900
rect 6043 8860 7144 8888
rect 8312 8860 9128 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 5166 8820 5172 8832
rect 4908 8792 5172 8820
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 8312 8820 8340 8860
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 6512 8792 8340 8820
rect 6512 8780 6518 8792
rect 8386 8780 8392 8832
rect 8444 8780 8450 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 10244 8829 10272 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 12452 8956 12480 8996
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 13372 9033 13400 9132
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13998 9160 14004 9172
rect 13504 9132 14004 9160
rect 13504 9120 13510 9132
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 14240 9132 14289 9160
rect 14240 9120 14246 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 12860 8996 13185 9024
rect 12860 8984 12866 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12452 8928 13093 8956
rect 10321 8919 10379 8925
rect 13081 8925 13093 8928
rect 13127 8956 13139 8959
rect 13446 8956 13452 8968
rect 13127 8928 13452 8956
rect 13127 8925 13139 8928
rect 13081 8919 13139 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 14182 8956 14188 8968
rect 14139 8928 14188 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8628 8792 8953 8820
rect 8628 8780 8634 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 10229 8823 10287 8829
rect 10229 8789 10241 8823
rect 10275 8789 10287 8823
rect 10229 8783 10287 8789
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 10888 8820 10916 8851
rect 10962 8848 10968 8900
rect 11020 8848 11026 8900
rect 12158 8848 12164 8900
rect 12216 8848 12222 8900
rect 12253 8891 12311 8897
rect 12253 8857 12265 8891
rect 12299 8888 12311 8891
rect 13817 8891 13875 8897
rect 13817 8888 13829 8891
rect 12299 8860 13829 8888
rect 12299 8857 12311 8860
rect 12253 8851 12311 8857
rect 13817 8857 13829 8860
rect 13863 8857 13875 8891
rect 13817 8851 13875 8857
rect 10744 8792 10916 8820
rect 10744 8780 10750 8792
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12268 8820 12296 8851
rect 11848 8792 12296 8820
rect 11848 8780 11854 8792
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 14550 8820 14556 8832
rect 12676 8792 14556 8820
rect 12676 8780 12682 8792
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2556 8588 2973 8616
rect 2556 8576 2562 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 2961 8579 3019 8585
rect 3620 8588 3832 8616
rect 3620 8548 3648 8588
rect 2884 8520 3648 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2314 8480 2320 8492
rect 1719 8452 2320 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2406 8440 2412 8492
rect 2464 8440 2470 8492
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2731 8452 2820 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2372 8316 2728 8344
rect 2372 8304 2378 8316
rect 2700 8288 2728 8316
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2556 8248 2605 8276
rect 2556 8236 2562 8248
rect 2593 8245 2605 8248
rect 2639 8245 2651 8279
rect 2593 8239 2651 8245
rect 2682 8236 2688 8288
rect 2740 8236 2746 8288
rect 2792 8276 2820 8452
rect 2884 8353 2912 8520
rect 3694 8508 3700 8560
rect 3752 8508 3758 8560
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 3712 8421 3740 8508
rect 3804 8480 3832 8588
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4212 8588 4353 8616
rect 4212 8576 4218 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4706 8616 4712 8628
rect 4663 8588 4712 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6178 8616 6184 8628
rect 6043 8588 6184 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6546 8576 6552 8628
rect 6604 8576 6610 8628
rect 6914 8576 6920 8628
rect 6972 8576 6978 8628
rect 8294 8576 8300 8628
rect 8352 8576 8358 8628
rect 8386 8576 8392 8628
rect 8444 8576 8450 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9858 8616 9864 8628
rect 9646 8588 9864 8616
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 5868 8520 6040 8548
rect 5868 8508 5874 8520
rect 4433 8483 4491 8489
rect 4433 8480 4445 8483
rect 3804 8452 4445 8480
rect 4433 8449 4445 8452
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4847 8452 5181 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3292 8384 3525 8412
rect 3292 8372 3298 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3878 8372 3884 8424
rect 3936 8372 3942 8424
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8313 2927 8347
rect 3786 8344 3792 8356
rect 2869 8307 2927 8313
rect 2976 8316 3792 8344
rect 2976 8276 3004 8316
rect 3786 8304 3792 8316
rect 3844 8344 3850 8356
rect 4724 8344 4752 8443
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6012 8480 6040 8520
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6932 8548 6960 8576
rect 7745 8551 7803 8557
rect 6144 8520 7696 8548
rect 6144 8508 6150 8520
rect 6380 8489 6408 8520
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 6012 8452 6193 8480
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 6932 8480 6960 8520
rect 7668 8489 7696 8520
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 8312 8548 8340 8576
rect 7791 8520 8340 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6932 8452 7113 8480
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7101 8443 7159 8449
rect 7300 8452 7389 8480
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 5368 8344 5396 8440
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 7300 8353 7328 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7834 8480 7840 8492
rect 7699 8452 7840 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8404 8480 8432 8576
rect 7975 8452 8432 8480
rect 9493 8483 9551 8489
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9646 8480 9674 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 11020 8588 11069 8616
rect 11020 8576 11026 8588
rect 11057 8585 11069 8588
rect 11103 8585 11115 8619
rect 11057 8579 11115 8585
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 13354 8616 13360 8628
rect 12676 8588 13360 8616
rect 12676 8576 12682 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 14274 8576 14280 8628
rect 14332 8576 14338 8628
rect 10042 8508 10048 8560
rect 10100 8508 10106 8560
rect 12820 8520 13492 8548
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9539 8452 9781 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 10060 8480 10088 8508
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 10060 8452 10977 8480
rect 9769 8443 9827 8449
rect 10965 8449 10977 8452
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8480 11299 8483
rect 11701 8483 11759 8489
rect 11287 8452 11560 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 3844 8316 5028 8344
rect 5368 8316 6653 8344
rect 3844 8304 3850 8316
rect 2792 8248 3004 8276
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 4890 8276 4896 8288
rect 3200 8248 4896 8276
rect 3200 8236 3206 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5000 8276 5028 8316
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 6641 8307 6699 8313
rect 7285 8347 7343 8353
rect 7285 8313 7297 8347
rect 7331 8313 7343 8347
rect 7285 8307 7343 8313
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 8128 8344 8156 8375
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 10008 8384 10057 8412
rect 10008 8372 10014 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10045 8375 10103 8381
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10275 8384 10885 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 10873 8381 10885 8384
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 7607 8316 8156 8344
rect 9677 8347 9735 8353
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 9858 8344 9864 8356
rect 9723 8316 9864 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 11532 8353 11560 8452
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 12066 8480 12072 8492
rect 11747 8452 12072 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12299 8452 12633 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 12820 8489 12848 8520
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 12943 8452 13369 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 13357 8449 13369 8452
rect 13403 8449 13415 8483
rect 13464 8480 13492 8520
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13872 8520 14228 8548
rect 13872 8508 13878 8520
rect 13722 8480 13728 8492
rect 13464 8452 13728 8480
rect 13357 8443 13415 8449
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 14200 8489 14228 8520
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13780 8452 13921 8480
rect 13780 8440 13786 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 11790 8304 11796 8356
rect 11848 8344 11854 8356
rect 12250 8344 12256 8356
rect 11848 8316 12256 8344
rect 11848 8304 11854 8316
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 12452 8344 12480 8375
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 13044 8384 13185 8412
rect 13044 8372 13050 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13262 8372 13268 8424
rect 13320 8372 13326 8424
rect 13280 8344 13308 8372
rect 12452 8316 13308 8344
rect 8386 8276 8392 8288
rect 5000 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 9180 8248 9321 8276
rect 9180 8236 9186 8248
rect 9309 8245 9321 8248
rect 9355 8245 9367 8279
rect 9309 8239 9367 8245
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 13538 8276 13544 8288
rect 13412 8248 13544 8276
rect 13412 8236 13418 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 14090 8236 14096 8288
rect 14148 8236 14154 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 3513 8075 3571 8081
rect 2464 8044 3464 8072
rect 2464 8032 2470 8044
rect 3436 8004 3464 8044
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3878 8072 3884 8084
rect 3559 8044 3884 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5258 8072 5264 8084
rect 5123 8044 5264 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10100 8044 12112 8072
rect 10100 8032 10106 8044
rect 4617 8007 4675 8013
rect 4617 8004 4629 8007
rect 3436 7976 4629 8004
rect 4617 7973 4629 7976
rect 4663 7973 4675 8007
rect 4617 7967 4675 7973
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 5552 7936 5580 8032
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 8113 8007 8171 8013
rect 8113 8004 8125 8007
rect 7432 7976 8125 8004
rect 7432 7964 7438 7976
rect 8113 7973 8125 7976
rect 8159 7973 8171 8007
rect 8113 7967 8171 7973
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 3099 7908 5580 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 3068 7868 3096 7899
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 9140 7936 9168 7967
rect 12084 7945 12112 8044
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12216 8044 12357 8072
rect 12216 8032 12222 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 12526 8032 12532 8084
rect 12584 8032 12590 8084
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 14458 8072 14464 8084
rect 13596 8044 14464 8072
rect 13596 8032 13602 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 7064 7908 8340 7936
rect 9140 7908 9413 7936
rect 7064 7896 7070 7908
rect 2280 7840 3096 7868
rect 2280 7828 2286 7840
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3694 7868 3700 7880
rect 3467 7840 3700 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4890 7868 4896 7880
rect 4847 7840 4896 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 6454 7868 6460 7880
rect 5031 7840 6460 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 2808 7803 2866 7809
rect 2808 7769 2820 7803
rect 2854 7800 2866 7803
rect 3050 7800 3056 7812
rect 2854 7772 3056 7800
rect 2854 7769 2866 7772
rect 2808 7763 2866 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 3160 7732 3188 7828
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 4341 7803 4399 7809
rect 3283 7772 3740 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 1719 7704 3188 7732
rect 3712 7732 3740 7772
rect 4341 7769 4353 7803
rect 4387 7769 4399 7803
rect 4341 7763 4399 7769
rect 4356 7732 4384 7763
rect 4430 7760 4436 7812
rect 4488 7760 4494 7812
rect 5000 7800 5028 7831
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6604 7840 7113 7868
rect 6604 7828 6610 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7708 7840 7757 7868
rect 7708 7828 7714 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7892 7840 8033 7868
rect 7892 7828 7898 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8312 7877 8340 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 12115 7908 12756 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12728 7880 12756 7908
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9122 7868 9128 7880
rect 8987 7840 9128 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11606 7868 11612 7880
rect 11471 7840 11612 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 12216 7840 12265 7868
rect 12216 7828 12222 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13504 7840 13553 7868
rect 13504 7828 13510 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 14148 7840 14289 7868
rect 14148 7828 14154 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 4908 7772 5028 7800
rect 7009 7803 7067 7809
rect 4908 7744 4936 7772
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 8220 7800 8248 7828
rect 9232 7800 9260 7828
rect 7055 7772 8248 7800
rect 8956 7772 9260 7800
rect 11180 7803 11238 7809
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 8956 7744 8984 7772
rect 11180 7769 11192 7803
rect 11226 7800 11238 7803
rect 12434 7800 12440 7812
rect 11226 7772 12440 7800
rect 11226 7769 11238 7772
rect 11180 7763 11238 7769
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 14182 7800 14188 7812
rect 13740 7772 14188 7800
rect 3712 7704 4384 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 4890 7692 4896 7744
rect 4948 7692 4954 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7524 7704 7849 7732
rect 7524 7692 7530 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7732 9919 7735
rect 9950 7732 9956 7744
rect 9907 7704 9956 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 10928 7704 11529 7732
rect 10928 7692 10934 7704
rect 11517 7701 11529 7704
rect 11563 7701 11575 7735
rect 11517 7695 11575 7701
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 13740 7741 13768 7772
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7701 13783 7735
rect 13725 7695 13783 7701
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 2314 7528 2320 7540
rect 1443 7500 2320 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2556 7500 3096 7528
rect 2556 7488 2562 7500
rect 2222 7420 2228 7472
rect 2280 7460 2286 7472
rect 3068 7469 3096 7500
rect 3510 7488 3516 7540
rect 3568 7488 3574 7540
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 4890 7528 4896 7540
rect 3936 7500 4896 7528
rect 3936 7488 3942 7500
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 3053 7463 3111 7469
rect 2280 7432 2820 7460
rect 2280 7420 2286 7432
rect 2792 7401 2820 7432
rect 3053 7429 3065 7463
rect 3099 7429 3111 7463
rect 3528 7460 3556 7488
rect 3528 7432 4660 7460
rect 3053 7423 3111 7429
rect 2521 7395 2579 7401
rect 2521 7361 2533 7395
rect 2567 7392 2579 7395
rect 2777 7395 2835 7401
rect 2567 7364 2728 7392
rect 2567 7361 2579 7364
rect 2521 7355 2579 7361
rect 2700 7324 2728 7364
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 3786 7392 3792 7404
rect 3651 7364 3792 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4632 7401 4660 7432
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 5810 7392 5816 7404
rect 4617 7355 4675 7361
rect 5552 7364 5816 7392
rect 2961 7327 3019 7333
rect 2700 7296 2912 7324
rect 2884 7256 2912 7296
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3234 7324 3240 7336
rect 3007 7296 3240 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 5552 7324 5580 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6380 7392 6408 7491
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7282 7528 7288 7540
rect 6963 7500 7288 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7466 7488 7472 7540
rect 7524 7488 7530 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 12158 7528 12164 7540
rect 11287 7500 12164 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 6840 7460 6868 7488
rect 6564 7432 6868 7460
rect 6564 7401 6592 7432
rect 6043 7364 6408 7392
rect 6549 7395 6607 7401
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6914 7392 6920 7404
rect 6871 7364 6920 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7484 7401 7512 7488
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8202 7460 8208 7472
rect 7883 7432 8208 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 9631 7432 11652 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 9876 7401 9904 7432
rect 11624 7404 11652 7432
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7248 7364 7297 7392
rect 7248 7352 7254 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10128 7395 10186 7401
rect 10128 7361 10140 7395
rect 10174 7392 10186 7395
rect 10870 7392 10876 7404
rect 10174 7364 10876 7392
rect 10174 7361 10186 7364
rect 10128 7355 10186 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11606 7352 11612 7404
rect 11664 7352 11670 7404
rect 12084 7401 12112 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12986 7528 12992 7540
rect 12667 7500 12992 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7497 13139 7531
rect 13081 7491 13139 7497
rect 13096 7460 13124 7491
rect 13354 7488 13360 7540
rect 13412 7488 13418 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 14182 7488 14188 7540
rect 14240 7488 14246 7540
rect 12406 7432 13124 7460
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12406 7392 12434 7432
rect 12299 7364 12434 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 12989 7395 13047 7401
rect 12584 7364 12848 7392
rect 12584 7352 12590 7364
rect 12820 7336 12848 7364
rect 12989 7361 13001 7395
rect 13035 7390 13047 7395
rect 13035 7362 13124 7390
rect 13035 7361 13047 7362
rect 12989 7355 13047 7361
rect 4387 7296 5580 7324
rect 5721 7327 5779 7333
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6454 7324 6460 7336
rect 5951 7296 6460 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 3142 7256 3148 7268
rect 2884 7228 3148 7256
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 5261 7259 5319 7265
rect 5261 7256 5273 7259
rect 4172 7228 5273 7256
rect 4172 7200 4200 7228
rect 5261 7225 5273 7228
rect 5307 7256 5319 7259
rect 5626 7256 5632 7268
rect 5307 7228 5632 7256
rect 5307 7225 5319 7228
rect 5261 7219 5319 7225
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 5736 7256 5764 7287
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 12802 7284 12808 7336
rect 12860 7284 12866 7336
rect 13096 7324 13124 7362
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 13228 7364 13277 7392
rect 13228 7352 13234 7364
rect 13265 7361 13277 7364
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 14108 7392 14136 7488
rect 13863 7364 14136 7392
rect 14200 7392 14228 7488
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 14200 7364 14289 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14001 7327 14059 7333
rect 13096 7296 13768 7324
rect 7101 7259 7159 7265
rect 7101 7256 7113 7259
rect 5736 7228 7113 7256
rect 7101 7225 7113 7228
rect 7147 7225 7159 7259
rect 7101 7219 7159 7225
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 11517 7259 11575 7265
rect 11517 7256 11529 7259
rect 11204 7228 11529 7256
rect 11204 7216 11210 7228
rect 11517 7225 11529 7228
rect 11563 7225 11575 7259
rect 12820 7256 12848 7284
rect 13170 7256 13176 7268
rect 12820 7228 13176 7256
rect 11517 7219 11575 7225
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 13740 7200 13768 7296
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14366 7324 14372 7336
rect 14047 7296 14372 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 2406 7148 2412 7200
rect 2464 7188 2470 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 2464 7160 3709 7188
rect 2464 7148 2470 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 4154 7148 4160 7200
rect 4212 7148 4218 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4304 7160 4813 7188
rect 4304 7148 4310 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 4801 7151 4859 7157
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6454 7188 6460 7200
rect 6227 7160 6460 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7653 7191 7711 7197
rect 7653 7157 7665 7191
rect 7699 7188 7711 7191
rect 8294 7188 8300 7200
rect 7699 7160 8300 7188
rect 7699 7157 7711 7160
rect 7653 7151 7711 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 12434 7148 12440 7200
rect 12492 7148 12498 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13630 7188 13636 7200
rect 12851 7160 13636 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13722 7148 13728 7200
rect 13780 7148 13786 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 14056 7160 14105 7188
rect 14056 7148 14062 7160
rect 14093 7157 14105 7160
rect 14139 7157 14151 7191
rect 14093 7151 14151 7157
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 3050 6944 3056 6996
rect 3108 6944 3114 6996
rect 4246 6944 4252 6996
rect 4304 6944 4310 6996
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 5902 6984 5908 6996
rect 5684 6956 5908 6984
rect 5684 6944 5690 6956
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7708 6956 7849 6984
rect 7708 6944 7714 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 9769 6987 9827 6993
rect 9769 6953 9781 6987
rect 9815 6984 9827 6987
rect 9950 6984 9956 6996
rect 9815 6956 9956 6984
rect 9815 6953 9827 6956
rect 9769 6947 9827 6953
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 13446 6944 13452 6996
rect 13504 6944 13510 6996
rect 3510 6876 3516 6928
rect 3568 6916 3574 6928
rect 8478 6916 8484 6928
rect 3568 6888 8484 6916
rect 3568 6876 3574 6888
rect 8478 6876 8484 6888
rect 8536 6876 8542 6928
rect 10321 6919 10379 6925
rect 10321 6885 10333 6919
rect 10367 6885 10379 6919
rect 10321 6879 10379 6885
rect 934 6808 940 6860
rect 992 6848 998 6860
rect 1397 6851 1455 6857
rect 1397 6848 1409 6851
rect 992 6820 1409 6848
rect 992 6808 998 6820
rect 1397 6817 1409 6820
rect 1443 6817 1455 6851
rect 1397 6811 1455 6817
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 2314 6808 2320 6860
rect 2372 6848 2378 6860
rect 2409 6851 2467 6857
rect 2409 6848 2421 6851
rect 2372 6820 2421 6848
rect 2372 6808 2378 6820
rect 2409 6817 2421 6820
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 3835 6820 4660 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 2556 6752 3341 6780
rect 2556 6740 2562 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 3988 6712 4016 6743
rect 4632 6721 4660 6820
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6848 6423 6851
rect 6454 6848 6460 6860
rect 6411 6820 6460 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6696 6820 6837 6848
rect 6696 6808 6702 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 7098 6808 7104 6860
rect 7156 6808 7162 6860
rect 8294 6808 8300 6860
rect 8352 6808 8358 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8496 6820 9137 6848
rect 5074 6740 5080 6792
rect 5132 6740 5138 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5960 6752 6009 6780
rect 5960 6740 5966 6752
rect 5997 6749 6009 6752
rect 6043 6780 6055 6783
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 6043 6752 6193 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 7282 6740 7288 6792
rect 7340 6740 7346 6792
rect 8496 6789 8524 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9858 6848 9864 6860
rect 9355 6820 9864 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10336 6848 10364 6879
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 11333 6919 11391 6925
rect 11333 6916 11345 6919
rect 10836 6888 11345 6916
rect 10836 6876 10842 6888
rect 11333 6885 11345 6888
rect 11379 6885 11391 6919
rect 12618 6916 12624 6928
rect 11333 6879 11391 6885
rect 12360 6888 12624 6916
rect 11054 6848 11060 6860
rect 10336 6820 11060 6848
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11790 6848 11796 6860
rect 11532 6820 11796 6848
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8404 6752 8493 6780
rect 3528 6684 4016 6712
rect 4617 6715 4675 6721
rect 3528 6653 3556 6684
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4663 6684 5365 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 8404 6656 8432 6752
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8597 6783 8655 6789
rect 8597 6749 8609 6783
rect 8643 6780 8655 6783
rect 8754 6780 8760 6792
rect 8643 6752 8760 6780
rect 8643 6749 8655 6752
rect 8597 6743 8655 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10410 6780 10416 6792
rect 10183 6752 10416 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10870 6780 10876 6792
rect 10735 6752 10876 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 11532 6789 11560 6820
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 11882 6808 11888 6860
rect 11940 6808 11946 6860
rect 12360 6848 12388 6888
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 11992 6820 12388 6848
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6780 11667 6783
rect 11698 6780 11704 6792
rect 11655 6752 11704 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 10980 6712 11008 6743
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11992 6712 12020 6820
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 12492 6820 13645 6848
rect 12492 6808 12498 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 13863 6820 14412 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 14384 6792 14412 6820
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12115 6752 12725 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13262 6780 13268 6792
rect 12943 6752 13268 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14292 6712 14320 6743
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 10336 6684 11008 6712
rect 11716 6684 12020 6712
rect 12406 6684 14320 6712
rect 10336 6656 10364 6684
rect 3513 6647 3571 6653
rect 3513 6613 3525 6647
rect 3559 6613 3571 6647
rect 3513 6607 3571 6613
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5442 6644 5448 6656
rect 5040 6616 5448 6644
rect 5040 6604 5046 6616
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 6822 6644 6828 6656
rect 5500 6616 6828 6644
rect 5500 6604 5506 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7708 6616 7757 6644
rect 7708 6604 7714 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8444 6616 8677 6644
rect 8444 6604 8450 6616
rect 8665 6613 8677 6616
rect 8711 6613 8723 6647
rect 8665 6607 8723 6613
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10226 6644 10232 6656
rect 9999 6616 10232 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10318 6604 10324 6656
rect 10376 6604 10382 6656
rect 10502 6604 10508 6656
rect 10560 6604 10566 6656
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 11716 6644 11744 6684
rect 10919 6616 11744 6644
rect 11793 6647 11851 6653
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 12406 6644 12434 6684
rect 11839 6616 12434 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12526 6604 12532 6656
rect 12584 6604 12590 6656
rect 13081 6647 13139 6653
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13814 6644 13820 6656
rect 13127 6616 13820 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13964 6616 14105 6644
rect 13964 6604 13970 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2498 6440 2504 6452
rect 1995 6412 2504 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 3142 6440 3148 6452
rect 2823 6412 3148 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3694 6400 3700 6452
rect 3752 6400 3758 6452
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 5074 6440 5080 6452
rect 4111 6412 5080 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5810 6440 5816 6452
rect 5184 6412 5816 6440
rect 2314 6372 2320 6384
rect 1780 6344 2320 6372
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1780 6313 1808 6344
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 3234 6372 3240 6384
rect 2731 6344 3240 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3712 6372 3740 6400
rect 4249 6375 4307 6381
rect 3712 6344 4200 6372
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1544 6276 1777 6304
rect 1544 6264 1550 6276
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 3421 6307 3479 6313
rect 2087 6276 2452 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2424 6248 2452 6276
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 3467 6276 3617 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3605 6273 3617 6276
rect 3651 6304 3663 6307
rect 3712 6304 3740 6344
rect 4172 6313 4200 6344
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 5184 6372 5212 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6638 6440 6644 6452
rect 6411 6412 6644 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6409 10011 6443
rect 9953 6403 10011 6409
rect 10612 6412 11836 6440
rect 4295 6344 5212 6372
rect 5552 6344 6224 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 5552 6316 5580 6344
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 3651 6276 3740 6304
rect 3804 6276 3893 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 2222 6196 2228 6248
rect 2280 6196 2286 6248
rect 2406 6196 2412 6248
rect 2464 6196 2470 6248
rect 3804 6177 3832 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4203 6276 4445 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 6196 6313 6224 6344
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 9968 6372 9996 6403
rect 10612 6384 10640 6412
rect 6512 6344 9996 6372
rect 6512 6332 6518 6344
rect 8680 6313 8708 6344
rect 10594 6332 10600 6384
rect 10652 6332 10658 6384
rect 11146 6372 11152 6384
rect 11072 6344 11152 6372
rect 5925 6307 5983 6313
rect 5925 6273 5937 6307
rect 5971 6304 5983 6307
rect 6181 6307 6239 6313
rect 5971 6276 6132 6304
rect 5971 6273 5983 6276
rect 5925 6267 5983 6273
rect 6104 6236 6132 6276
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 6181 6267 6239 6273
rect 6288 6276 8033 6304
rect 6288 6236 6316 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 11072 6313 11100 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 11698 6372 11704 6384
rect 11296 6344 11704 6372
rect 11296 6332 11302 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 11808 6372 11836 6412
rect 13446 6400 13452 6452
rect 13504 6400 13510 6452
rect 11974 6372 11980 6384
rect 11808 6344 11980 6372
rect 11974 6332 11980 6344
rect 12032 6372 12038 6384
rect 12032 6344 12296 6372
rect 12032 6332 12038 6344
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9272 6276 9689 6304
rect 9272 6264 9278 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 11066 6307 11124 6313
rect 11066 6273 11078 6307
rect 11112 6273 11124 6307
rect 11066 6267 11124 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11606 6304 11612 6316
rect 11379 6276 11612 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11606 6264 11612 6276
rect 11664 6304 11670 6316
rect 12268 6304 12296 6344
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 12768 6344 13001 6372
rect 12768 6332 12774 6344
rect 12989 6341 13001 6344
rect 13035 6341 13047 6375
rect 13464 6372 13492 6400
rect 12989 6335 13047 6341
rect 13280 6344 13492 6372
rect 13280 6313 13308 6344
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11664 6276 12204 6304
rect 12268 6276 12449 6304
rect 11664 6264 11670 6276
rect 12176 6248 12204 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13446 6264 13452 6316
rect 13504 6264 13510 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 6104 6208 6316 6236
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 3789 6171 3847 6177
rect 3789 6137 3801 6171
rect 3835 6137 3847 6171
rect 3789 6131 3847 6137
rect 4617 6171 4675 6177
rect 4617 6137 4629 6171
rect 4663 6168 4675 6171
rect 4663 6140 5304 6168
rect 4663 6137 4675 6140
rect 4617 6131 4675 6137
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 1854 6100 1860 6112
rect 1627 6072 1860 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 4982 6100 4988 6112
rect 4847 6072 4988 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5276 6100 5304 6140
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 7024 6168 7052 6199
rect 7190 6196 7196 6248
rect 7248 6196 7254 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8386 6236 8392 6248
rect 7975 6208 8392 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 6696 6140 7052 6168
rect 6696 6128 6702 6140
rect 7208 6100 7236 6196
rect 7760 6168 7788 6199
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 11440 6208 11529 6236
rect 9769 6171 9827 6177
rect 9769 6168 9781 6171
rect 7760 6140 9781 6168
rect 9769 6137 9781 6140
rect 9815 6137 9827 6171
rect 9769 6131 9827 6137
rect 5276 6072 7236 6100
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 9306 6100 9312 6112
rect 7607 6072 9312 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11440 6100 11468 6208
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6236 13139 6239
rect 13354 6236 13360 6248
rect 13127 6208 13360 6236
rect 13127 6205 13139 6208
rect 13081 6199 13139 6205
rect 13354 6196 13360 6208
rect 13412 6236 13418 6248
rect 13412 6208 13676 6236
rect 13412 6196 13418 6208
rect 11885 6171 11943 6177
rect 11885 6168 11897 6171
rect 11532 6140 11897 6168
rect 11532 6112 11560 6140
rect 11885 6137 11897 6140
rect 11931 6168 11943 6171
rect 12618 6168 12624 6180
rect 11931 6140 12624 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 13648 6177 13676 6208
rect 13633 6171 13691 6177
rect 13633 6137 13645 6171
rect 13679 6137 13691 6171
rect 13633 6131 13691 6137
rect 11020 6072 11468 6100
rect 11020 6060 11026 6072
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 12066 6100 12072 6112
rect 11664 6072 12072 6100
rect 11664 6060 11670 6072
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13872 6072 14197 6100
rect 13872 6060 13878 6072
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14185 6063 14243 6069
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3234 5896 3240 5908
rect 2731 5868 3240 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3752 5868 3893 5896
rect 3752 5856 3758 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5626 5896 5632 5908
rect 5316 5868 5632 5896
rect 5316 5856 5322 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6638 5896 6644 5908
rect 6319 5868 6644 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6880 5868 7205 5896
rect 6880 5856 6886 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7340 5868 7481 5896
rect 7340 5856 7346 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 8113 5899 8171 5905
rect 7469 5859 7527 5865
rect 7576 5868 8064 5896
rect 1872 5828 1900 5856
rect 1872 5800 2774 5828
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1636 5732 1685 5760
rect 1636 5720 1642 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 2746 5760 2774 5800
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 3786 5828 3792 5840
rect 2924 5800 3792 5828
rect 2924 5788 2930 5800
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 7576 5828 7604 5868
rect 6840 5800 7604 5828
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 2746 5732 3065 5760
rect 1673 5723 1731 5729
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 4154 5760 4160 5772
rect 3283 5732 4160 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5534 5760 5540 5772
rect 5307 5732 5540 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 1486 5692 1492 5704
rect 1443 5664 1492 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1486 5652 1492 5664
rect 1544 5652 1550 5704
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2958 5692 2964 5704
rect 1903 5664 2964 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5692 5411 5695
rect 5399 5664 5580 5692
rect 5399 5661 5411 5664
rect 5353 5655 5411 5661
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 3620 5624 3648 5655
rect 1360 5596 3648 5624
rect 5016 5627 5074 5633
rect 1360 5584 1366 5596
rect 5016 5593 5028 5627
rect 5062 5624 5074 5627
rect 5442 5624 5448 5636
rect 5062 5596 5448 5624
rect 5062 5593 5074 5596
rect 5016 5587 5074 5593
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 5552 5624 5580 5664
rect 5626 5652 5632 5704
rect 5684 5652 5690 5704
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6840 5701 6868 5800
rect 7834 5788 7840 5840
rect 7892 5788 7898 5840
rect 8036 5828 8064 5868
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 9122 5896 9128 5908
rect 8159 5868 9128 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 10560 5868 11468 5896
rect 10560 5856 10566 5868
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 8036 5800 8217 5828
rect 8205 5797 8217 5800
rect 8251 5797 8263 5831
rect 9232 5828 9260 5856
rect 8205 5791 8263 5797
rect 8588 5800 9260 5828
rect 9677 5831 9735 5837
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 8294 5760 8300 5772
rect 6972 5732 7144 5760
rect 6972 5720 6978 5732
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7116 5701 7144 5732
rect 7668 5732 8300 5760
rect 7668 5701 7696 5732
rect 8294 5720 8300 5732
rect 8352 5760 8358 5772
rect 8588 5760 8616 5800
rect 9677 5797 9689 5831
rect 9723 5828 9735 5831
rect 10134 5828 10140 5840
rect 9723 5800 10140 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 10873 5831 10931 5837
rect 10873 5797 10885 5831
rect 10919 5797 10931 5831
rect 10873 5791 10931 5797
rect 8352 5732 8616 5760
rect 8352 5720 8358 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7607 5664 7665 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8588 5701 8616 5732
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 8711 5732 9229 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 10888 5760 10916 5791
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 10888 5732 11161 5760
rect 9217 5723 9275 5729
rect 11149 5729 11161 5732
rect 11195 5729 11207 5763
rect 11440 5760 11468 5868
rect 11514 5856 11520 5908
rect 11572 5856 11578 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 11756 5868 12725 5896
rect 11756 5856 11762 5868
rect 12713 5865 12725 5868
rect 12759 5865 12771 5899
rect 12713 5859 12771 5865
rect 13354 5856 13360 5908
rect 13412 5856 13418 5908
rect 14274 5856 14280 5908
rect 14332 5856 14338 5908
rect 12526 5788 12532 5840
rect 12584 5788 12590 5840
rect 13262 5760 13268 5772
rect 11440 5732 13268 5760
rect 11149 5723 11207 5729
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 14292 5760 14320 5856
rect 13372 5732 14320 5760
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7892 5664 7941 5692
rect 7892 5652 7898 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 7929 5655 7987 5661
rect 8036 5664 8401 5692
rect 6472 5624 6500 5652
rect 5552 5596 6500 5624
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2406 5556 2412 5568
rect 2363 5528 2412 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 3418 5516 3424 5568
rect 3476 5516 3482 5568
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 8036 5556 8064 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8573 5655 8631 5661
rect 8680 5664 9045 5692
rect 8680 5636 8708 5664
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 9858 5692 9864 5704
rect 9815 5664 9864 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 8662 5584 8668 5636
rect 8720 5584 8726 5636
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 9968 5624 9996 5655
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10796 5664 10977 5692
rect 10796 5624 10824 5664
rect 10965 5661 10977 5664
rect 11011 5692 11023 5695
rect 11606 5692 11612 5704
rect 11011 5664 11612 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 11882 5652 11888 5704
rect 11940 5652 11946 5704
rect 12066 5652 12072 5704
rect 12124 5652 12130 5704
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 9732 5596 9996 5624
rect 10244 5596 10824 5624
rect 9732 5584 9738 5596
rect 5583 5528 8064 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 9582 5556 9588 5568
rect 8536 5528 9588 5556
rect 8536 5516 8542 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10244 5556 10272 5596
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11698 5624 11704 5636
rect 10928 5596 11704 5624
rect 10928 5584 10934 5596
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12820 5624 12848 5652
rect 12492 5596 12848 5624
rect 12492 5584 12498 5596
rect 9824 5528 10272 5556
rect 9824 5516 9830 5528
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 10962 5556 10968 5568
rect 10376 5528 10968 5556
rect 10376 5516 10382 5528
rect 10962 5516 10968 5528
rect 11020 5556 11026 5568
rect 13372 5556 13400 5732
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13688 5664 13737 5692
rect 13688 5652 13694 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 11020 5528 13400 5556
rect 11020 5516 11026 5528
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 2406 5312 2412 5364
rect 2464 5312 2470 5364
rect 2958 5312 2964 5364
rect 3016 5312 3022 5364
rect 3605 5355 3663 5361
rect 3605 5321 3617 5355
rect 3651 5321 3663 5355
rect 4062 5352 4068 5364
rect 3605 5315 3663 5321
rect 3804 5324 4068 5352
rect 2866 5284 2872 5296
rect 2424 5256 2872 5284
rect 2424 5228 2452 5256
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 2976 5284 3004 5312
rect 3620 5284 3648 5315
rect 2976 5256 3648 5284
rect 1670 5176 1676 5228
rect 1728 5176 1734 5228
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3234 5216 3240 5228
rect 3099 5188 3240 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3418 5216 3424 5228
rect 3375 5188 3424 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 3804 5225 3832 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4798 5352 4804 5364
rect 4479 5324 4804 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5350 5312 5356 5364
rect 5408 5312 5414 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5500 5324 5764 5352
rect 5500 5312 5506 5324
rect 4982 5284 4988 5296
rect 4356 5256 4988 5284
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 4356 5225 4384 5256
rect 4982 5244 4988 5256
rect 5040 5244 5046 5296
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 5368 5284 5396 5312
rect 5736 5284 5764 5324
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 5905 5355 5963 5361
rect 5905 5352 5917 5355
rect 5868 5324 5917 5352
rect 5868 5312 5874 5324
rect 5905 5321 5917 5324
rect 5951 5321 5963 5355
rect 5905 5315 5963 5321
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 7708 5324 8125 5352
rect 7708 5312 7714 5324
rect 8113 5321 8125 5324
rect 8159 5352 8171 5355
rect 8202 5352 8208 5364
rect 8159 5324 8208 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9674 5352 9680 5364
rect 8803 5324 9680 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 5224 5256 5488 5284
rect 5736 5256 7880 5284
rect 5224 5244 5230 5256
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 5000 5216 5028 5244
rect 5460 5225 5488 5256
rect 5353 5219 5411 5225
rect 5000 5214 5304 5216
rect 5353 5214 5365 5219
rect 5000 5188 5365 5214
rect 5276 5186 5365 5188
rect 4341 5179 4399 5185
rect 5353 5185 5365 5186
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6454 5216 6460 5228
rect 6043 5188 6460 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6638 5216 6644 5228
rect 6595 5188 6644 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 6779 5188 7052 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 992 5120 1409 5148
rect 992 5108 998 5120
rect 1397 5117 1409 5120
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3528 5148 3556 5176
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 2915 5120 3556 5148
rect 4540 5120 4905 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 4065 5083 4123 5089
rect 2746 5052 3740 5080
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 2746 5012 2774 5052
rect 1820 4984 2774 5012
rect 1820 4972 1826 4984
rect 3418 4972 3424 5024
rect 3476 4972 3482 5024
rect 3712 5012 3740 5052
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4540 5080 4568 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5537 5151 5595 5157
rect 5123 5120 5304 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5276 5089 5304 5120
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5920 5148 5948 5176
rect 7024 5160 7052 5188
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 7248 5188 7788 5216
rect 7248 5176 7254 5188
rect 5583 5120 6684 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 4111 5052 4568 5080
rect 5261 5083 5319 5089
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 5261 5049 5273 5083
rect 5307 5080 5319 5083
rect 5307 5052 5672 5080
rect 5307 5049 5319 5052
rect 5261 5043 5319 5049
rect 5644 5024 5672 5052
rect 6656 5024 6684 5120
rect 6914 5108 6920 5160
rect 6972 5108 6978 5160
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 7116 5120 7481 5148
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 3712 4984 4169 5012
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 4157 4975 4215 4981
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4890 5012 4896 5024
rect 4672 4984 4896 5012
rect 4672 4972 4678 4984
rect 4890 4972 4896 4984
rect 4948 5012 4954 5024
rect 5350 5012 5356 5024
rect 4948 4984 5356 5012
rect 4948 4972 4954 4984
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6638 4972 6644 5024
rect 6696 4972 6702 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7116 5021 7144 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 7760 5080 7788 5188
rect 7852 5148 7880 5256
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 8496 5216 8524 5315
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 11057 5355 11115 5361
rect 11057 5352 11069 5355
rect 10744 5324 11069 5352
rect 10744 5312 10750 5324
rect 11057 5321 11069 5324
rect 11103 5321 11115 5355
rect 11057 5315 11115 5321
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 12066 5352 12072 5364
rect 11747 5324 12072 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12584 5324 14044 5352
rect 12584 5312 12590 5324
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 12345 5287 12403 5293
rect 12345 5284 12357 5287
rect 8996 5256 12357 5284
rect 8996 5244 9002 5256
rect 12345 5253 12357 5256
rect 12391 5253 12403 5287
rect 12345 5247 12403 5253
rect 12437 5287 12495 5293
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 12483 5256 13277 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 13265 5253 13277 5256
rect 13311 5284 13323 5287
rect 13357 5287 13415 5293
rect 13357 5284 13369 5287
rect 13311 5256 13369 5284
rect 13311 5253 13323 5256
rect 13265 5247 13323 5253
rect 13357 5253 13369 5256
rect 13403 5253 13415 5287
rect 13357 5247 13415 5253
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8496 5188 8585 5216
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 9364 5188 9597 5216
rect 9364 5176 9370 5188
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 9692 5188 9996 5216
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 7852 5120 8861 5148
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9692 5148 9720 5188
rect 9447 5120 9720 5148
rect 9769 5151 9827 5157
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 9769 5117 9781 5151
rect 9815 5148 9827 5151
rect 9858 5148 9864 5160
rect 9815 5120 9864 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 9416 5080 9444 5111
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 9968 5148 9996 5188
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10192 5188 10333 5216
rect 10192 5176 10198 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10428 5188 10640 5216
rect 10428 5148 10456 5188
rect 9968 5120 10456 5148
rect 10502 5108 10508 5160
rect 10560 5108 10566 5160
rect 10612 5148 10640 5188
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 11514 5176 11520 5228
rect 11572 5176 11578 5228
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5216 13875 5219
rect 13906 5216 13912 5228
rect 13863 5188 13912 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14016 5225 14044 5324
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14826 5216 14832 5228
rect 14415 5188 14832 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 11606 5148 11612 5160
rect 10612 5120 11612 5148
rect 11606 5108 11612 5120
rect 11664 5108 11670 5160
rect 11974 5108 11980 5160
rect 12032 5108 12038 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 13354 5148 13360 5160
rect 12851 5120 13360 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 7760 5052 9444 5080
rect 9582 5040 9588 5092
rect 9640 5080 9646 5092
rect 12710 5080 12716 5092
rect 9640 5040 9674 5080
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6788 4984 7113 5012
rect 6788 4972 6794 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 9646 5012 9674 5040
rect 9876 5052 12716 5080
rect 9876 5012 9904 5052
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 14182 5040 14188 5092
rect 14240 5040 14246 5092
rect 9646 4984 9904 5012
rect 7101 4975 7159 4981
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10689 5015 10747 5021
rect 10689 5012 10701 5015
rect 10192 4984 10701 5012
rect 10192 4972 10198 4984
rect 10689 4981 10701 4984
rect 10735 4981 10747 5015
rect 10689 4975 10747 4981
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 12066 5012 12072 5024
rect 11296 4984 12072 5012
rect 11296 4972 11302 4984
rect 12066 4972 12072 4984
rect 12124 5012 12130 5024
rect 12434 5012 12440 5024
rect 12124 4984 12440 5012
rect 12124 4972 12130 4984
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2222 4808 2228 4820
rect 1995 4780 2228 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 3568 4780 5549 4808
rect 3568 4768 3574 4780
rect 5537 4777 5549 4780
rect 5583 4777 5595 4811
rect 5537 4771 5595 4777
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 6086 4808 6092 4820
rect 5776 4780 6092 4808
rect 5776 4768 5782 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 6825 4811 6883 4817
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 6914 4808 6920 4820
rect 6871 4780 6920 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7469 4811 7527 4817
rect 7469 4777 7481 4811
rect 7515 4808 7527 4811
rect 7650 4808 7656 4820
rect 7515 4780 7656 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4808 8079 4811
rect 8478 4808 8484 4820
rect 8067 4780 8484 4808
rect 8067 4777 8079 4780
rect 8021 4771 8079 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 8938 4808 8944 4820
rect 8803 4780 8944 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9030 4768 9036 4820
rect 9088 4768 9094 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9766 4808 9772 4820
rect 9723 4780 9772 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10502 4808 10508 4820
rect 10091 4780 10508 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11514 4808 11520 4820
rect 11379 4780 11520 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 11664 4780 13400 4808
rect 11664 4768 11670 4780
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 3234 4740 3240 4752
rect 2823 4712 3240 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 3970 4740 3976 4752
rect 3476 4712 3976 4740
rect 3476 4700 3482 4712
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 4985 4743 5043 4749
rect 4985 4740 4997 4743
rect 4764 4712 4997 4740
rect 4764 4700 4770 4712
rect 4985 4709 4997 4712
rect 5031 4709 5043 4743
rect 4985 4703 5043 4709
rect 5261 4743 5319 4749
rect 5261 4709 5273 4743
rect 5307 4709 5319 4743
rect 5261 4703 5319 4709
rect 2130 4632 2136 4684
rect 2188 4632 2194 4684
rect 2314 4632 2320 4684
rect 2372 4632 2378 4684
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 3142 4672 3148 4684
rect 3099 4644 3148 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 5276 4672 5304 4703
rect 5350 4700 5356 4752
rect 5408 4700 5414 4752
rect 5813 4743 5871 4749
rect 5813 4709 5825 4743
rect 5859 4709 5871 4743
rect 5813 4703 5871 4709
rect 7101 4743 7159 4749
rect 7101 4709 7113 4743
rect 7147 4709 7159 4743
rect 7101 4703 7159 4709
rect 3620 4644 5304 4672
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1636 4576 1777 4604
rect 1636 4564 1642 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 1765 4567 1823 4573
rect 2746 4576 2881 4604
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 2746 4536 2774 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 1719 4508 2774 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 3620 4468 3648 4644
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 3752 4576 3893 4604
rect 3752 4564 3758 4576
rect 3881 4573 3893 4576
rect 3927 4604 3939 4607
rect 4614 4604 4620 4616
rect 3927 4576 4620 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4614 4564 4620 4576
rect 4672 4604 4678 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4672 4576 4721 4604
rect 4672 4564 4678 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 4948 4576 5181 4604
rect 4948 4564 4954 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5368 4604 5396 4700
rect 5828 4672 5856 4703
rect 5736 4644 5856 4672
rect 5736 4613 5764 4644
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5960 4644 6101 4672
rect 5960 4632 5966 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6454 4672 6460 4684
rect 6319 4644 6460 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6822 4632 6828 4684
rect 6880 4632 6886 4684
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5368 4576 5457 4604
rect 5169 4567 5227 4573
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5721 4567 5779 4573
rect 5828 4576 6009 4604
rect 4798 4496 4804 4548
rect 4856 4496 4862 4548
rect 5460 4536 5488 4567
rect 5828 4536 5856 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 5460 4508 5856 4536
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6840 4536 6868 4632
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7116 4604 7144 4703
rect 8294 4700 8300 4752
rect 8352 4700 8358 4752
rect 10873 4743 10931 4749
rect 10873 4740 10885 4743
rect 9140 4712 10885 4740
rect 8312 4672 8340 4700
rect 8312 4644 8432 4672
rect 7055 4576 7144 4604
rect 7285 4607 7343 4613
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 7300 4536 7328 4567
rect 5960 4508 7328 4536
rect 7668 4536 7696 4567
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8404 4613 8432 4644
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8478 4604 8484 4616
rect 8435 4576 8484 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9140 4604 9168 4712
rect 10873 4709 10885 4712
rect 10919 4709 10931 4743
rect 13372 4740 13400 4780
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13596 4780 14197 4808
rect 13596 4768 13602 4780
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 14185 4771 14243 4777
rect 13817 4743 13875 4749
rect 13817 4740 13829 4743
rect 13372 4712 13829 4740
rect 10873 4703 10931 4709
rect 13817 4709 13829 4712
rect 13863 4709 13875 4743
rect 13817 4703 13875 4709
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 9766 4672 9772 4684
rect 9539 4644 9772 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 12216 4644 12480 4672
rect 12216 4632 12222 4644
rect 8619 4576 9168 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9582 4564 9588 4616
rect 9640 4564 9646 4616
rect 9869 4603 9927 4609
rect 9869 4569 9881 4603
rect 9915 4600 9927 4603
rect 9915 4572 9996 4600
rect 9915 4569 9927 4572
rect 9869 4563 9927 4569
rect 9968 4536 9996 4572
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 10376 4576 10609 4604
rect 10376 4564 10382 4576
rect 10597 4573 10609 4576
rect 10643 4573 10655 4607
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10597 4567 10655 4573
rect 10980 4576 11069 4604
rect 10980 4536 11008 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4604 11207 4607
rect 11256 4604 11284 4632
rect 11698 4604 11704 4616
rect 11195 4576 11284 4604
rect 11348 4576 11704 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 11348 4536 11376 4576
rect 11698 4564 11704 4576
rect 11756 4604 11762 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11756 4576 11805 4604
rect 11756 4564 11762 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 12452 4613 12480 4644
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 12483 4576 12940 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 7668 4508 8248 4536
rect 9968 4508 10456 4536
rect 5960 4496 5966 4508
rect 1912 4440 3648 4468
rect 1912 4428 1918 4440
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 8220 4477 8248 4508
rect 4433 4471 4491 4477
rect 4433 4468 4445 4471
rect 4304 4440 4445 4468
rect 4304 4428 4310 4440
rect 4433 4437 4445 4440
rect 4479 4437 4491 4471
rect 4433 4431 4491 4437
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10428 4477 10456 4508
rect 10980 4508 11376 4536
rect 11609 4539 11667 4545
rect 10980 4480 11008 4508
rect 11609 4505 11621 4539
rect 11655 4536 11667 4539
rect 11900 4536 11928 4564
rect 11655 4508 11928 4536
rect 12345 4539 12403 4545
rect 11655 4505 11667 4508
rect 11609 4499 11667 4505
rect 12345 4505 12357 4539
rect 12391 4536 12403 4539
rect 12682 4539 12740 4545
rect 12682 4536 12694 4539
rect 12391 4508 12694 4536
rect 12391 4505 12403 4508
rect 12345 4499 12403 4505
rect 12682 4505 12694 4508
rect 12728 4505 12740 4539
rect 12682 4499 12740 4505
rect 12912 4480 12940 4576
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 10229 4471 10287 4477
rect 10229 4468 10241 4471
rect 10008 4440 10241 4468
rect 10008 4428 10014 4440
rect 10229 4437 10241 4440
rect 10275 4437 10287 4471
rect 10229 4431 10287 4437
rect 10413 4471 10471 4477
rect 10413 4437 10425 4471
rect 10459 4437 10471 4471
rect 10413 4431 10471 4437
rect 10962 4428 10968 4480
rect 11020 4428 11026 4480
rect 12894 4428 12900 4480
rect 12952 4428 12958 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 3878 4224 3884 4276
rect 3936 4264 3942 4276
rect 3973 4267 4031 4273
rect 3973 4264 3985 4267
rect 3936 4236 3985 4264
rect 3936 4224 3942 4236
rect 3973 4233 3985 4236
rect 4019 4233 4031 4267
rect 3973 4227 4031 4233
rect 5905 4267 5963 4273
rect 5905 4233 5917 4267
rect 5951 4233 5963 4267
rect 5905 4227 5963 4233
rect 3418 4196 3424 4208
rect 2700 4168 3424 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1544 4100 1685 4128
rect 1544 4088 1550 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2700 4137 2728 4168
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 4706 4196 4712 4208
rect 4571 4168 4712 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 4798 4156 4804 4208
rect 4856 4196 4862 4208
rect 4856 4168 5672 4196
rect 4856 4156 4862 4168
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 2188 4100 2513 4128
rect 2188 4088 2194 4100
rect 2501 4097 2513 4100
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 3142 4128 3148 4140
rect 2685 4091 2743 4097
rect 2884 4100 3148 4128
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 992 4032 1409 4060
rect 992 4020 998 4032
rect 1397 4029 1409 4032
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 2130 3952 2136 4004
rect 2188 3992 2194 4004
rect 2884 3992 2912 4100
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5442 4128 5448 4140
rect 5123 4100 5448 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5644 4137 5672 4168
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5920 4128 5948 4227
rect 6086 4224 6092 4276
rect 6144 4224 6150 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7193 4267 7251 4273
rect 7193 4264 7205 4267
rect 7064 4236 7205 4264
rect 7064 4224 7070 4236
rect 7193 4233 7205 4236
rect 7239 4233 7251 4267
rect 7193 4227 7251 4233
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 12250 4264 12256 4276
rect 9272 4236 12256 4264
rect 9272 4224 9278 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12989 4267 13047 4273
rect 12989 4233 13001 4267
rect 13035 4233 13047 4267
rect 12989 4227 13047 4233
rect 6104 4137 6132 4224
rect 6638 4156 6644 4208
rect 6696 4196 6702 4208
rect 6696 4168 6960 4196
rect 6696 4156 6702 4168
rect 5629 4091 5687 4097
rect 5736 4100 5948 4128
rect 6089 4131 6147 4137
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3510 4060 3516 4072
rect 3467 4032 3516 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 3620 4032 4445 4060
rect 3620 4001 3648 4032
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5736 4060 5764 4100
rect 6089 4097 6101 4131
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6730 4088 6736 4140
rect 6788 4088 6794 4140
rect 5316 4032 5764 4060
rect 5813 4063 5871 4069
rect 5316 4020 5322 4032
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5994 4060 6000 4072
rect 5859 4032 6000 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6932 4060 6960 4168
rect 7484 4168 7696 4196
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7484 4128 7512 4168
rect 7331 4100 7512 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7668 4128 7696 4168
rect 8496 4168 8708 4196
rect 8496 4128 8524 4168
rect 7668 4100 8524 4128
rect 8570 4088 8576 4140
rect 8628 4088 8634 4140
rect 8680 4128 8708 4168
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 10689 4199 10747 4205
rect 9640 4168 9996 4196
rect 9640 4156 9646 4168
rect 9858 4128 9864 4140
rect 8680 4100 9864 4128
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9968 4072 9996 4168
rect 10689 4165 10701 4199
rect 10735 4196 10747 4199
rect 11057 4199 11115 4205
rect 11057 4196 11069 4199
rect 10735 4168 11069 4196
rect 10735 4165 10747 4168
rect 10689 4159 10747 4165
rect 11057 4165 11069 4168
rect 11103 4165 11115 4199
rect 11057 4159 11115 4165
rect 11698 4156 11704 4208
rect 11756 4196 11762 4208
rect 13004 4196 13032 4227
rect 11756 4168 13032 4196
rect 14016 4168 14228 4196
rect 11756 4156 11762 4168
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10100 4100 10149 4128
rect 10100 4088 10106 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 6932 4032 7665 4060
rect 6825 4023 6883 4029
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8260 4032 8677 4060
rect 8260 4020 8266 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9674 4060 9680 4072
rect 8895 4032 9680 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10318 4060 10324 4072
rect 10008 4032 10324 4060
rect 10008 4020 10014 4032
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 2188 3964 2912 3992
rect 3145 3995 3203 4001
rect 2188 3952 2194 3964
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3605 3995 3663 4001
rect 3605 3992 3617 3995
rect 3191 3964 3617 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 3605 3961 3617 3964
rect 3651 3961 3663 3995
rect 3605 3955 3663 3961
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 7248 3964 8401 3992
rect 7248 3952 7254 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 9306 3952 9312 4004
rect 9364 3992 9370 4004
rect 10796 3992 10824 4023
rect 9364 3964 10824 3992
rect 9364 3952 9370 3964
rect 5166 3884 5172 3936
rect 5224 3884 5230 3936
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 7098 3924 7104 3936
rect 5776 3896 7104 3924
rect 5776 3884 5782 3896
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7374 3884 7380 3936
rect 7432 3884 7438 3936
rect 8110 3884 8116 3936
rect 8168 3884 8174 3936
rect 9398 3884 9404 3936
rect 9456 3884 9462 3936
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10980 3924 11008 4091
rect 12618 4088 12624 4140
rect 12676 4137 12682 4140
rect 12676 4091 12688 4137
rect 12676 4088 12682 4091
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 14016 4128 14044 4168
rect 12952 4100 14044 4128
rect 12952 4088 12958 4100
rect 14090 4088 14096 4140
rect 14148 4137 14154 4140
rect 14148 4091 14160 4137
rect 14200 4128 14228 4168
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 14200 4100 14381 4128
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14148 4088 14154 4091
rect 10468 3896 11008 3924
rect 10468 3884 10474 3896
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11514 3924 11520 3936
rect 11204 3896 11520 3924
rect 11204 3884 11210 3896
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 2958 3720 2964 3732
rect 1903 3692 2964 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 6638 3720 6644 3732
rect 3200 3692 6644 3720
rect 3200 3680 3206 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7892 3692 7941 3720
rect 7892 3680 7898 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8570 3680 8576 3732
rect 8628 3680 8634 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 9306 3720 9312 3732
rect 8803 3692 9312 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9916 3692 12434 3720
rect 9916 3680 9922 3692
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 2038 3652 2044 3664
rect 1627 3624 2044 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 2038 3612 2044 3624
rect 2096 3612 2102 3664
rect 2130 3612 2136 3664
rect 2188 3612 2194 3664
rect 3605 3655 3663 3661
rect 3605 3621 3617 3655
rect 3651 3652 3663 3655
rect 3694 3652 3700 3664
rect 3651 3624 3700 3652
rect 3651 3621 3663 3624
rect 3605 3615 3663 3621
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 3970 3612 3976 3664
rect 4028 3612 4034 3664
rect 4430 3612 4436 3664
rect 4488 3612 4494 3664
rect 5813 3655 5871 3661
rect 5813 3621 5825 3655
rect 5859 3652 5871 3655
rect 5902 3652 5908 3664
rect 5859 3624 5908 3652
rect 5859 3621 5871 3624
rect 5813 3615 5871 3621
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 8588 3652 8616 3680
rect 7708 3624 8616 3652
rect 7708 3612 7714 3624
rect 4154 3584 4160 3596
rect 4080 3556 4160 3584
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1854 3516 1860 3528
rect 1719 3488 1860 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1412 3448 1440 3479
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2271 3488 2774 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 1964 3448 1992 3479
rect 2498 3457 2504 3460
rect 1412 3420 1900 3448
rect 1964 3420 2360 3448
rect 1872 3380 1900 3420
rect 2130 3380 2136 3392
rect 1872 3352 2136 3380
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 2332 3380 2360 3420
rect 2492 3411 2504 3457
rect 2498 3408 2504 3411
rect 2556 3408 2562 3460
rect 2746 3448 2774 3488
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4080 3525 4108 3556
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 4448 3584 4476 3612
rect 4212 3556 4476 3584
rect 4212 3544 4218 3556
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 5592 3556 6285 3584
rect 5592 3544 5598 3556
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 5552 3516 5580 3544
rect 4479 3488 5580 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 4448 3448 4476 3479
rect 5994 3476 6000 3528
rect 6052 3476 6058 3528
rect 8036 3525 8064 3624
rect 8846 3612 8852 3664
rect 8904 3612 8910 3664
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 10468 3624 10517 3652
rect 10468 3612 10474 3624
rect 10505 3621 10517 3624
rect 10551 3621 10563 3655
rect 10505 3615 10563 3621
rect 12066 3612 12072 3664
rect 12124 3612 12130 3664
rect 12406 3652 12434 3692
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12676 3692 12909 3720
rect 12676 3680 12682 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14090 3720 14096 3732
rect 13955 3692 14096 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14366 3680 14372 3732
rect 14424 3680 14430 3732
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12406 3624 13001 3652
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 14274 3612 14280 3664
rect 14332 3612 14338 3664
rect 8110 3544 8116 3596
rect 8168 3544 8174 3596
rect 8864 3584 8892 3612
rect 12802 3584 12808 3596
rect 8220 3556 8892 3584
rect 11716 3556 12808 3584
rect 8021 3519 8079 3525
rect 6104 3488 6684 3516
rect 4706 3457 4712 3460
rect 2746 3420 4476 3448
rect 4700 3411 4712 3457
rect 4706 3408 4712 3411
rect 4764 3408 4770 3460
rect 4890 3408 4896 3460
rect 4948 3408 4954 3460
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 6104 3448 6132 3488
rect 5040 3420 6132 3448
rect 5040 3408 5046 3420
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 6518 3451 6576 3457
rect 6518 3448 6530 3451
rect 6420 3420 6530 3448
rect 6420 3408 6426 3420
rect 6518 3417 6530 3420
rect 6564 3417 6576 3451
rect 6656 3448 6684 3488
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8220 3448 8248 3556
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 6656 3420 8248 3448
rect 6518 3411 6576 3417
rect 3510 3380 3516 3392
rect 2332 3352 3516 3380
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 4908 3380 4936 3408
rect 4295 3352 4936 3380
rect 6089 3383 6147 3389
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 6638 3380 6644 3392
rect 6135 3352 6644 3380
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 8312 3380 8340 3479
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 9180 3488 10701 3516
rect 9180 3476 9186 3488
rect 10689 3485 10701 3488
rect 10735 3516 10747 3519
rect 11716 3516 11744 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 14292 3584 14320 3612
rect 13188 3556 14320 3584
rect 10735 3488 11744 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 13188 3525 13216 3556
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12124 3488 12265 3516
rect 12124 3476 12130 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14182 3516 14188 3528
rect 13403 3488 14188 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 9398 3457 9404 3460
rect 9392 3448 9404 3457
rect 9359 3420 9404 3448
rect 9392 3411 9404 3420
rect 9398 3408 9404 3411
rect 9456 3408 9462 3460
rect 10956 3451 11014 3457
rect 10428 3420 10916 3448
rect 10428 3380 10456 3420
rect 8312 3352 10456 3380
rect 10888 3380 10916 3420
rect 10956 3417 10968 3451
rect 11002 3448 11014 3451
rect 11146 3448 11152 3460
rect 11002 3420 11152 3448
rect 11002 3417 11014 3420
rect 10956 3411 11014 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 13372 3448 13400 3479
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14550 3516 14556 3528
rect 14323 3488 14556 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 11572 3420 13400 3448
rect 11572 3408 11578 3420
rect 11606 3380 11612 3392
rect 10888 3352 11612 3380
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 14182 3380 14188 3392
rect 11940 3352 14188 3380
rect 11940 3340 11946 3352
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 2682 3136 2688 3188
rect 2740 3136 2746 3188
rect 2774 3136 2780 3188
rect 2832 3136 2838 3188
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 2976 3148 3249 3176
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2700 3040 2728 3136
rect 2455 3012 2728 3040
rect 2869 3043 2927 3049
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2976 3040 3004 3148
rect 3237 3145 3249 3148
rect 3283 3176 3295 3179
rect 4154 3176 4160 3188
rect 3283 3148 4160 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5534 3176 5540 3188
rect 4632 3148 5540 3176
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 3099 3080 4200 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2976 3012 3157 3040
rect 2869 3003 2927 3009
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 4062 3040 4068 3052
rect 3145 3003 3203 3009
rect 3252 3012 4068 3040
rect 1394 2932 1400 2984
rect 1452 2932 1458 2984
rect 2884 2972 2912 3003
rect 3252 2972 3280 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4172 3040 4200 3080
rect 4246 3068 4252 3120
rect 4304 3108 4310 3120
rect 4350 3111 4408 3117
rect 4350 3108 4362 3111
rect 4304 3080 4362 3108
rect 4304 3068 4310 3080
rect 4350 3077 4362 3080
rect 4396 3077 4408 3111
rect 4350 3071 4408 3077
rect 4632 3049 4660 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 7190 3136 7196 3188
rect 7248 3136 7254 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 10594 3176 10600 3188
rect 9907 3148 10600 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11204 3148 11529 3176
rect 11204 3136 11210 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 11664 3148 12940 3176
rect 11664 3136 11670 3148
rect 5261 3111 5319 3117
rect 5261 3108 5273 3111
rect 4724 3080 5273 3108
rect 4617 3043 4675 3049
rect 4172 3012 4568 3040
rect 2884 2944 3280 2972
rect 4540 2972 4568 3012
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4724 2972 4752 3080
rect 5261 3077 5273 3080
rect 5307 3077 5319 3111
rect 5261 3071 5319 3077
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 7006 3108 7012 3120
rect 5408 3080 7012 3108
rect 5408 3068 5414 3080
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4540 2944 4752 2972
rect 2746 2876 3188 2904
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2746 2836 2774 2876
rect 3160 2848 3188 2876
rect 2639 2808 2774 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 3142 2796 3148 2848
rect 3200 2796 3206 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4816 2836 4844 3003
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 7208 3040 7236 3136
rect 7392 3049 7420 3136
rect 7561 3111 7619 3117
rect 7561 3077 7573 3111
rect 7607 3108 7619 3111
rect 8754 3108 8760 3120
rect 7607 3080 8760 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 9272 3080 9413 3108
rect 9272 3068 9278 3080
rect 9401 3077 9413 3080
rect 9447 3077 9459 3111
rect 10612 3108 10640 3136
rect 12802 3108 12808 3120
rect 10612 3080 11100 3108
rect 9401 3071 9459 3077
rect 6043 3012 7236 3040
rect 7377 3043 7435 3049
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 5442 2932 5448 2984
rect 5500 2932 5506 2984
rect 5920 2972 5948 3000
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 5920 2944 6929 2972
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 5460 2904 5488 2932
rect 7484 2904 7512 3003
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8858 3043 8916 3049
rect 8858 3040 8870 3043
rect 8536 3012 8870 3040
rect 8536 3000 8542 3012
rect 8858 3009 8870 3012
rect 8904 3009 8916 3043
rect 8858 3003 8916 3009
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 10962 3000 10968 3052
rect 11020 3049 11026 3052
rect 11020 3003 11032 3049
rect 11072 3040 11100 3080
rect 11256 3080 12808 3108
rect 11256 3049 11284 3080
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 12912 3108 12940 3148
rect 13173 3111 13231 3117
rect 12912 3080 13124 3108
rect 11241 3043 11299 3049
rect 11072 3012 11192 3040
rect 11020 3000 11026 3003
rect 11164 2972 11192 3012
rect 11241 3009 11253 3043
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11164 2944 12081 2972
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 13004 2972 13032 3003
rect 12216 2944 13032 2972
rect 12216 2932 12222 2944
rect 9950 2904 9956 2916
rect 5460 2876 7512 2904
rect 9324 2876 9956 2904
rect 4304 2808 4844 2836
rect 6181 2839 6239 2845
rect 4304 2796 4310 2808
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6914 2836 6920 2848
rect 6227 2808 6920 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 7248 2808 7297 2836
rect 7248 2796 7254 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 8386 2836 8392 2848
rect 7791 2808 8392 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 8386 2796 8392 2808
rect 8444 2836 8450 2848
rect 9324 2836 9352 2876
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13096 2904 13124 3080
rect 13173 3077 13185 3111
rect 13219 3108 13231 3111
rect 13262 3108 13268 3120
rect 13219 3080 13268 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 14182 3000 14188 3052
rect 14240 3000 14246 3052
rect 14458 3000 14464 3052
rect 14516 3000 14522 3052
rect 12851 2876 13124 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 8444 2808 9352 2836
rect 8444 2796 8450 2808
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9456 2808 9505 2836
rect 9456 2796 9462 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 10928 2808 12449 2836
rect 10928 2796 10934 2808
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 14550 2836 14556 2848
rect 13495 2808 14556 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 4706 2592 4712 2644
rect 4764 2592 4770 2644
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8202 2632 8208 2644
rect 7791 2604 8208 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2632 8815 2635
rect 8803 2604 10916 2632
rect 8803 2601 8815 2604
rect 8757 2595 8815 2601
rect 2038 2524 2044 2576
rect 2096 2524 2102 2576
rect 2406 2524 2412 2576
rect 2464 2524 2470 2576
rect 4522 2564 4528 2576
rect 3160 2536 4528 2564
rect 3160 2505 3188 2536
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 4617 2567 4675 2573
rect 4617 2533 4629 2567
rect 4663 2564 4675 2567
rect 5184 2564 5212 2592
rect 4663 2536 5212 2564
rect 5813 2567 5871 2573
rect 4663 2533 4675 2536
rect 4617 2527 4675 2533
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5859 2536 6377 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 10042 2564 10048 2576
rect 9631 2536 10048 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2465 3203 2499
rect 3145 2459 3203 2465
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 3973 2499 4031 2505
rect 3292 2468 3556 2496
rect 3292 2456 3298 2468
rect 566 2388 572 2440
rect 624 2428 630 2440
rect 3421 2431 3479 2437
rect 624 2400 1900 2428
rect 624 2388 630 2400
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 1360 2332 1501 2360
rect 1360 2320 1366 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 1670 2320 1676 2372
rect 1728 2320 1734 2372
rect 1872 2369 1900 2400
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3528 2428 3556 2468
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 5828 2496 5856 2527
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 10226 2524 10232 2576
rect 10284 2564 10290 2576
rect 10888 2564 10916 2604
rect 10962 2592 10968 2644
rect 11020 2592 11026 2644
rect 12158 2592 12164 2644
rect 12216 2592 12222 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13817 2635 13875 2641
rect 13817 2632 13829 2635
rect 13412 2604 13829 2632
rect 13412 2592 13418 2604
rect 13817 2601 13829 2604
rect 13863 2601 13875 2635
rect 13817 2595 13875 2601
rect 14090 2592 14096 2644
rect 14148 2592 14154 2644
rect 12176 2564 12204 2592
rect 10284 2536 10824 2564
rect 10888 2536 12204 2564
rect 10284 2524 10290 2536
rect 4019 2468 5856 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6696 2468 6837 2496
rect 6696 2456 6702 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6972 2468 7297 2496
rect 6972 2456 6978 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7708 2468 7849 2496
rect 7708 2456 7714 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 10134 2456 10140 2508
rect 10192 2456 10198 2508
rect 10410 2456 10416 2508
rect 10468 2456 10474 2508
rect 10796 2496 10824 2536
rect 14108 2496 14136 2592
rect 10796 2468 12204 2496
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 3528 2400 4169 2428
rect 3421 2391 3479 2397
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 1857 2363 1915 2369
rect 1857 2329 1869 2363
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2222 2320 2228 2372
rect 2280 2320 2286 2372
rect 3436 2360 3464 2391
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4856 2400 5273 2428
rect 4856 2388 4862 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6454 2428 6460 2440
rect 6227 2400 6460 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 4982 2360 4988 2372
rect 3436 2332 4988 2360
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 6012 2292 6040 2391
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2428 7159 2431
rect 7190 2428 7196 2440
rect 7147 2400 7196 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 7024 2360 7052 2391
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8444 2400 8585 2428
rect 8444 2388 8450 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8812 2400 9045 2428
rect 8812 2388 8818 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 12176 2437 12204 2468
rect 13924 2468 14136 2496
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11112 2400 11345 2428
rect 11112 2388 11118 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13924 2437 13952 2468
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12492 2400 13277 2428
rect 12492 2388 12498 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 7282 2360 7288 2372
rect 7024 2332 7288 2360
rect 7282 2320 7288 2332
rect 7340 2360 7346 2372
rect 8220 2360 8248 2388
rect 7340 2332 8248 2360
rect 10045 2363 10103 2369
rect 7340 2320 7346 2332
rect 10045 2329 10057 2363
rect 10091 2329 10103 2363
rect 10045 2323 10103 2329
rect 3200 2264 6040 2292
rect 3200 2252 3206 2264
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8904 2264 9137 2292
rect 8904 2252 8910 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 10060 2292 10088 2323
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 10468 2332 11284 2360
rect 10468 2320 10474 2332
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 10060 2264 11161 2292
rect 9125 2255 9183 2261
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11256 2292 11284 2332
rect 11606 2320 11612 2372
rect 11664 2320 11670 2372
rect 12710 2320 12716 2372
rect 12768 2320 12774 2372
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11256 2264 11713 2292
rect 11149 2255 11207 2261
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 11940 2264 12265 2292
rect 11940 2252 11946 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12253 2255 12311 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12400 2264 12817 2292
rect 12400 2252 12406 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13136 2264 13369 2292
rect 13136 2252 13142 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 14182 2252 14188 2304
rect 14240 2252 14246 2304
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 6178 2088 6184 2100
rect 2372 2060 6184 2088
rect 2372 2048 2378 2060
rect 6178 2048 6184 2060
rect 6236 2048 6242 2100
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 14182 2088 14188 2100
rect 8260 2060 14188 2088
rect 8260 2048 8266 2060
rect 14182 2048 14188 2060
rect 14240 2048 14246 2100
rect 2774 1980 2780 2032
rect 2832 2020 2838 2032
rect 5258 2020 5264 2032
rect 2832 1992 5264 2020
rect 2832 1980 2838 1992
rect 5258 1980 5264 1992
rect 5316 1980 5322 2032
<< via1 >>
rect 9864 22108 9916 22160
rect 11428 22108 11480 22160
rect 3792 21972 3844 22024
rect 5264 21972 5316 22024
rect 3976 21904 4028 21956
rect 9220 21904 9272 21956
rect 3056 21836 3108 21888
rect 8576 21836 8628 21888
rect 4376 21734 4428 21786
rect 4440 21734 4492 21786
rect 4504 21734 4556 21786
rect 4568 21734 4620 21786
rect 4632 21734 4684 21786
rect 7803 21734 7855 21786
rect 7867 21734 7919 21786
rect 7931 21734 7983 21786
rect 7995 21734 8047 21786
rect 8059 21734 8111 21786
rect 11230 21734 11282 21786
rect 11294 21734 11346 21786
rect 11358 21734 11410 21786
rect 11422 21734 11474 21786
rect 11486 21734 11538 21786
rect 14657 21734 14709 21786
rect 14721 21734 14773 21786
rect 14785 21734 14837 21786
rect 14849 21734 14901 21786
rect 14913 21734 14965 21786
rect 2780 21632 2832 21684
rect 3056 21675 3108 21684
rect 3056 21641 3065 21675
rect 3065 21641 3099 21675
rect 3099 21641 3108 21675
rect 3056 21632 3108 21641
rect 2044 21564 2096 21616
rect 1400 21496 1452 21548
rect 940 21428 992 21480
rect 2136 21539 2188 21548
rect 2136 21505 2145 21539
rect 2145 21505 2179 21539
rect 2179 21505 2188 21539
rect 2136 21496 2188 21505
rect 4068 21564 4120 21616
rect 5540 21632 5592 21684
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 3792 21539 3844 21548
rect 3792 21505 3801 21539
rect 3801 21505 3835 21539
rect 3835 21505 3844 21539
rect 3792 21496 3844 21505
rect 4252 21471 4304 21480
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 4804 21496 4856 21548
rect 5264 21564 5316 21616
rect 5172 21539 5224 21548
rect 5172 21505 5181 21539
rect 5181 21505 5215 21539
rect 5215 21505 5224 21539
rect 5172 21496 5224 21505
rect 5816 21632 5868 21684
rect 6828 21564 6880 21616
rect 6920 21564 6972 21616
rect 6092 21428 6144 21480
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 3424 21292 3476 21344
rect 3976 21335 4028 21344
rect 3976 21301 3985 21335
rect 3985 21301 4019 21335
rect 4019 21301 4028 21335
rect 3976 21292 4028 21301
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 7656 21632 7708 21684
rect 8484 21675 8536 21684
rect 8484 21641 8493 21675
rect 8493 21641 8527 21675
rect 8527 21641 8536 21675
rect 8484 21632 8536 21641
rect 8576 21632 8628 21684
rect 9036 21632 9088 21684
rect 9772 21632 9824 21684
rect 10784 21675 10836 21684
rect 10784 21641 10793 21675
rect 10793 21641 10827 21675
rect 10827 21641 10836 21675
rect 10784 21632 10836 21641
rect 11152 21632 11204 21684
rect 13360 21632 13412 21684
rect 7288 21496 7340 21548
rect 8484 21496 8536 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 10140 21428 10192 21480
rect 14464 21496 14516 21548
rect 7380 21360 7432 21412
rect 7932 21360 7984 21412
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 12808 21428 12860 21480
rect 4712 21292 4764 21344
rect 4988 21292 5040 21344
rect 5356 21335 5408 21344
rect 5356 21301 5365 21335
rect 5365 21301 5399 21335
rect 5399 21301 5408 21335
rect 5356 21292 5408 21301
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 7104 21292 7156 21344
rect 7196 21335 7248 21344
rect 7196 21301 7205 21335
rect 7205 21301 7239 21335
rect 7239 21301 7248 21335
rect 7196 21292 7248 21301
rect 11060 21292 11112 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 13544 21292 13596 21344
rect 14004 21292 14056 21344
rect 2663 21190 2715 21242
rect 2727 21190 2779 21242
rect 2791 21190 2843 21242
rect 2855 21190 2907 21242
rect 2919 21190 2971 21242
rect 6090 21190 6142 21242
rect 6154 21190 6206 21242
rect 6218 21190 6270 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 9517 21190 9569 21242
rect 9581 21190 9633 21242
rect 9645 21190 9697 21242
rect 9709 21190 9761 21242
rect 9773 21190 9825 21242
rect 12944 21190 12996 21242
rect 13008 21190 13060 21242
rect 13072 21190 13124 21242
rect 13136 21190 13188 21242
rect 13200 21190 13252 21242
rect 1492 21131 1544 21140
rect 1492 21097 1501 21131
rect 1501 21097 1535 21131
rect 1535 21097 1544 21131
rect 1492 21088 1544 21097
rect 4252 21088 4304 21140
rect 5908 21088 5960 21140
rect 7932 21131 7984 21140
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 9956 21088 10008 21140
rect 10876 21088 10928 21140
rect 12164 21088 12216 21140
rect 2228 20884 2280 20936
rect 3516 20995 3568 21004
rect 3516 20961 3525 20995
rect 3525 20961 3559 20995
rect 3559 20961 3568 20995
rect 3516 20952 3568 20961
rect 3608 20952 3660 21004
rect 2872 20884 2924 20936
rect 3976 20884 4028 20936
rect 1768 20859 1820 20868
rect 1768 20825 1777 20859
rect 1777 20825 1811 20859
rect 1811 20825 1820 20859
rect 1768 20816 1820 20825
rect 1860 20748 1912 20800
rect 2320 20791 2372 20800
rect 2320 20757 2329 20791
rect 2329 20757 2363 20791
rect 2363 20757 2372 20791
rect 2320 20748 2372 20757
rect 3332 20748 3384 20800
rect 4804 20791 4856 20800
rect 4804 20757 4813 20791
rect 4813 20757 4847 20791
rect 4847 20757 4856 20791
rect 4804 20748 4856 20757
rect 5264 20952 5316 21004
rect 5448 20952 5500 21004
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6184 20884 6236 20936
rect 5724 20859 5776 20868
rect 5724 20825 5733 20859
rect 5733 20825 5767 20859
rect 5767 20825 5776 20859
rect 5724 20816 5776 20825
rect 11612 21020 11664 21072
rect 7104 20884 7156 20936
rect 7380 20884 7432 20936
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 8852 20884 8904 20936
rect 9956 20884 10008 20936
rect 5264 20748 5316 20800
rect 5448 20748 5500 20800
rect 6460 20791 6512 20800
rect 6460 20757 6469 20791
rect 6469 20757 6503 20791
rect 6503 20757 6512 20791
rect 6460 20748 6512 20757
rect 7012 20748 7064 20800
rect 7656 20748 7708 20800
rect 8668 20816 8720 20868
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10968 20884 11020 20936
rect 15016 21088 15068 21140
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 12256 20884 12308 20936
rect 14096 20884 14148 20936
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 11152 20791 11204 20800
rect 11152 20757 11161 20791
rect 11161 20757 11195 20791
rect 11195 20757 11204 20791
rect 11152 20748 11204 20757
rect 12532 20748 12584 20800
rect 12808 20816 12860 20868
rect 14004 20816 14056 20868
rect 13820 20748 13872 20800
rect 4376 20646 4428 20698
rect 4440 20646 4492 20698
rect 4504 20646 4556 20698
rect 4568 20646 4620 20698
rect 4632 20646 4684 20698
rect 7803 20646 7855 20698
rect 7867 20646 7919 20698
rect 7931 20646 7983 20698
rect 7995 20646 8047 20698
rect 8059 20646 8111 20698
rect 11230 20646 11282 20698
rect 11294 20646 11346 20698
rect 11358 20646 11410 20698
rect 11422 20646 11474 20698
rect 11486 20646 11538 20698
rect 14657 20646 14709 20698
rect 14721 20646 14773 20698
rect 14785 20646 14837 20698
rect 14849 20646 14901 20698
rect 14913 20646 14965 20698
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2412 20544 2464 20596
rect 3424 20544 3476 20596
rect 3976 20587 4028 20596
rect 3976 20553 3985 20587
rect 3985 20553 4019 20587
rect 4019 20553 4028 20587
rect 3976 20544 4028 20553
rect 5540 20544 5592 20596
rect 6184 20587 6236 20596
rect 6184 20553 6193 20587
rect 6193 20553 6227 20587
rect 6227 20553 6236 20587
rect 6184 20544 6236 20553
rect 9036 20544 9088 20596
rect 10324 20544 10376 20596
rect 10968 20544 11020 20596
rect 2228 20408 2280 20460
rect 2504 20451 2556 20460
rect 2504 20417 2513 20451
rect 2513 20417 2547 20451
rect 2547 20417 2556 20451
rect 2504 20408 2556 20417
rect 2872 20451 2924 20460
rect 2872 20417 2906 20451
rect 2906 20417 2924 20451
rect 2872 20408 2924 20417
rect 4804 20476 4856 20528
rect 6460 20476 6512 20528
rect 7196 20408 7248 20460
rect 9036 20408 9088 20460
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 11060 20408 11112 20460
rect 11152 20408 11204 20460
rect 14188 20544 14240 20596
rect 11612 20476 11664 20528
rect 13544 20476 13596 20528
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 5632 20340 5684 20392
rect 940 20204 992 20256
rect 5724 20204 5776 20256
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 7472 20272 7524 20324
rect 9680 20272 9732 20324
rect 6552 20204 6604 20256
rect 7380 20204 7432 20256
rect 8208 20204 8260 20256
rect 8760 20204 8812 20256
rect 9128 20247 9180 20256
rect 9128 20213 9137 20247
rect 9137 20213 9171 20247
rect 9171 20213 9180 20247
rect 9128 20204 9180 20213
rect 9864 20204 9916 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 13452 20204 13504 20256
rect 13728 20204 13780 20256
rect 2663 20102 2715 20154
rect 2727 20102 2779 20154
rect 2791 20102 2843 20154
rect 2855 20102 2907 20154
rect 2919 20102 2971 20154
rect 6090 20102 6142 20154
rect 6154 20102 6206 20154
rect 6218 20102 6270 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 9517 20102 9569 20154
rect 9581 20102 9633 20154
rect 9645 20102 9697 20154
rect 9709 20102 9761 20154
rect 9773 20102 9825 20154
rect 12944 20102 12996 20154
rect 13008 20102 13060 20154
rect 13072 20102 13124 20154
rect 13136 20102 13188 20154
rect 13200 20102 13252 20154
rect 3884 20000 3936 20052
rect 4712 19932 4764 19984
rect 6000 20000 6052 20052
rect 6644 20000 6696 20052
rect 8116 20000 8168 20052
rect 8208 19932 8260 19984
rect 9772 20000 9824 20052
rect 9864 20000 9916 20052
rect 10692 20000 10744 20052
rect 10876 20043 10928 20052
rect 10876 20009 10885 20043
rect 10885 20009 10919 20043
rect 10919 20009 10928 20043
rect 10876 20000 10928 20009
rect 11980 20000 12032 20052
rect 3240 19864 3292 19916
rect 4068 19864 4120 19916
rect 6552 19864 6604 19916
rect 9312 19932 9364 19984
rect 10416 19932 10468 19984
rect 13728 19932 13780 19984
rect 3516 19796 3568 19848
rect 3884 19796 3936 19848
rect 4160 19796 4212 19848
rect 2228 19728 2280 19780
rect 2780 19728 2832 19780
rect 4068 19728 4120 19780
rect 4252 19771 4304 19780
rect 4252 19737 4261 19771
rect 4261 19737 4295 19771
rect 4295 19737 4304 19771
rect 4252 19728 4304 19737
rect 4804 19771 4856 19780
rect 4804 19737 4813 19771
rect 4813 19737 4847 19771
rect 4847 19737 4856 19771
rect 4804 19728 4856 19737
rect 4896 19771 4948 19780
rect 4896 19737 4905 19771
rect 4905 19737 4939 19771
rect 4939 19737 4948 19771
rect 4896 19728 4948 19737
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 1952 19660 2004 19712
rect 3056 19660 3108 19712
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 8760 19796 8812 19848
rect 6460 19728 6512 19780
rect 7012 19728 7064 19780
rect 7656 19728 7708 19780
rect 8668 19728 8720 19780
rect 10508 19796 10560 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 10784 19864 10836 19916
rect 11796 19864 11848 19916
rect 13360 19864 13412 19916
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 12532 19796 12584 19848
rect 15292 19796 15344 19848
rect 10784 19728 10836 19780
rect 11152 19728 11204 19780
rect 13268 19771 13320 19780
rect 13268 19737 13277 19771
rect 13277 19737 13311 19771
rect 13311 19737 13320 19771
rect 13268 19728 13320 19737
rect 6736 19660 6788 19712
rect 7564 19660 7616 19712
rect 8300 19660 8352 19712
rect 10232 19660 10284 19712
rect 10416 19660 10468 19712
rect 14096 19660 14148 19712
rect 14372 19660 14424 19712
rect 4376 19558 4428 19610
rect 4440 19558 4492 19610
rect 4504 19558 4556 19610
rect 4568 19558 4620 19610
rect 4632 19558 4684 19610
rect 7803 19558 7855 19610
rect 7867 19558 7919 19610
rect 7931 19558 7983 19610
rect 7995 19558 8047 19610
rect 8059 19558 8111 19610
rect 11230 19558 11282 19610
rect 11294 19558 11346 19610
rect 11358 19558 11410 19610
rect 11422 19558 11474 19610
rect 11486 19558 11538 19610
rect 14657 19558 14709 19610
rect 14721 19558 14773 19610
rect 14785 19558 14837 19610
rect 14849 19558 14901 19610
rect 14913 19558 14965 19610
rect 3976 19456 4028 19508
rect 4068 19456 4120 19508
rect 4896 19456 4948 19508
rect 6092 19499 6144 19508
rect 6092 19465 6101 19499
rect 6101 19465 6135 19499
rect 6135 19465 6144 19499
rect 6092 19456 6144 19465
rect 6920 19456 6972 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 2780 19388 2832 19440
rect 3332 19388 3384 19440
rect 7656 19499 7708 19508
rect 7656 19465 7665 19499
rect 7665 19465 7699 19499
rect 7699 19465 7708 19499
rect 7656 19456 7708 19465
rect 8484 19456 8536 19508
rect 9404 19499 9456 19508
rect 9404 19465 9413 19499
rect 9413 19465 9447 19499
rect 9447 19465 9456 19499
rect 9404 19456 9456 19465
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 9772 19456 9824 19508
rect 10692 19456 10744 19508
rect 11520 19456 11572 19508
rect 11704 19456 11756 19508
rect 12624 19456 12676 19508
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 14188 19499 14240 19508
rect 14188 19465 14197 19499
rect 14197 19465 14231 19499
rect 14231 19465 14240 19499
rect 14188 19456 14240 19465
rect 14556 19456 14608 19508
rect 8300 19431 8352 19440
rect 4712 19320 4764 19372
rect 2412 19252 2464 19304
rect 3516 19295 3568 19304
rect 3516 19261 3525 19295
rect 3525 19261 3559 19295
rect 3559 19261 3568 19295
rect 3516 19252 3568 19261
rect 4344 19295 4396 19304
rect 4344 19261 4353 19295
rect 4353 19261 4387 19295
rect 4387 19261 4396 19295
rect 4344 19252 4396 19261
rect 4896 19252 4948 19304
rect 5724 19320 5776 19372
rect 8300 19397 8309 19431
rect 8309 19397 8343 19431
rect 8343 19397 8352 19431
rect 8300 19388 8352 19397
rect 8576 19388 8628 19440
rect 2228 19184 2280 19236
rect 3608 19184 3660 19236
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 6552 19252 6604 19304
rect 7564 19252 7616 19304
rect 9864 19388 9916 19440
rect 10140 19388 10192 19440
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 11612 19388 11664 19440
rect 12072 19388 12124 19440
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 10140 19252 10192 19304
rect 10416 19252 10468 19304
rect 11060 19320 11112 19372
rect 12256 19320 12308 19372
rect 12348 19320 12400 19372
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 14004 19320 14056 19372
rect 14556 19320 14608 19372
rect 7840 19184 7892 19236
rect 7932 19184 7984 19236
rect 940 19116 992 19168
rect 2136 19159 2188 19168
rect 2136 19125 2145 19159
rect 2145 19125 2179 19159
rect 2179 19125 2188 19159
rect 2136 19116 2188 19125
rect 5908 19116 5960 19168
rect 8300 19116 8352 19168
rect 8392 19116 8444 19168
rect 8944 19116 8996 19168
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 11888 19252 11940 19304
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 2663 19014 2715 19066
rect 2727 19014 2779 19066
rect 2791 19014 2843 19066
rect 2855 19014 2907 19066
rect 2919 19014 2971 19066
rect 6090 19014 6142 19066
rect 6154 19014 6206 19066
rect 6218 19014 6270 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 9517 19014 9569 19066
rect 9581 19014 9633 19066
rect 9645 19014 9697 19066
rect 9709 19014 9761 19066
rect 9773 19014 9825 19066
rect 12944 19014 12996 19066
rect 13008 19014 13060 19066
rect 13072 19014 13124 19066
rect 13136 19014 13188 19066
rect 13200 19014 13252 19066
rect 1952 18912 2004 18964
rect 2044 18912 2096 18964
rect 3516 18912 3568 18964
rect 4160 18955 4212 18964
rect 4160 18921 4169 18955
rect 4169 18921 4203 18955
rect 4203 18921 4212 18955
rect 4160 18912 4212 18921
rect 4436 18955 4488 18964
rect 4436 18921 4445 18955
rect 4445 18921 4479 18955
rect 4479 18921 4488 18955
rect 4436 18912 4488 18921
rect 2320 18776 2372 18828
rect 3424 18776 3476 18828
rect 1860 18751 1912 18760
rect 1860 18717 1869 18751
rect 1869 18717 1903 18751
rect 1903 18717 1912 18751
rect 1860 18708 1912 18717
rect 2228 18708 2280 18760
rect 2320 18572 2372 18624
rect 3792 18708 3844 18760
rect 3884 18708 3936 18760
rect 8392 18912 8444 18964
rect 5632 18776 5684 18828
rect 6644 18776 6696 18828
rect 7932 18887 7984 18896
rect 7932 18853 7941 18887
rect 7941 18853 7975 18887
rect 7975 18853 7984 18887
rect 7932 18844 7984 18853
rect 8116 18776 8168 18828
rect 7564 18708 7616 18760
rect 7656 18708 7708 18760
rect 7840 18708 7892 18760
rect 8576 18844 8628 18896
rect 9864 18912 9916 18964
rect 11612 18955 11664 18964
rect 11612 18921 11621 18955
rect 11621 18921 11655 18955
rect 11655 18921 11664 18955
rect 11612 18912 11664 18921
rect 12164 18912 12216 18964
rect 12348 18912 12400 18964
rect 12716 18912 12768 18964
rect 13912 18912 13964 18964
rect 8944 18844 8996 18896
rect 10140 18776 10192 18828
rect 10324 18776 10376 18828
rect 10692 18776 10744 18828
rect 8944 18708 8996 18760
rect 9680 18708 9732 18760
rect 10600 18708 10652 18760
rect 10968 18751 11020 18760
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 11060 18708 11112 18760
rect 14096 18844 14148 18896
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 13728 18708 13780 18760
rect 15200 18708 15252 18760
rect 5540 18640 5592 18692
rect 6276 18683 6328 18692
rect 6276 18649 6285 18683
rect 6285 18649 6319 18683
rect 6319 18649 6328 18683
rect 6276 18640 6328 18649
rect 7288 18640 7340 18692
rect 6000 18615 6052 18624
rect 6000 18581 6009 18615
rect 6009 18581 6043 18615
rect 6043 18581 6052 18615
rect 6000 18572 6052 18581
rect 7196 18572 7248 18624
rect 8484 18572 8536 18624
rect 12072 18572 12124 18624
rect 12900 18683 12952 18692
rect 12900 18649 12909 18683
rect 12909 18649 12943 18683
rect 12943 18649 12952 18683
rect 12900 18640 12952 18649
rect 14188 18572 14240 18624
rect 14464 18572 14516 18624
rect 4376 18470 4428 18522
rect 4440 18470 4492 18522
rect 4504 18470 4556 18522
rect 4568 18470 4620 18522
rect 4632 18470 4684 18522
rect 7803 18470 7855 18522
rect 7867 18470 7919 18522
rect 7931 18470 7983 18522
rect 7995 18470 8047 18522
rect 8059 18470 8111 18522
rect 11230 18470 11282 18522
rect 11294 18470 11346 18522
rect 11358 18470 11410 18522
rect 11422 18470 11474 18522
rect 11486 18470 11538 18522
rect 14657 18470 14709 18522
rect 14721 18470 14773 18522
rect 14785 18470 14837 18522
rect 14849 18470 14901 18522
rect 14913 18470 14965 18522
rect 2320 18411 2372 18420
rect 2320 18377 2329 18411
rect 2329 18377 2363 18411
rect 2363 18377 2372 18411
rect 2320 18368 2372 18377
rect 3608 18368 3660 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 1584 18232 1636 18284
rect 2136 18232 2188 18284
rect 6276 18300 6328 18352
rect 6460 18343 6512 18352
rect 6460 18309 6469 18343
rect 6469 18309 6503 18343
rect 6503 18309 6512 18343
rect 6460 18300 6512 18309
rect 6552 18343 6604 18352
rect 6552 18309 6561 18343
rect 6561 18309 6595 18343
rect 6595 18309 6604 18343
rect 6552 18300 6604 18309
rect 7196 18300 7248 18352
rect 3516 18232 3568 18284
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 5540 18232 5592 18284
rect 2228 18164 2280 18216
rect 3240 18164 3292 18216
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2412 18028 2464 18080
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 3332 18028 3384 18080
rect 6000 18164 6052 18216
rect 6460 18164 6512 18216
rect 8300 18368 8352 18420
rect 10968 18368 11020 18420
rect 12164 18368 12216 18420
rect 8944 18300 8996 18352
rect 5908 18096 5960 18148
rect 4068 18028 4120 18080
rect 5540 18071 5592 18080
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 7288 18096 7340 18148
rect 8116 18096 8168 18148
rect 9220 18232 9272 18284
rect 11060 18300 11112 18352
rect 9404 18164 9456 18216
rect 10416 18232 10468 18284
rect 10600 18232 10652 18284
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 10324 18164 10376 18216
rect 9680 18096 9732 18148
rect 10876 18207 10928 18216
rect 10876 18173 10885 18207
rect 10885 18173 10919 18207
rect 10919 18173 10928 18207
rect 10876 18164 10928 18173
rect 11060 18164 11112 18216
rect 11704 18232 11756 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 13912 18343 13964 18352
rect 13912 18309 13921 18343
rect 13921 18309 13955 18343
rect 13955 18309 13964 18343
rect 13912 18300 13964 18309
rect 11612 18164 11664 18216
rect 12532 18232 12584 18284
rect 12348 18164 12400 18216
rect 13452 18164 13504 18216
rect 10968 18096 11020 18148
rect 11888 18096 11940 18148
rect 12256 18139 12308 18148
rect 12256 18105 12265 18139
rect 12265 18105 12299 18139
rect 12299 18105 12308 18139
rect 12256 18096 12308 18105
rect 6828 18028 6880 18080
rect 8024 18028 8076 18080
rect 9864 18028 9916 18080
rect 11704 18028 11756 18080
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14464 18028 14516 18080
rect 2663 17926 2715 17978
rect 2727 17926 2779 17978
rect 2791 17926 2843 17978
rect 2855 17926 2907 17978
rect 2919 17926 2971 17978
rect 6090 17926 6142 17978
rect 6154 17926 6206 17978
rect 6218 17926 6270 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 9517 17926 9569 17978
rect 9581 17926 9633 17978
rect 9645 17926 9697 17978
rect 9709 17926 9761 17978
rect 9773 17926 9825 17978
rect 12944 17926 12996 17978
rect 13008 17926 13060 17978
rect 13072 17926 13124 17978
rect 13136 17926 13188 17978
rect 13200 17926 13252 17978
rect 2412 17867 2464 17876
rect 2412 17833 2421 17867
rect 2421 17833 2455 17867
rect 2455 17833 2464 17867
rect 2412 17824 2464 17833
rect 3332 17824 3384 17876
rect 3884 17824 3936 17876
rect 7656 17824 7708 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9312 17824 9364 17876
rect 10048 17824 10100 17876
rect 10140 17824 10192 17876
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 3240 17688 3292 17740
rect 8300 17688 8352 17740
rect 940 17620 992 17672
rect 2872 17620 2924 17672
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 1768 17595 1820 17604
rect 1768 17561 1777 17595
rect 1777 17561 1811 17595
rect 1811 17561 1820 17595
rect 1768 17552 1820 17561
rect 4160 17620 4212 17672
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 7104 17620 7156 17672
rect 8024 17620 8076 17672
rect 5540 17552 5592 17604
rect 10232 17756 10284 17808
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 9864 17620 9916 17672
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 2964 17484 3016 17536
rect 3608 17484 3660 17536
rect 3884 17484 3936 17536
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 7012 17484 7064 17536
rect 7196 17484 7248 17536
rect 8668 17484 8720 17536
rect 10140 17552 10192 17604
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 12624 17824 12676 17876
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 10876 17552 10928 17604
rect 11980 17552 12032 17604
rect 12348 17620 12400 17672
rect 12164 17552 12216 17604
rect 10232 17527 10284 17536
rect 10232 17493 10241 17527
rect 10241 17493 10275 17527
rect 10275 17493 10284 17527
rect 10232 17484 10284 17493
rect 10692 17484 10744 17536
rect 13636 17663 13688 17672
rect 13636 17629 13645 17663
rect 13645 17629 13679 17663
rect 13679 17629 13688 17663
rect 13636 17620 13688 17629
rect 14004 17620 14056 17672
rect 12716 17484 12768 17536
rect 13452 17484 13504 17536
rect 13728 17527 13780 17536
rect 13728 17493 13737 17527
rect 13737 17493 13771 17527
rect 13771 17493 13780 17527
rect 13728 17484 13780 17493
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 1400 17280 1452 17332
rect 3424 17280 3476 17332
rect 4252 17280 4304 17332
rect 4896 17280 4948 17332
rect 6552 17280 6604 17332
rect 6920 17280 6972 17332
rect 9128 17280 9180 17332
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 2964 17187 3016 17196
rect 2964 17153 2998 17187
rect 2998 17153 3016 17187
rect 2964 17144 3016 17153
rect 7104 17212 7156 17264
rect 5816 17144 5868 17196
rect 10416 17255 10468 17264
rect 10416 17221 10425 17255
rect 10425 17221 10459 17255
rect 10459 17221 10468 17255
rect 10416 17212 10468 17221
rect 10508 17212 10560 17264
rect 10968 17212 11020 17264
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 5632 17008 5684 17060
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 8024 17076 8076 17128
rect 8300 17076 8352 17128
rect 940 16940 992 16992
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 4804 16940 4856 16992
rect 6920 16940 6972 16992
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 7564 16940 7616 16992
rect 9864 17076 9916 17128
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11428 17212 11480 17264
rect 11980 17280 12032 17332
rect 12440 17280 12492 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 13268 17212 13320 17264
rect 10508 17076 10560 17128
rect 11520 17187 11572 17196
rect 11520 17153 11537 17187
rect 11537 17153 11571 17187
rect 11571 17153 11572 17187
rect 11520 17144 11572 17153
rect 14372 17144 14424 17196
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 12164 17076 12216 17128
rect 12348 17076 12400 17128
rect 10876 17051 10928 17060
rect 10876 17017 10885 17051
rect 10885 17017 10919 17051
rect 10919 17017 10928 17051
rect 10876 17008 10928 17017
rect 11060 17008 11112 17060
rect 11980 17008 12032 17060
rect 12808 17119 12860 17128
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 12348 16940 12400 16992
rect 12440 16940 12492 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 3700 16736 3752 16788
rect 3884 16736 3936 16788
rect 3148 16668 3200 16720
rect 4068 16668 4120 16720
rect 4160 16668 4212 16720
rect 1584 16600 1636 16652
rect 2504 16507 2556 16516
rect 2504 16473 2522 16507
rect 2522 16473 2556 16507
rect 2504 16464 2556 16473
rect 2964 16532 3016 16584
rect 1400 16439 1452 16448
rect 1400 16405 1409 16439
rect 1409 16405 1443 16439
rect 1443 16405 1452 16439
rect 1400 16396 1452 16405
rect 2964 16396 3016 16448
rect 3700 16532 3752 16584
rect 3884 16575 3936 16584
rect 3884 16541 3893 16575
rect 3893 16541 3927 16575
rect 3927 16541 3936 16575
rect 3884 16532 3936 16541
rect 4252 16532 4304 16584
rect 7380 16736 7432 16788
rect 9128 16736 9180 16788
rect 10232 16736 10284 16788
rect 5632 16600 5684 16652
rect 4804 16532 4856 16584
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 7472 16600 7524 16652
rect 8024 16600 8076 16652
rect 6736 16532 6788 16584
rect 4712 16396 4764 16448
rect 4988 16439 5040 16448
rect 4988 16405 4997 16439
rect 4997 16405 5031 16439
rect 5031 16405 5040 16439
rect 4988 16396 5040 16405
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 5724 16396 5776 16448
rect 6000 16396 6052 16448
rect 6644 16464 6696 16516
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 7656 16396 7708 16448
rect 8760 16532 8812 16584
rect 11520 16668 11572 16720
rect 12808 16736 12860 16788
rect 13268 16736 13320 16788
rect 12072 16643 12124 16652
rect 9956 16532 10008 16584
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 9036 16464 9088 16516
rect 12348 16532 12400 16584
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 8668 16396 8720 16448
rect 10140 16507 10192 16516
rect 10140 16473 10174 16507
rect 10174 16473 10192 16507
rect 10140 16464 10192 16473
rect 12164 16464 12216 16516
rect 13452 16464 13504 16516
rect 14280 16532 14332 16584
rect 15016 16532 15068 16584
rect 9588 16439 9640 16448
rect 9588 16405 9597 16439
rect 9597 16405 9631 16439
rect 9631 16405 9640 16439
rect 9588 16396 9640 16405
rect 11796 16396 11848 16448
rect 12348 16439 12400 16448
rect 12348 16405 12357 16439
rect 12357 16405 12391 16439
rect 12391 16405 12400 16439
rect 12348 16396 12400 16405
rect 13268 16396 13320 16448
rect 13912 16396 13964 16448
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 1400 16192 1452 16244
rect 2780 16192 2832 16244
rect 3884 16192 3936 16244
rect 4712 16192 4764 16244
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 3424 16056 3476 16108
rect 4344 16124 4396 16176
rect 4804 16167 4856 16176
rect 4804 16133 4813 16167
rect 4813 16133 4847 16167
rect 4847 16133 4856 16167
rect 4804 16124 4856 16133
rect 4988 16192 5040 16244
rect 6736 16192 6788 16244
rect 7380 16192 7432 16244
rect 9312 16192 9364 16244
rect 9588 16192 9640 16244
rect 12532 16192 12584 16244
rect 12716 16192 12768 16244
rect 13452 16192 13504 16244
rect 13912 16192 13964 16244
rect 5724 16124 5776 16176
rect 9956 16124 10008 16176
rect 8392 16056 8444 16108
rect 10324 16099 10376 16108
rect 10324 16065 10342 16099
rect 10342 16065 10376 16099
rect 10324 16056 10376 16065
rect 10876 16099 10928 16108
rect 10876 16065 10885 16099
rect 10885 16065 10919 16099
rect 10919 16065 10928 16099
rect 10876 16056 10928 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 13820 16124 13872 16176
rect 11796 16099 11848 16108
rect 11796 16065 11830 16099
rect 11830 16065 11848 16099
rect 11796 16056 11848 16065
rect 2964 15988 3016 16040
rect 3148 15920 3200 15972
rect 3608 15920 3660 15972
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 7564 15988 7616 16040
rect 8300 16031 8352 16040
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 10968 15988 11020 16040
rect 940 15852 992 15904
rect 2412 15852 2464 15904
rect 3056 15852 3108 15904
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 8760 15852 8812 15904
rect 9220 15895 9272 15904
rect 9220 15861 9229 15895
rect 9229 15861 9263 15895
rect 9263 15861 9272 15895
rect 9220 15852 9272 15861
rect 13636 16056 13688 16108
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 13268 15988 13320 16040
rect 12716 15920 12768 15972
rect 13268 15852 13320 15904
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 2504 15648 2556 15700
rect 3148 15648 3200 15700
rect 3608 15648 3660 15700
rect 3700 15648 3752 15700
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 4252 15648 4304 15700
rect 4804 15691 4856 15700
rect 4804 15657 4813 15691
rect 4813 15657 4847 15691
rect 4847 15657 4856 15691
rect 4804 15648 4856 15657
rect 5172 15648 5224 15700
rect 6644 15648 6696 15700
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 7656 15648 7708 15700
rect 8392 15648 8444 15700
rect 8576 15648 8628 15700
rect 13360 15648 13412 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2228 15512 2280 15564
rect 2504 15444 2556 15496
rect 2136 15376 2188 15428
rect 3424 15376 3476 15428
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 3792 15376 3844 15428
rect 6000 15580 6052 15632
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 10784 15623 10836 15632
rect 10784 15589 10793 15623
rect 10793 15589 10827 15623
rect 10827 15589 10836 15623
rect 10784 15580 10836 15589
rect 11152 15580 11204 15632
rect 12348 15580 12400 15632
rect 12808 15623 12860 15632
rect 12808 15589 12817 15623
rect 12817 15589 12851 15623
rect 12851 15589 12860 15623
rect 12808 15580 12860 15589
rect 9036 15444 9088 15496
rect 9220 15444 9272 15496
rect 10232 15512 10284 15564
rect 10416 15512 10468 15564
rect 10968 15444 11020 15496
rect 11612 15512 11664 15564
rect 11888 15512 11940 15564
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 9680 15376 9732 15428
rect 11060 15376 11112 15428
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 13268 15376 13320 15428
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9128 15308 9180 15360
rect 10048 15308 10100 15360
rect 11612 15308 11664 15360
rect 13912 15419 13964 15428
rect 13912 15385 13921 15419
rect 13921 15385 13955 15419
rect 13955 15385 13964 15419
rect 13912 15376 13964 15385
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 2044 15104 2096 15156
rect 1584 14968 1636 15020
rect 2228 15036 2280 15088
rect 2412 15036 2464 15088
rect 3608 15104 3660 15156
rect 4896 15104 4948 15156
rect 8392 15104 8444 15156
rect 9680 15104 9732 15156
rect 10140 15104 10192 15156
rect 11704 15104 11756 15156
rect 12440 15104 12492 15156
rect 13728 15104 13780 15156
rect 3056 14968 3108 15020
rect 3240 14968 3292 15020
rect 3792 14968 3844 15020
rect 5264 15036 5316 15088
rect 10784 15036 10836 15088
rect 11152 15079 11204 15088
rect 11152 15045 11161 15079
rect 11161 15045 11195 15079
rect 11195 15045 11204 15079
rect 11152 15036 11204 15045
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 7564 14968 7616 15020
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 13636 15079 13688 15088
rect 13636 15045 13654 15079
rect 13654 15045 13688 15079
rect 13636 15036 13688 15045
rect 12072 14968 12124 15020
rect 12532 14968 12584 15020
rect 13820 14968 13872 15020
rect 1124 14832 1176 14884
rect 3240 14832 3292 14884
rect 2504 14764 2556 14816
rect 6920 14900 6972 14952
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8576 14943 8628 14952
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 9404 14900 9456 14952
rect 9864 14900 9916 14952
rect 10968 14900 11020 14952
rect 14280 14832 14332 14884
rect 4252 14764 4304 14816
rect 4712 14807 4764 14816
rect 4712 14773 4721 14807
rect 4721 14773 4755 14807
rect 4755 14773 4764 14807
rect 4712 14764 4764 14773
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 11704 14764 11756 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 1492 14560 1544 14612
rect 4252 14560 4304 14612
rect 4344 14560 4396 14612
rect 4896 14560 4948 14612
rect 7472 14560 7524 14612
rect 7840 14560 7892 14612
rect 8300 14560 8352 14612
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 9864 14560 9916 14612
rect 11704 14560 11756 14612
rect 12440 14560 12492 14612
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 940 14356 992 14408
rect 2412 14356 2464 14408
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 3332 14424 3384 14476
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 7564 14424 7616 14476
rect 4252 14288 4304 14340
rect 4528 14288 4580 14340
rect 5540 14356 5592 14408
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 10048 14492 10100 14544
rect 8944 14356 8996 14408
rect 10416 14424 10468 14476
rect 10876 14424 10928 14476
rect 11612 14424 11664 14476
rect 12716 14424 12768 14476
rect 13912 14492 13964 14544
rect 10048 14356 10100 14408
rect 12164 14356 12216 14408
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 2872 14220 2924 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 3608 14220 3660 14272
rect 4804 14263 4856 14272
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 5724 14220 5776 14272
rect 7104 14220 7156 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 11612 14220 11664 14272
rect 11980 14220 12032 14272
rect 13728 14220 13780 14272
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 1400 14016 1452 14068
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4804 14016 4856 14068
rect 4160 13948 4212 14000
rect 5540 14016 5592 14068
rect 7472 14016 7524 14068
rect 7564 14059 7616 14068
rect 7564 14025 7573 14059
rect 7573 14025 7607 14059
rect 7607 14025 7616 14059
rect 7564 14016 7616 14025
rect 1584 13812 1636 13864
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 4712 13880 4764 13932
rect 4896 13787 4948 13796
rect 4896 13753 4905 13787
rect 4905 13753 4939 13787
rect 4939 13753 4948 13787
rect 4896 13744 4948 13753
rect 6460 13880 6512 13932
rect 8760 14016 8812 14068
rect 10048 14016 10100 14068
rect 10324 14016 10376 14068
rect 10876 14016 10928 14068
rect 10968 14016 11020 14068
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 7748 13880 7800 13889
rect 9128 13880 9180 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9312 13880 9364 13932
rect 9956 13880 10008 13932
rect 11152 13948 11204 14000
rect 11612 14016 11664 14068
rect 12440 14016 12492 14068
rect 13360 14016 13412 14068
rect 14096 14016 14148 14068
rect 11244 13880 11296 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 6736 13812 6788 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7196 13812 7248 13864
rect 7380 13812 7432 13864
rect 10784 13812 10836 13864
rect 11152 13812 11204 13864
rect 11888 13812 11940 13864
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 12624 13812 12676 13864
rect 13268 13812 13320 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 5724 13676 5776 13728
rect 14464 13676 14516 13728
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 2044 13472 2096 13524
rect 2228 13472 2280 13524
rect 3516 13472 3568 13524
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 1952 13404 2004 13456
rect 2412 13336 2464 13388
rect 4068 13404 4120 13456
rect 6644 13472 6696 13524
rect 6736 13472 6788 13524
rect 4988 13404 5040 13456
rect 7012 13404 7064 13456
rect 1952 13268 2004 13320
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 3516 13268 3568 13320
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4804 13268 4856 13320
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 7288 13336 7340 13388
rect 7748 13472 7800 13524
rect 8484 13472 8536 13524
rect 10140 13472 10192 13524
rect 10968 13515 11020 13524
rect 10968 13481 10977 13515
rect 10977 13481 11011 13515
rect 11011 13481 11020 13515
rect 10968 13472 11020 13481
rect 12624 13472 12676 13524
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 10048 13404 10100 13456
rect 10784 13404 10836 13456
rect 8760 13336 8812 13388
rect 9312 13336 9364 13388
rect 8208 13268 8260 13320
rect 11244 13336 11296 13388
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 1584 13200 1636 13252
rect 1676 13200 1728 13252
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 5264 13132 5316 13184
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 7472 13200 7524 13252
rect 7656 13243 7708 13252
rect 7656 13209 7690 13243
rect 7690 13209 7708 13243
rect 7656 13200 7708 13209
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 11888 13268 11940 13320
rect 12072 13268 12124 13320
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 13268 13268 13320 13320
rect 8576 13132 8628 13184
rect 8944 13132 8996 13184
rect 9128 13132 9180 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 11980 13132 12032 13184
rect 13544 13200 13596 13252
rect 14004 13200 14056 13252
rect 13820 13132 13872 13184
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 1860 12928 1912 12980
rect 2320 12928 2372 12980
rect 3240 12928 3292 12980
rect 3332 12928 3384 12980
rect 3976 12928 4028 12980
rect 4252 12928 4304 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 2412 12860 2464 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2504 12724 2556 12776
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 4528 12792 4580 12844
rect 5632 12792 5684 12844
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 3056 12724 3108 12733
rect 3608 12724 3660 12776
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 6828 12928 6880 12980
rect 7104 12928 7156 12980
rect 7288 12928 7340 12980
rect 7472 12928 7524 12980
rect 9220 12928 9272 12980
rect 9680 12928 9732 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11060 12928 11112 12980
rect 8300 12860 8352 12912
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 8944 12792 8996 12844
rect 11888 12928 11940 12980
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 10232 12792 10284 12844
rect 12072 12860 12124 12912
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 10968 12724 11020 12776
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 11888 12724 11940 12776
rect 12440 12724 12492 12776
rect 15200 12792 15252 12844
rect 15292 12656 15344 12708
rect 4068 12588 4120 12640
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 11980 12588 12032 12640
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 12808 12588 12860 12640
rect 14924 12588 14976 12640
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 2136 12384 2188 12436
rect 12440 12384 12492 12436
rect 12532 12384 12584 12436
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 940 12180 992 12232
rect 4436 12316 4488 12368
rect 4620 12359 4672 12368
rect 4620 12325 4629 12359
rect 4629 12325 4663 12359
rect 4663 12325 4672 12359
rect 4620 12316 4672 12325
rect 5356 12316 5408 12368
rect 5632 12316 5684 12368
rect 7840 12359 7892 12368
rect 7840 12325 7849 12359
rect 7849 12325 7883 12359
rect 7883 12325 7892 12359
rect 7840 12316 7892 12325
rect 10324 12316 10376 12368
rect 10416 12359 10468 12368
rect 10416 12325 10425 12359
rect 10425 12325 10459 12359
rect 10459 12325 10468 12359
rect 10416 12316 10468 12325
rect 12348 12316 12400 12368
rect 1860 12248 1912 12300
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 5172 12248 5224 12300
rect 5540 12248 5592 12300
rect 6092 12248 6144 12300
rect 7380 12248 7432 12300
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8576 12248 8628 12300
rect 9220 12248 9272 12300
rect 1952 12180 2004 12232
rect 2044 12112 2096 12164
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 1492 12044 1544 12096
rect 2504 12044 2556 12096
rect 3700 12044 3752 12096
rect 4528 12112 4580 12164
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5908 12180 5960 12232
rect 6460 12180 6512 12232
rect 5080 12044 5132 12096
rect 5264 12155 5316 12164
rect 5264 12121 5273 12155
rect 5273 12121 5307 12155
rect 5307 12121 5316 12155
rect 5264 12112 5316 12121
rect 5356 12112 5408 12164
rect 6000 12112 6052 12164
rect 6736 12112 6788 12164
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 9220 12112 9272 12164
rect 11060 12180 11112 12232
rect 11704 12180 11756 12232
rect 12532 12248 12584 12300
rect 13452 12248 13504 12300
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 8852 12044 8904 12096
rect 9404 12044 9456 12096
rect 11888 12112 11940 12164
rect 12624 12180 12676 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13360 12112 13412 12164
rect 12440 12044 12492 12096
rect 15016 12180 15068 12232
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3148 11840 3200 11892
rect 5080 11840 5132 11892
rect 1860 11704 1912 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2964 11704 3016 11756
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 6092 11747 6144 11756
rect 6092 11713 6101 11747
rect 6101 11713 6135 11747
rect 6135 11713 6144 11747
rect 6092 11704 6144 11713
rect 6276 11704 6328 11756
rect 7288 11840 7340 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 10968 11840 11020 11892
rect 6644 11772 6696 11824
rect 8760 11704 8812 11756
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12532 11840 12584 11892
rect 12992 11840 13044 11892
rect 13360 11840 13412 11892
rect 13636 11840 13688 11892
rect 5080 11568 5132 11620
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5908 11500 5960 11552
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 8852 11636 8904 11688
rect 12440 11704 12492 11756
rect 12716 11704 12768 11756
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 12164 11636 12216 11688
rect 12624 11636 12676 11688
rect 13268 11636 13320 11688
rect 7196 11568 7248 11620
rect 8300 11568 8352 11620
rect 9220 11568 9272 11620
rect 11060 11568 11112 11620
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 14004 11500 14056 11552
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 1676 11296 1728 11348
rect 1860 11296 1912 11348
rect 2228 11296 2280 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 4804 11228 4856 11280
rect 7012 11228 7064 11280
rect 2504 11160 2556 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 1952 11092 2004 11144
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 1860 11024 1912 11076
rect 2228 11024 2280 11076
rect 2412 11024 2464 11076
rect 5080 11024 5132 11076
rect 5540 11092 5592 11144
rect 7012 11092 7064 11144
rect 10324 11296 10376 11348
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 11520 11296 11572 11348
rect 11888 11296 11940 11348
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 12440 11160 12492 11212
rect 10232 11092 10284 11144
rect 5724 11067 5776 11076
rect 5724 11033 5758 11067
rect 5758 11033 5776 11067
rect 5724 11024 5776 11033
rect 2136 10956 2188 11008
rect 3976 10956 4028 11008
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 7288 10956 7340 11008
rect 8208 10956 8260 11008
rect 11428 11092 11480 11144
rect 12072 11092 12124 11144
rect 12808 11160 12860 11212
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 12624 11024 12676 11076
rect 14096 11092 14148 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 13728 11024 13780 11076
rect 14372 11160 14424 11212
rect 14464 11024 14516 11076
rect 11612 10956 11664 11008
rect 13360 10956 13412 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 2044 10752 2096 10804
rect 2504 10752 2556 10804
rect 3148 10752 3200 10804
rect 5724 10752 5776 10804
rect 8760 10752 8812 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 1308 10548 1360 10600
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 1952 10548 2004 10600
rect 2136 10548 2188 10600
rect 3056 10548 3108 10600
rect 4344 10616 4396 10668
rect 4528 10616 4580 10668
rect 5908 10616 5960 10668
rect 3976 10548 4028 10600
rect 5356 10480 5408 10532
rect 7472 10684 7524 10736
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 14004 10752 14056 10804
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 6920 10548 6972 10600
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 8760 10548 8812 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 1768 10412 1820 10464
rect 3516 10412 3568 10464
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4252 10412 4304 10464
rect 4528 10412 4580 10464
rect 5264 10412 5316 10464
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 14556 10684 14608 10736
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 11796 10616 11848 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 11428 10548 11480 10600
rect 13268 10616 13320 10668
rect 13820 10616 13872 10668
rect 14280 10616 14332 10668
rect 12992 10523 13044 10532
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13636 10412 13688 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 1584 10208 1636 10260
rect 3332 10208 3384 10260
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 3976 10208 4028 10260
rect 4068 10140 4120 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 2504 9979 2556 9988
rect 2504 9945 2538 9979
rect 2538 9945 2556 9979
rect 2504 9936 2556 9945
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5448 10208 5500 10260
rect 7656 10208 7708 10260
rect 8576 10208 8628 10260
rect 8668 10208 8720 10260
rect 9864 10208 9916 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 11428 10208 11480 10260
rect 12532 10208 12584 10260
rect 12716 10208 12768 10260
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 5632 10004 5684 10056
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 8484 10072 8536 10124
rect 13636 10208 13688 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 4344 9868 4396 9920
rect 5172 9868 5224 9920
rect 7196 9936 7248 9988
rect 7656 9936 7708 9988
rect 8852 10004 8904 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 8668 9868 8720 9920
rect 9864 10004 9916 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10140 9911 10192 9920
rect 10140 9877 10149 9911
rect 10149 9877 10183 9911
rect 10183 9877 10192 9911
rect 10140 9868 10192 9877
rect 11612 10004 11664 10056
rect 13912 10004 13964 10056
rect 13360 9936 13412 9988
rect 12164 9868 12216 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 3240 9664 3292 9716
rect 3792 9664 3844 9716
rect 3976 9664 4028 9716
rect 1860 9528 1912 9580
rect 940 9460 992 9512
rect 2136 9460 2188 9512
rect 3332 9392 3384 9444
rect 3884 9528 3936 9580
rect 5724 9596 5776 9648
rect 6460 9664 6512 9716
rect 7472 9664 7524 9716
rect 8760 9664 8812 9716
rect 9220 9664 9272 9716
rect 10232 9664 10284 9716
rect 4160 9324 4212 9376
rect 5448 9528 5500 9580
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 5080 9460 5132 9512
rect 5632 9460 5684 9512
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 8392 9528 8444 9580
rect 8484 9528 8536 9580
rect 9864 9596 9916 9648
rect 13912 9664 13964 9716
rect 7656 9392 7708 9444
rect 10140 9528 10192 9580
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12624 9528 12676 9580
rect 14004 9528 14056 9580
rect 12532 9460 12584 9512
rect 13452 9503 13504 9512
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 13544 9460 13596 9512
rect 13912 9460 13964 9512
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 5264 9324 5316 9376
rect 5816 9324 5868 9376
rect 6460 9324 6512 9376
rect 7196 9324 7248 9376
rect 7288 9324 7340 9376
rect 8576 9324 8628 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 3240 9120 3292 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 3884 9120 3936 9172
rect 4712 9120 4764 9172
rect 4988 9120 5040 9172
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 6460 9120 6512 9172
rect 7196 9120 7248 9172
rect 3056 9052 3108 9104
rect 3332 9052 3384 9104
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 2136 8780 2188 8832
rect 2688 8848 2740 8900
rect 3240 8916 3292 8968
rect 4160 8984 4212 9036
rect 5264 9052 5316 9104
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 3608 8916 3660 8925
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4712 8916 4764 8968
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5264 8916 5316 8968
rect 4344 8848 4396 8900
rect 3516 8780 3568 8832
rect 3976 8780 4028 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 4988 8891 5040 8900
rect 4988 8857 4997 8891
rect 4997 8857 5031 8891
rect 5031 8857 5040 8891
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 8760 9120 8812 9172
rect 10416 9120 10468 9172
rect 11888 9120 11940 9172
rect 8300 8984 8352 9036
rect 9220 8984 9272 9036
rect 4988 8848 5040 8857
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 8392 8916 8444 8968
rect 10324 9052 10376 9104
rect 11152 9052 11204 9104
rect 12164 8984 12216 9036
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 5172 8780 5224 8832
rect 6460 8780 6512 8832
rect 9128 8848 9180 8900
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8576 8780 8628 8832
rect 12808 8984 12860 9036
rect 13452 9120 13504 9172
rect 14004 9120 14056 9172
rect 14188 9120 14240 9172
rect 13452 8916 13504 8968
rect 14188 8916 14240 8968
rect 10692 8780 10744 8832
rect 10968 8891 11020 8900
rect 10968 8857 10977 8891
rect 10977 8857 11011 8891
rect 11011 8857 11020 8891
rect 10968 8848 11020 8857
rect 12164 8891 12216 8900
rect 12164 8857 12173 8891
rect 12173 8857 12207 8891
rect 12207 8857 12216 8891
rect 12164 8848 12216 8857
rect 11796 8780 11848 8832
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 12624 8780 12676 8832
rect 14556 8780 14608 8832
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 2504 8576 2556 8628
rect 2320 8440 2372 8492
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2320 8304 2372 8356
rect 2504 8236 2556 8288
rect 2688 8236 2740 8288
rect 3700 8508 3752 8560
rect 3240 8372 3292 8424
rect 4160 8576 4212 8628
rect 4712 8576 4764 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6184 8576 6236 8628
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 6920 8576 6972 8628
rect 8300 8576 8352 8628
rect 8392 8576 8444 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 5816 8508 5868 8560
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 3792 8304 3844 8356
rect 5356 8440 5408 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6092 8508 6144 8560
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 7840 8440 7892 8492
rect 9864 8576 9916 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 10968 8576 11020 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 12624 8576 12676 8628
rect 13360 8576 13412 8628
rect 14280 8619 14332 8628
rect 14280 8585 14289 8619
rect 14289 8585 14323 8619
rect 14323 8585 14332 8619
rect 14280 8576 14332 8585
rect 10048 8508 10100 8560
rect 3148 8236 3200 8288
rect 4896 8236 4948 8288
rect 9956 8372 10008 8424
rect 9864 8304 9916 8356
rect 12072 8440 12124 8492
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 13820 8508 13872 8560
rect 13728 8440 13780 8492
rect 11796 8304 11848 8356
rect 12256 8304 12308 8356
rect 12992 8372 13044 8424
rect 13268 8372 13320 8424
rect 8392 8236 8444 8288
rect 9128 8236 9180 8288
rect 13360 8236 13412 8288
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 13544 8236 13596 8245
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 2412 8032 2464 8084
rect 3884 8032 3936 8084
rect 5264 8032 5316 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 7380 7964 7432 8016
rect 2228 7828 2280 7880
rect 7012 7896 7064 7948
rect 12164 8032 12216 8084
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13544 8032 13596 8084
rect 14464 8032 14516 8084
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3700 7828 3752 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4896 7828 4948 7880
rect 3056 7760 3108 7812
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 6460 7828 6512 7880
rect 6552 7828 6604 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7656 7828 7708 7880
rect 7840 7828 7892 7880
rect 8208 7828 8260 7880
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 9128 7828 9180 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 11612 7828 11664 7880
rect 12164 7828 12216 7880
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13452 7828 13504 7880
rect 14096 7828 14148 7880
rect 12440 7760 12492 7812
rect 4896 7692 4948 7744
rect 7472 7692 7524 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 8944 7692 8996 7744
rect 9956 7692 10008 7744
rect 10876 7692 10928 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 14188 7760 14240 7812
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2320 7488 2372 7540
rect 2504 7488 2556 7540
rect 2228 7420 2280 7472
rect 3516 7488 3568 7540
rect 3884 7488 3936 7540
rect 4896 7488 4948 7540
rect 3792 7352 3844 7404
rect 4160 7352 4212 7404
rect 3240 7284 3292 7336
rect 5816 7352 5868 7404
rect 6828 7488 6880 7540
rect 7288 7488 7340 7540
rect 7472 7488 7524 7540
rect 6920 7352 6972 7404
rect 7196 7352 7248 7404
rect 8208 7420 8260 7472
rect 10876 7352 10928 7404
rect 11612 7352 11664 7404
rect 12164 7488 12216 7540
rect 12992 7488 13044 7540
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 14096 7488 14148 7540
rect 14188 7488 14240 7540
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 3148 7216 3200 7268
rect 5632 7216 5684 7268
rect 6460 7284 6512 7336
rect 12808 7284 12860 7336
rect 13176 7352 13228 7404
rect 11152 7216 11204 7268
rect 13176 7216 13228 7268
rect 14372 7284 14424 7336
rect 2412 7148 2464 7200
rect 4160 7148 4212 7200
rect 4252 7148 4304 7200
rect 6460 7148 6512 7200
rect 8300 7148 8352 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 13636 7148 13688 7200
rect 13728 7148 13780 7200
rect 14004 7148 14056 7200
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 3056 6987 3108 6996
rect 3056 6953 3065 6987
rect 3065 6953 3099 6987
rect 3099 6953 3108 6987
rect 3056 6944 3108 6953
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 5632 6944 5684 6996
rect 5908 6944 5960 6996
rect 7656 6944 7708 6996
rect 9956 6944 10008 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 3516 6876 3568 6928
rect 8484 6876 8536 6928
rect 940 6808 992 6860
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 2320 6808 2372 6860
rect 2504 6740 2556 6792
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 6460 6808 6512 6860
rect 6644 6808 6696 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 8300 6851 8352 6860
rect 8300 6817 8309 6851
rect 8309 6817 8343 6851
rect 8343 6817 8352 6851
rect 8300 6808 8352 6817
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 5908 6740 5960 6792
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 9864 6808 9916 6860
rect 10784 6876 10836 6928
rect 11060 6808 11112 6860
rect 8760 6740 8812 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10416 6740 10468 6792
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 10876 6740 10928 6792
rect 11796 6808 11848 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12624 6876 12676 6928
rect 11704 6740 11756 6792
rect 12440 6808 12492 6860
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 13268 6740 13320 6792
rect 14372 6740 14424 6792
rect 4988 6604 5040 6656
rect 5448 6604 5500 6656
rect 6828 6604 6880 6656
rect 7656 6604 7708 6656
rect 8392 6604 8444 6656
rect 10232 6604 10284 6656
rect 10324 6604 10376 6656
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 13820 6604 13872 6656
rect 13912 6604 13964 6656
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2504 6400 2556 6452
rect 3148 6400 3200 6452
rect 3700 6400 3752 6452
rect 5080 6400 5132 6452
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 2320 6332 2372 6384
rect 3240 6332 3292 6384
rect 1492 6264 1544 6273
rect 5816 6400 5868 6452
rect 6644 6400 6696 6452
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 2228 6196 2280 6205
rect 2412 6196 2464 6248
rect 5540 6264 5592 6316
rect 6460 6332 6512 6384
rect 10600 6332 10652 6384
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9220 6264 9272 6316
rect 11152 6332 11204 6384
rect 11244 6332 11296 6384
rect 11704 6332 11756 6384
rect 13452 6400 13504 6452
rect 11980 6332 12032 6384
rect 11612 6264 11664 6316
rect 12716 6332 12768 6384
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 1860 6060 1912 6112
rect 4988 6060 5040 6112
rect 6644 6128 6696 6180
rect 7196 6196 7248 6248
rect 8392 6196 8444 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 10968 6060 11020 6112
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 12164 6196 12216 6248
rect 13360 6196 13412 6248
rect 12624 6128 12676 6180
rect 11520 6060 11572 6112
rect 11612 6060 11664 6112
rect 12072 6060 12124 6112
rect 13820 6060 13872 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 1860 5856 1912 5908
rect 3240 5856 3292 5908
rect 3700 5856 3752 5908
rect 5264 5856 5316 5908
rect 5632 5856 5684 5908
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 6828 5856 6880 5908
rect 7288 5856 7340 5908
rect 1584 5720 1636 5772
rect 2872 5788 2924 5840
rect 3792 5788 3844 5840
rect 4160 5720 4212 5772
rect 5540 5720 5592 5772
rect 1492 5652 1544 5704
rect 2964 5652 3016 5704
rect 1308 5584 1360 5636
rect 5448 5584 5500 5636
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6460 5652 6512 5704
rect 7840 5831 7892 5840
rect 7840 5797 7849 5831
rect 7849 5797 7883 5831
rect 7883 5797 7892 5831
rect 7840 5788 7892 5797
rect 9128 5856 9180 5908
rect 9220 5856 9272 5908
rect 10508 5856 10560 5908
rect 6920 5720 6972 5772
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 8300 5720 8352 5772
rect 10140 5831 10192 5840
rect 10140 5797 10149 5831
rect 10149 5797 10183 5831
rect 10183 5797 10192 5831
rect 10140 5788 10192 5797
rect 7840 5652 7892 5704
rect 11520 5899 11572 5908
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 11704 5856 11756 5908
rect 13360 5899 13412 5908
rect 13360 5865 13369 5899
rect 13369 5865 13403 5899
rect 13403 5865 13412 5899
rect 13360 5856 13412 5865
rect 14280 5856 14332 5908
rect 12532 5831 12584 5840
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 12532 5788 12584 5797
rect 13268 5720 13320 5772
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 2412 5516 2464 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 9864 5652 9916 5704
rect 8668 5584 8720 5636
rect 9680 5584 9732 5636
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 11612 5652 11664 5704
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 8484 5516 8536 5568
rect 9588 5516 9640 5568
rect 9772 5516 9824 5568
rect 10876 5584 10928 5636
rect 11704 5584 11756 5636
rect 12440 5584 12492 5636
rect 10324 5516 10376 5568
rect 10968 5516 11020 5568
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13636 5652 13688 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 2964 5312 3016 5364
rect 2872 5244 2924 5296
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 2412 5176 2464 5228
rect 3240 5176 3292 5228
rect 3424 5176 3476 5228
rect 3516 5176 3568 5228
rect 4068 5312 4120 5364
rect 4804 5312 4856 5364
rect 5356 5312 5408 5364
rect 5448 5312 5500 5364
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4988 5244 5040 5296
rect 5172 5244 5224 5296
rect 5816 5312 5868 5364
rect 7656 5312 7708 5364
rect 8208 5312 8260 5364
rect 5908 5176 5960 5228
rect 6460 5176 6512 5228
rect 6644 5176 6696 5228
rect 940 5108 992 5160
rect 1768 4972 1820 5024
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 7196 5176 7248 5228
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7012 5108 7064 5160
rect 4620 4972 4672 5024
rect 4896 4972 4948 5024
rect 5356 4972 5408 5024
rect 5632 4972 5684 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 6644 4972 6696 5024
rect 6736 4972 6788 5024
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 9680 5312 9732 5364
rect 10692 5312 10744 5364
rect 12072 5312 12124 5364
rect 12532 5312 12584 5364
rect 8944 5244 8996 5296
rect 9312 5176 9364 5228
rect 9864 5108 9916 5160
rect 10140 5176 10192 5228
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13912 5176 13964 5228
rect 14832 5176 14884 5228
rect 11612 5108 11664 5160
rect 11980 5151 12032 5160
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 13360 5108 13412 5160
rect 9588 5040 9640 5092
rect 12716 5040 12768 5092
rect 14188 5083 14240 5092
rect 14188 5049 14197 5083
rect 14197 5049 14231 5083
rect 14231 5049 14240 5083
rect 14188 5040 14240 5049
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 11244 4972 11296 5024
rect 12072 4972 12124 5024
rect 12440 4972 12492 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 2228 4768 2280 4820
rect 3516 4768 3568 4820
rect 5724 4768 5776 4820
rect 6092 4768 6144 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 6920 4768 6972 4820
rect 7656 4768 7708 4820
rect 8484 4768 8536 4820
rect 8944 4768 8996 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9772 4768 9824 4820
rect 10508 4768 10560 4820
rect 11520 4768 11572 4820
rect 11612 4768 11664 4820
rect 3240 4743 3292 4752
rect 3240 4709 3249 4743
rect 3249 4709 3283 4743
rect 3283 4709 3292 4743
rect 3240 4700 3292 4709
rect 3424 4700 3476 4752
rect 3976 4700 4028 4752
rect 4712 4700 4764 4752
rect 2136 4675 2188 4684
rect 2136 4641 2145 4675
rect 2145 4641 2179 4675
rect 2179 4641 2188 4675
rect 2136 4632 2188 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3148 4632 3200 4684
rect 5356 4700 5408 4752
rect 1584 4564 1636 4616
rect 1860 4428 1912 4480
rect 3700 4564 3752 4616
rect 4620 4564 4672 4616
rect 4896 4564 4948 4616
rect 5908 4632 5960 4684
rect 6460 4632 6512 4684
rect 6828 4632 6880 4684
rect 4804 4539 4856 4548
rect 4804 4505 4813 4539
rect 4813 4505 4847 4539
rect 4847 4505 4856 4539
rect 4804 4496 4856 4505
rect 5908 4496 5960 4548
rect 8300 4700 8352 4752
rect 8300 4564 8352 4616
rect 8484 4564 8536 4616
rect 13544 4768 13596 4820
rect 9772 4632 9824 4684
rect 11244 4632 11296 4684
rect 12164 4632 12216 4684
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9588 4607 9640 4616
rect 9588 4573 9597 4607
rect 9597 4573 9631 4607
rect 9631 4573 9640 4607
rect 9588 4564 9640 4573
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11704 4564 11756 4616
rect 11888 4564 11940 4616
rect 4252 4428 4304 4480
rect 9956 4428 10008 4480
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 10968 4428 11020 4480
rect 12900 4428 12952 4480
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 3884 4224 3936 4276
rect 1492 4088 1544 4140
rect 2136 4088 2188 4140
rect 3424 4156 3476 4208
rect 4712 4156 4764 4208
rect 4804 4156 4856 4208
rect 940 4020 992 4072
rect 2136 3952 2188 4004
rect 3148 4088 3200 4140
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 5448 4088 5500 4140
rect 6092 4224 6144 4276
rect 7012 4224 7064 4276
rect 9220 4224 9272 4276
rect 12256 4224 12308 4276
rect 6644 4156 6696 4208
rect 3516 4020 3568 4072
rect 5264 4020 5316 4072
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 6000 4020 6052 4072
rect 6644 4020 6696 4072
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9588 4156 9640 4208
rect 9864 4088 9916 4140
rect 11704 4156 11756 4208
rect 10048 4088 10100 4140
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8208 4020 8260 4072
rect 9680 4020 9732 4072
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 10324 4020 10376 4072
rect 7196 3952 7248 4004
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 5724 3884 5776 3936
rect 7104 3884 7156 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 10416 3884 10468 3936
rect 12624 4131 12676 4140
rect 12624 4097 12642 4131
rect 12642 4097 12676 4131
rect 12624 4088 12676 4097
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 14096 4131 14148 4140
rect 14096 4097 14114 4131
rect 14114 4097 14148 4131
rect 14096 4088 14148 4097
rect 11152 3884 11204 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 2964 3680 3016 3732
rect 3148 3680 3200 3732
rect 6644 3680 6696 3732
rect 7840 3680 7892 3732
rect 8576 3680 8628 3732
rect 9312 3680 9364 3732
rect 9864 3680 9916 3732
rect 2044 3612 2096 3664
rect 2136 3655 2188 3664
rect 2136 3621 2145 3655
rect 2145 3621 2179 3655
rect 2179 3621 2188 3655
rect 2136 3612 2188 3621
rect 3700 3612 3752 3664
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 4436 3612 4488 3664
rect 5908 3612 5960 3664
rect 7656 3655 7708 3664
rect 7656 3621 7665 3655
rect 7665 3621 7699 3655
rect 7699 3621 7708 3655
rect 7656 3612 7708 3621
rect 1860 3476 1912 3528
rect 2136 3340 2188 3392
rect 2504 3451 2556 3460
rect 2504 3417 2538 3451
rect 2538 3417 2556 3451
rect 2504 3408 2556 3417
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 4160 3544 4212 3596
rect 5540 3544 5592 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 8852 3612 8904 3664
rect 10416 3612 10468 3664
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 12624 3680 12676 3732
rect 14096 3680 14148 3732
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 14280 3612 14332 3664
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 4712 3451 4764 3460
rect 4712 3417 4746 3451
rect 4746 3417 4764 3451
rect 4712 3408 4764 3417
rect 4896 3408 4948 3460
rect 4988 3408 5040 3460
rect 6368 3408 6420 3460
rect 3516 3340 3568 3392
rect 6644 3340 6696 3392
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 12808 3544 12860 3596
rect 12072 3476 12124 3528
rect 9404 3451 9456 3460
rect 9404 3417 9438 3451
rect 9438 3417 9456 3451
rect 9404 3408 9456 3417
rect 11152 3408 11204 3460
rect 11520 3408 11572 3460
rect 14188 3476 14240 3528
rect 14556 3476 14608 3528
rect 11612 3340 11664 3392
rect 11888 3340 11940 3392
rect 14188 3340 14240 3392
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 2688 3136 2740 3188
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 4160 3136 4212 3188
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 4068 3000 4120 3052
rect 4252 3068 4304 3120
rect 5540 3136 5592 3188
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 7196 3136 7248 3188
rect 7380 3136 7432 3188
rect 10600 3136 10652 3188
rect 11152 3136 11204 3188
rect 11612 3136 11664 3188
rect 5356 3068 5408 3120
rect 7012 3068 7064 3120
rect 3148 2796 3200 2848
rect 4252 2796 4304 2848
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 5908 3000 5960 3052
rect 8760 3068 8812 3120
rect 9220 3068 9272 3120
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 8484 3000 8536 3052
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 10968 3043 11020 3052
rect 10968 3009 10986 3043
rect 10986 3009 11020 3043
rect 10968 3000 11020 3009
rect 12808 3068 12860 3120
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 12164 2932 12216 2984
rect 6920 2796 6972 2848
rect 7196 2796 7248 2848
rect 8392 2796 8444 2848
rect 9956 2864 10008 2916
rect 13268 3068 13320 3120
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 9404 2796 9456 2848
rect 10876 2796 10928 2848
rect 14556 2796 14608 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 4712 2592 4764 2601
rect 5172 2592 5224 2644
rect 8208 2592 8260 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 2044 2567 2096 2576
rect 2044 2533 2053 2567
rect 2053 2533 2087 2567
rect 2087 2533 2096 2567
rect 2044 2524 2096 2533
rect 2412 2567 2464 2576
rect 2412 2533 2421 2567
rect 2421 2533 2455 2567
rect 2455 2533 2464 2567
rect 2412 2524 2464 2533
rect 4528 2524 4580 2576
rect 3240 2456 3292 2508
rect 572 2388 624 2440
rect 1308 2320 1360 2372
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 10048 2524 10100 2576
rect 10232 2524 10284 2576
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 12164 2592 12216 2644
rect 13360 2592 13412 2644
rect 14096 2592 14148 2644
rect 6644 2456 6696 2508
rect 6920 2456 6972 2508
rect 7656 2456 7708 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 4804 2388 4856 2440
rect 4988 2320 5040 2372
rect 3148 2252 3200 2304
rect 6460 2388 6512 2440
rect 7196 2388 7248 2440
rect 8208 2388 8260 2440
rect 8392 2388 8444 2440
rect 8760 2388 8812 2440
rect 11060 2388 11112 2440
rect 12440 2388 12492 2440
rect 14004 2388 14056 2440
rect 7288 2320 7340 2372
rect 8852 2252 8904 2304
rect 10416 2320 10468 2372
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 11612 2320 11664 2329
rect 12716 2363 12768 2372
rect 12716 2329 12725 2363
rect 12725 2329 12759 2363
rect 12759 2329 12768 2363
rect 12716 2320 12768 2329
rect 11888 2252 11940 2304
rect 12348 2252 12400 2304
rect 13084 2252 13136 2304
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 2320 2048 2372 2100
rect 6184 2048 6236 2100
rect 8208 2048 8260 2100
rect 14188 2048 14240 2100
rect 2780 1980 2832 2032
rect 5264 1980 5316 2032
<< metal2 >>
rect 938 23338 994 24000
rect 938 23310 1164 23338
rect 938 23200 994 23310
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 952 21049 980 21422
rect 938 21040 994 21049
rect 938 20975 994 20984
rect 940 20256 992 20262
rect 940 20198 992 20204
rect 952 19961 980 20198
rect 938 19952 994 19961
rect 938 19887 994 19896
rect 940 19168 992 19174
rect 940 19110 992 19116
rect 952 18873 980 19110
rect 938 18864 994 18873
rect 938 18799 994 18808
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 952 17678 980 17711
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 940 16992 992 16998
rect 940 16934 992 16940
rect 952 16697 980 16934
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15609 980 15846
rect 938 15600 994 15609
rect 938 15535 994 15544
rect 1136 14890 1164 23310
rect 1674 23202 1730 24000
rect 1780 23310 1992 23338
rect 1780 23202 1808 23310
rect 1674 23200 1808 23202
rect 1688 23174 1808 23200
rect 1490 22128 1546 22137
rect 1490 22063 1546 22072
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 20448 1440 21490
rect 1504 21146 1532 22063
rect 1584 21344 1636 21350
rect 1636 21304 1716 21332
rect 1584 21286 1636 21292
rect 1492 21140 1544 21146
rect 1492 21082 1544 21088
rect 1412 20420 1532 20448
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17338 1440 18226
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 16250 1440 16390
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1124 14884 1176 14890
rect 1124 14826 1176 14832
rect 938 14512 994 14521
rect 938 14447 994 14456
rect 952 14414 980 14447
rect 940 14408 992 14414
rect 940 14350 992 14356
rect 1412 14074 1440 15438
rect 1504 14618 1532 20420
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1596 18290 1624 19654
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 16658 1624 18022
rect 1688 17490 1716 21304
rect 1768 20868 1820 20874
rect 1768 20810 1820 20816
rect 1780 20777 1808 20810
rect 1860 20800 1912 20806
rect 1766 20768 1822 20777
rect 1860 20742 1912 20748
rect 1766 20703 1822 20712
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 17762 1808 19314
rect 1872 18766 1900 20742
rect 1964 19718 1992 23310
rect 2410 23200 2466 24000
rect 2778 23216 2834 23225
rect 2044 21616 2096 21622
rect 2044 21558 2096 21564
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1964 18970 1992 19314
rect 2056 18970 2084 21558
rect 2136 21548 2188 21554
rect 2136 21490 2188 21496
rect 2148 20777 2176 21490
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2134 20768 2190 20777
rect 2134 20703 2190 20712
rect 2240 20602 2268 20878
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2240 19786 2268 20402
rect 2228 19780 2280 19786
rect 2228 19722 2280 19728
rect 2240 19242 2268 19722
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 2148 18290 2176 19110
rect 2240 18766 2268 19178
rect 2332 18834 2360 20742
rect 2424 20602 2452 23200
rect 3146 23200 3202 24000
rect 3882 23200 3938 24000
rect 4264 23310 4568 23338
rect 2778 23151 2834 23160
rect 2792 21690 2820 23151
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3068 21690 3096 21830
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 2663 21244 2971 21253
rect 2663 21242 2669 21244
rect 2725 21242 2749 21244
rect 2805 21242 2829 21244
rect 2885 21242 2909 21244
rect 2965 21242 2971 21244
rect 2725 21190 2727 21242
rect 2907 21190 2909 21242
rect 2663 21188 2669 21190
rect 2725 21188 2749 21190
rect 2805 21188 2829 21190
rect 2885 21188 2909 21190
rect 2965 21188 2971 21190
rect 2663 21179 2971 21188
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2884 20466 2912 20878
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2516 19417 2544 20402
rect 2663 20156 2971 20165
rect 2663 20154 2669 20156
rect 2725 20154 2749 20156
rect 2805 20154 2829 20156
rect 2885 20154 2909 20156
rect 2965 20154 2971 20156
rect 2725 20102 2727 20154
rect 2907 20102 2909 20154
rect 2663 20100 2669 20102
rect 2725 20100 2749 20102
rect 2805 20100 2829 20102
rect 2885 20100 2909 20102
rect 2965 20100 2971 20102
rect 2663 20091 2971 20100
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2792 19446 2820 19722
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2780 19440 2832 19446
rect 2502 19408 2558 19417
rect 2780 19382 2832 19388
rect 2502 19343 2558 19352
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18426 2360 18566
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 1780 17734 1992 17762
rect 1766 17640 1822 17649
rect 1766 17575 1768 17584
rect 1820 17575 1822 17584
rect 1768 17546 1820 17552
rect 1688 17462 1900 17490
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16946 1808 17138
rect 1688 16918 1808 16946
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15026 1624 15302
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13258 1624 13806
rect 1688 13258 1716 16918
rect 1872 16574 1900 17462
rect 1964 16776 1992 17734
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 1964 16748 2084 16776
rect 1872 16546 1992 16574
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1584 13252 1636 13258
rect 1584 13194 1636 13200
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1596 12850 1624 13194
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 938 12336 994 12345
rect 938 12271 994 12280
rect 952 12238 980 12271
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 10169 1348 10542
rect 1306 10160 1362 10169
rect 1306 10095 1362 10104
rect 1412 10062 1440 11047
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 940 9512 992 9518
rect 940 9454 992 9460
rect 952 9081 980 9454
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 8106 1532 12038
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10266 1624 10610
rect 1780 10554 1808 16050
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 12986 1900 13806
rect 1964 13462 1992 16546
rect 2056 15162 2084 16748
rect 2148 15434 2176 17138
rect 2240 17082 2268 18158
rect 2424 18086 2452 19246
rect 2663 19068 2971 19077
rect 2663 19066 2669 19068
rect 2725 19066 2749 19068
rect 2805 19066 2829 19068
rect 2885 19066 2909 19068
rect 2965 19066 2971 19068
rect 2725 19014 2727 19066
rect 2907 19014 2909 19066
rect 2663 19012 2669 19014
rect 2725 19012 2749 19014
rect 2805 19012 2829 19014
rect 2885 19012 2909 19014
rect 2965 19012 2971 19014
rect 2663 19003 2971 19012
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2424 17882 2452 18022
rect 2663 17980 2971 17989
rect 2663 17978 2669 17980
rect 2725 17978 2749 17980
rect 2805 17978 2829 17980
rect 2885 17978 2909 17980
rect 2965 17978 2971 17980
rect 2725 17926 2727 17978
rect 2907 17926 2909 17978
rect 2663 17924 2669 17926
rect 2725 17924 2749 17926
rect 2805 17924 2829 17926
rect 2885 17924 2909 17926
rect 2965 17924 2971 17926
rect 2663 17915 2971 17924
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2240 17054 2360 17082
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 15570 2268 16934
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13530 2084 13806
rect 2240 13530 2268 15030
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1872 12306 1900 12922
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11762 1900 12242
rect 1964 12238 1992 13262
rect 2332 12986 2360 17054
rect 2424 16674 2452 17138
rect 2884 17082 2912 17614
rect 2964 17536 3016 17542
rect 3068 17524 3096 19654
rect 3160 17626 3188 23200
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 21554 3832 21966
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3332 20800 3384 20806
rect 3436 20777 3464 21286
rect 3620 21010 3648 21490
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3332 20742 3384 20748
rect 3422 20768 3478 20777
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3252 18222 3280 19858
rect 3344 19446 3372 20742
rect 3422 20703 3478 20712
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3436 18834 3464 20538
rect 3528 19854 3556 20946
rect 3896 20058 3924 23200
rect 4264 22094 4292 23310
rect 4540 23202 4568 23310
rect 4618 23202 4674 24000
rect 4540 23200 4674 23202
rect 5354 23200 5410 24000
rect 6090 23200 6146 24000
rect 6826 23200 6882 24000
rect 7562 23338 7618 24000
rect 7562 23310 7696 23338
rect 7562 23200 7618 23310
rect 4540 23174 4660 23200
rect 5368 22094 5396 23200
rect 4080 22066 4292 22094
rect 5276 22066 5396 22094
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3988 21350 4016 21898
rect 4080 21622 4108 22066
rect 5276 22030 5304 22066
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4376 21788 4684 21797
rect 4376 21786 4382 21788
rect 4438 21786 4462 21788
rect 4518 21786 4542 21788
rect 4598 21786 4622 21788
rect 4678 21786 4684 21788
rect 4438 21734 4440 21786
rect 4620 21734 4622 21786
rect 4376 21732 4382 21734
rect 4438 21732 4462 21734
rect 4518 21732 4542 21734
rect 4598 21732 4622 21734
rect 4678 21732 4684 21734
rect 4376 21723 4684 21732
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 4068 21616 4120 21622
rect 5264 21616 5316 21622
rect 4068 21558 4120 21564
rect 4816 21554 5120 21570
rect 5264 21558 5316 21564
rect 4804 21548 5120 21554
rect 4856 21542 5120 21548
rect 4804 21490 4856 21496
rect 4252 21480 4304 21486
rect 4252 21422 4304 21428
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 4264 21146 4292 21422
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20602 4016 20878
rect 4376 20700 4684 20709
rect 4376 20698 4382 20700
rect 4438 20698 4462 20700
rect 4518 20698 4542 20700
rect 4598 20698 4622 20700
rect 4678 20698 4684 20700
rect 4438 20646 4440 20698
rect 4620 20646 4622 20698
rect 4376 20644 4382 20646
rect 4438 20644 4462 20646
rect 4518 20644 4542 20646
rect 4598 20644 4622 20646
rect 4678 20644 4684 20646
rect 4376 20635 4684 20644
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4724 20346 4752 21286
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 20534 4844 20742
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 4080 19922 4108 20334
rect 4724 20318 4844 20346
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18970 3556 19246
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3620 18426 3648 19178
rect 3896 18766 3924 19790
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 4080 19514 4108 19722
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3252 17746 3280 18022
rect 3344 17882 3372 18022
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3424 17672 3476 17678
rect 3160 17598 3372 17626
rect 3424 17614 3476 17620
rect 3068 17496 3280 17524
rect 2964 17478 3016 17484
rect 2976 17202 3004 17478
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2884 17054 3096 17082
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 3068 16674 3096 17054
rect 3148 16720 3200 16726
rect 2424 16646 2820 16674
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15094 2452 15846
rect 2516 15706 2544 16458
rect 2792 16250 2820 16646
rect 2976 16668 3148 16674
rect 2976 16662 3200 16668
rect 2976 16646 3188 16662
rect 2976 16590 3004 16646
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2976 16046 3004 16390
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2516 14822 2544 15438
rect 3068 15026 3096 15846
rect 3160 15706 3188 15914
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3252 15026 3280 17496
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14408 2464 14414
rect 2410 14376 2412 14385
rect 2464 14376 2466 14385
rect 2410 14311 2466 14320
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 13394 2452 14214
rect 2516 14074 2544 14758
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2608 13682 2636 14350
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 14074 2912 14214
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2516 13654 2636 13682
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2148 12442 2176 12786
rect 2424 12730 2452 12854
rect 2516 12782 2544 13654
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 3056 13320 3108 13326
rect 3108 13280 3188 13308
rect 3056 13262 3108 13268
rect 2332 12702 2452 12730
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11354 1900 11494
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1964 11150 1992 12174
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1688 10526 1808 10554
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1688 8786 1716 10526
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 8974 1808 10406
rect 1872 10062 1900 11018
rect 1964 10606 1992 11086
rect 2056 10810 2084 12106
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11354 2268 11630
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10606 2176 10950
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2240 10418 2268 11018
rect 2056 10390 2268 10418
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9586 1900 9998
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1688 8758 1808 8786
rect 1412 8078 1532 8106
rect 938 6896 994 6905
rect 938 6831 940 6840
rect 992 6831 994 6840
rect 940 6802 992 6808
rect 1306 5808 1362 5817
rect 1306 5743 1362 5752
rect 1320 5642 1348 5743
rect 1308 5636 1360 5642
rect 1308 5578 1360 5584
rect 1412 5522 1440 8078
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1504 5710 1532 6258
rect 1596 5778 1624 7686
rect 1674 6896 1730 6905
rect 1674 6831 1676 6840
rect 1728 6831 1730 6840
rect 1676 6802 1728 6808
rect 1674 6216 1730 6225
rect 1674 6151 1730 6160
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1584 5568 1636 5574
rect 1412 5494 1532 5522
rect 1584 5510 1636 5516
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1504 4146 1532 5494
rect 1596 4622 1624 5510
rect 1688 5234 1716 6151
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1780 5030 1808 8758
rect 1950 7848 2006 7857
rect 1950 7783 2006 7792
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5914 1900 6054
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 952 3641 980 4014
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 1872 3534 1900 4422
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1674 3088 1730 3097
rect 1674 3023 1676 3032
rect 1728 3023 1730 3032
rect 1676 2994 1728 3000
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2689 1440 2926
rect 1398 2680 1454 2689
rect 1398 2615 1454 2624
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 584 800 612 2382
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 1320 800 1348 2314
rect 1688 1873 1716 2314
rect 1674 1864 1730 1873
rect 1674 1799 1730 1808
rect 1964 1465 1992 7783
rect 2056 4570 2084 10390
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2148 8838 2176 9454
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 4690 2176 8774
rect 2240 7886 2268 9998
rect 2332 8498 2360 12702
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 3068 12434 3096 12718
rect 2976 12406 3096 12434
rect 3160 12434 3188 13280
rect 3252 12986 3280 14826
rect 3344 14482 3372 17598
rect 3436 17338 3464 17614
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15434 3464 16050
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 12986 3372 14214
rect 3528 13530 3556 18226
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17241 3648 17478
rect 3606 17232 3662 17241
rect 3606 17167 3662 17176
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3712 16590 3740 16730
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15706 3648 15914
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15706 3740 15846
rect 3804 15706 3832 18702
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3896 17542 3924 17818
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3896 16794 3924 17478
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3896 16250 3924 16526
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3620 15162 3648 15642
rect 3988 15502 4016 19450
rect 4172 18970 4200 19790
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4264 19292 4292 19722
rect 4376 19612 4684 19621
rect 4376 19610 4382 19612
rect 4438 19610 4462 19612
rect 4518 19610 4542 19612
rect 4598 19610 4622 19612
rect 4678 19610 4684 19612
rect 4438 19558 4440 19610
rect 4620 19558 4622 19610
rect 4376 19556 4382 19558
rect 4438 19556 4462 19558
rect 4518 19556 4542 19558
rect 4598 19556 4622 19558
rect 4678 19556 4684 19558
rect 4376 19547 4684 19556
rect 4724 19378 4752 19926
rect 4816 19786 4844 20318
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4908 19514 4936 19722
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 5000 19394 5028 21286
rect 5092 19496 5120 21542
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 20788 5212 21490
rect 5276 21010 5304 21558
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5264 20800 5316 20806
rect 5184 20760 5264 20788
rect 5368 20777 5396 21286
rect 5460 21010 5488 21286
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5552 20856 5580 21626
rect 5828 20942 5856 21626
rect 6104 21486 6132 23200
rect 6840 21622 6868 23200
rect 7668 21690 7696 23310
rect 8298 23200 8354 24000
rect 9034 23200 9090 24000
rect 9770 23200 9826 24000
rect 10506 23338 10562 24000
rect 10506 23310 10824 23338
rect 10506 23200 10562 23310
rect 8312 22094 8340 23200
rect 8312 22066 8524 22094
rect 7803 21788 8111 21797
rect 7803 21786 7809 21788
rect 7865 21786 7889 21788
rect 7945 21786 7969 21788
rect 8025 21786 8049 21788
rect 8105 21786 8111 21788
rect 7865 21734 7867 21786
rect 8047 21734 8049 21786
rect 7803 21732 7809 21734
rect 7865 21732 7889 21734
rect 7945 21732 7969 21734
rect 8025 21732 8049 21734
rect 8105 21732 8111 21734
rect 7803 21723 8111 21732
rect 8496 21690 8524 22066
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8588 21690 8616 21830
rect 9048 21690 9076 23200
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6090 21244 6398 21253
rect 6090 21242 6096 21244
rect 6152 21242 6176 21244
rect 6232 21242 6256 21244
rect 6312 21242 6336 21244
rect 6392 21242 6398 21244
rect 6152 21190 6154 21242
rect 6334 21190 6336 21242
rect 6090 21188 6096 21190
rect 6152 21188 6176 21190
rect 6232 21188 6256 21190
rect 6312 21188 6336 21190
rect 6392 21188 6398 21190
rect 6090 21179 6398 21188
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5724 20868 5776 20874
rect 5552 20828 5672 20856
rect 5448 20800 5500 20806
rect 5264 20742 5316 20748
rect 5354 20768 5410 20777
rect 5092 19468 5212 19496
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4816 19366 5028 19394
rect 4344 19304 4396 19310
rect 4264 19264 4344 19292
rect 4816 19258 4844 19366
rect 5184 19334 5212 19468
rect 4344 19246 4396 19252
rect 4724 19230 4844 19258
rect 4896 19304 4948 19310
rect 5092 19306 5212 19334
rect 4948 19264 5028 19292
rect 4896 19246 4948 19252
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4436 18964 4488 18970
rect 4436 18906 4488 18912
rect 4448 18873 4476 18906
rect 4434 18864 4490 18873
rect 4434 18799 4490 18808
rect 4724 18737 4752 19230
rect 4710 18728 4766 18737
rect 4710 18663 4766 18672
rect 4376 18524 4684 18533
rect 4376 18522 4382 18524
rect 4438 18522 4462 18524
rect 4518 18522 4542 18524
rect 4598 18522 4622 18524
rect 4678 18522 4684 18524
rect 4438 18470 4440 18522
rect 4620 18470 4622 18522
rect 4376 18468 4382 18470
rect 4438 18468 4462 18470
rect 4518 18468 4542 18470
rect 4598 18468 4622 18470
rect 4678 18468 4684 18470
rect 4376 18459 4684 18468
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4080 17864 4108 18022
rect 4080 17836 4200 17864
rect 4172 17678 4200 17836
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4172 17134 4200 17614
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4264 17338 4292 17478
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16726 4200 17070
rect 4816 16998 4844 17614
rect 4908 17338 4936 18226
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 5000 17218 5028 19264
rect 4908 17190 5028 17218
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3804 15026 3832 15370
rect 4080 15314 4108 16662
rect 3896 15286 4108 15314
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3804 14414 3832 14962
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3528 12434 3556 13262
rect 3620 12782 3648 14214
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3160 12406 3280 12434
rect 2976 12306 3004 12406
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11082 2452 11494
rect 2516 11218 2544 12038
rect 3160 11898 3188 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2976 11762 3004 11834
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2516 10810 2544 11154
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10810 3188 11086
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 8634 2544 9930
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 3068 9110 3096 10542
rect 3252 9874 3280 12406
rect 3344 12406 3556 12434
rect 3344 11762 3372 12406
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3712 11558 3740 12038
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3160 9846 3280 9874
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7478 2268 7822
rect 2332 7546 2360 8298
rect 2424 8090 2452 8434
rect 2700 8294 2728 8842
rect 3160 8294 3188 9846
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3252 9178 3280 9658
rect 3344 9450 3372 10202
rect 3422 9616 3478 9625
rect 3422 9551 3478 9560
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3436 9178 3464 9551
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8430 3280 8910
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2516 7546 2544 8230
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 3160 7886 3188 8230
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2332 6866 2360 7482
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 6390 2360 6802
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2424 6338 2452 7142
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 3068 7002 3096 7754
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6458 2544 6734
rect 3160 6458 3188 7210
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3252 6390 3280 7278
rect 3240 6384 3292 6390
rect 2424 6310 2544 6338
rect 3240 6326 3292 6332
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2240 4826 2268 6190
rect 2318 5808 2374 5817
rect 2318 5743 2374 5752
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2332 4690 2360 5743
rect 2424 5574 2452 6190
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5370 2452 5510
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2056 4542 2176 4570
rect 2042 4176 2098 4185
rect 2148 4146 2176 4542
rect 2042 4111 2098 4120
rect 2136 4140 2188 4146
rect 2056 3670 2084 4111
rect 2136 4082 2188 4088
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 2148 3670 2176 3946
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 2136 3664 2188 3670
rect 2136 3606 2188 3612
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 2774 2176 3334
rect 2148 2746 2360 2774
rect 2044 2576 2096 2582
rect 2042 2544 2044 2553
rect 2096 2544 2098 2553
rect 2042 2479 2098 2488
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 1950 1456 2006 1465
rect 1950 1391 2006 1400
rect 2240 1170 2268 2314
rect 2332 2106 2360 2746
rect 2424 2582 2452 5170
rect 2516 3466 2544 6310
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 3252 5914 3280 6326
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 2872 5840 2924 5846
rect 3344 5794 3372 9046
rect 3528 8922 3556 10406
rect 3620 10266 3648 10610
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 2872 5782 2924 5788
rect 2884 5302 2912 5782
rect 3160 5766 3372 5794
rect 3436 8894 3556 8922
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2976 5370 3004 5646
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 3160 4690 3188 5766
rect 3436 5658 3464 8894
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 7546 3556 8774
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3252 5630 3464 5658
rect 3252 5234 3280 5630
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 5234 3464 5510
rect 3528 5234 3556 6870
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3422 5128 3478 5137
rect 3422 5063 3478 5072
rect 3436 5030 3464 5063
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3252 4146 3280 4694
rect 3436 4214 3464 4694
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 3160 3738 3188 4082
rect 3528 4078 3556 4762
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2964 3732 3016 3738
rect 3148 3732 3200 3738
rect 3016 3692 3096 3720
rect 2964 3674 3016 3680
rect 2778 3632 2834 3641
rect 2700 3590 2778 3618
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2700 3194 2728 3590
rect 3068 3618 3096 3692
rect 3148 3674 3200 3680
rect 3068 3590 3280 3618
rect 2778 3567 2834 3576
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 2792 3194 2820 3431
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 3160 2310 3188 2790
rect 3252 2514 3280 3590
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3097 3556 3334
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3620 2774 3648 8910
rect 3712 8566 3740 11494
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9722 3832 9998
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3896 9586 3924 15286
rect 4172 14006 4200 16662
rect 4816 16590 4844 16934
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4264 15706 4292 16526
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4724 16250 4752 16390
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15450 4384 16118
rect 4816 15706 4844 16118
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4264 15422 4384 15450
rect 4264 14906 4292 15422
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4908 15162 4936 17190
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 16250 5028 16390
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4264 14878 4384 14906
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14618 4292 14758
rect 4356 14618 4384 14878
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4540 14346 4568 14962
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 4264 13530 4292 14282
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4724 13938 4752 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14074 4844 14214
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4908 13802 4936 14554
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 5092 13682 5120 19306
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5184 15706 5212 16390
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5276 15094 5304 20742
rect 5500 20760 5580 20788
rect 5448 20742 5500 20748
rect 5354 20703 5410 20712
rect 5552 20602 5580 20760
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5644 20398 5672 20828
rect 5724 20810 5776 20816
rect 5736 20777 5764 20810
rect 5722 20768 5778 20777
rect 5722 20703 5778 20712
rect 5828 20482 5856 20878
rect 5736 20454 5856 20482
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5644 18834 5672 20334
rect 5736 20262 5764 20454
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 19378 5764 20198
rect 5920 19854 5948 21082
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 20602 6224 20878
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6184 20596 6236 20602
rect 6012 20556 6184 20584
rect 6012 20058 6040 20556
rect 6184 20538 6236 20544
rect 6472 20534 6500 20742
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6090 20156 6398 20165
rect 6090 20154 6096 20156
rect 6152 20154 6176 20156
rect 6232 20154 6256 20156
rect 6312 20154 6336 20156
rect 6392 20154 6398 20156
rect 6152 20102 6154 20154
rect 6334 20102 6336 20154
rect 6090 20100 6096 20102
rect 6152 20100 6176 20102
rect 6232 20100 6256 20102
rect 6312 20100 6336 20102
rect 6392 20100 6398 20102
rect 6090 20091 6398 20100
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6564 19922 6592 20198
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19514 6132 19790
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5552 18290 5580 18634
rect 5540 18284 5592 18290
rect 5592 18244 5672 18272
rect 5540 18226 5592 18232
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17610 5580 18022
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5644 17066 5672 18244
rect 5920 18154 5948 19110
rect 6090 19068 6398 19077
rect 6090 19066 6096 19068
rect 6152 19066 6176 19068
rect 6232 19066 6256 19068
rect 6312 19066 6336 19068
rect 6392 19066 6398 19068
rect 6152 19014 6154 19066
rect 6334 19014 6336 19066
rect 6090 19012 6096 19014
rect 6152 19012 6176 19014
rect 6232 19012 6256 19014
rect 6312 19012 6336 19014
rect 6392 19012 6398 19014
rect 6090 19003 6398 19012
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6012 18222 6040 18566
rect 6288 18358 6316 18634
rect 6472 18358 6500 19722
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6564 18714 6592 19246
rect 6656 18834 6684 19994
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6564 18686 6684 18714
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6472 18222 6500 18294
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 6090 17980 6398 17989
rect 6090 17978 6096 17980
rect 6152 17978 6176 17980
rect 6232 17978 6256 17980
rect 6312 17978 6336 17980
rect 6392 17978 6398 17980
rect 6152 17926 6154 17978
rect 6334 17926 6336 17978
rect 6090 17924 6096 17926
rect 6152 17924 6176 17926
rect 6232 17924 6256 17926
rect 6312 17924 6336 17926
rect 6392 17924 6398 17926
rect 6090 17915 6398 17924
rect 6564 17338 6592 18294
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5630 16688 5686 16697
rect 5630 16623 5632 16632
rect 5684 16623 5686 16632
rect 5632 16594 5684 16600
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16182 5764 16390
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14074 5580 14350
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 4908 13654 5120 13682
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4068 13456 4120 13462
rect 4066 13424 4068 13433
rect 4120 13424 4122 13433
rect 4066 13359 4122 13368
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12986 4016 13262
rect 4264 12986 4292 13466
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4724 12889 4752 13126
rect 4710 12880 4766 12889
rect 4528 12844 4580 12850
rect 4710 12815 4766 12824
rect 4528 12786 4580 12792
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4068 12640 4120 12646
rect 4066 12608 4068 12617
rect 4120 12608 4122 12617
rect 4066 12543 4122 12552
rect 4448 12374 4476 12718
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4540 12170 4568 12786
rect 4816 12764 4844 13262
rect 4724 12736 4844 12764
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4632 12374 4660 12582
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4724 11558 4752 12736
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10606 4016 10950
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4528 10668 4580 10674
rect 4724 10656 4752 11494
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4580 10628 4752 10656
rect 4528 10610 4580 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10266 4016 10542
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4080 10282 4108 10406
rect 3976 10260 4028 10266
rect 4080 10254 4200 10282
rect 3976 10202 4028 10208
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9722 4016 9998
rect 3976 9716 4028 9722
rect 4080 9697 4108 10134
rect 3976 9658 4028 9664
rect 4066 9688 4122 9697
rect 4066 9623 4122 9632
rect 4172 9602 4200 10254
rect 4264 9674 4292 10406
rect 4356 9926 4384 10610
rect 4540 10470 4568 10610
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4264 9646 4476 9674
rect 3884 9580 3936 9586
rect 4172 9574 4384 9602
rect 3884 9522 3936 9528
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 3804 9178 3924 9194
rect 3804 9172 3936 9178
rect 3804 9166 3884 9172
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3804 8362 3832 9166
rect 3884 9114 3936 9120
rect 3976 8968 4028 8974
rect 3974 8936 3976 8945
rect 4028 8936 4030 8945
rect 3974 8871 4030 8880
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 8356 3844 8362
rect 3712 8316 3792 8344
rect 3712 7886 3740 8316
rect 3792 8298 3844 8304
rect 3790 8256 3846 8265
rect 3790 8191 3846 8200
rect 3804 7886 3832 8191
rect 3896 8090 3924 8366
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3712 6458 3740 7822
rect 3804 7410 3832 7822
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3896 7290 3924 7482
rect 3804 7262 3924 7290
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3712 5914 3740 6394
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3804 5846 3832 7262
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 3670 3740 4558
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3804 3534 3832 4655
rect 3896 4282 3924 5170
rect 3988 4758 4016 8774
rect 4080 5370 4108 9415
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 9042 4200 9318
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4356 8906 4384 9574
rect 4448 9353 4476 9646
rect 4434 9344 4490 9353
rect 4434 9279 4490 9288
rect 4724 9178 4752 9998
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8974 4844 11222
rect 4908 8974 4936 13654
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 5000 12238 5028 13398
rect 5552 13190 5580 14010
rect 5736 13734 5764 14214
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12306 5212 12582
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11218 5028 12174
rect 5276 12170 5304 13126
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5368 12170 5396 12310
rect 5552 12306 5580 13126
rect 5736 12850 5764 13670
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5644 12374 5672 12786
rect 5828 12434 5856 17138
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6000 16448 6052 16454
rect 6380 16436 6408 16526
rect 6656 16522 6684 18686
rect 6748 16590 6776 19654
rect 6932 19514 6960 21558
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 7024 20806 7052 21490
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7116 20942 7144 21286
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7024 19514 7052 19722
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6840 17134 6868 18022
rect 7116 17678 7144 20878
rect 7208 20466 7236 21286
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7300 18816 7328 21490
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7932 21412 7984 21418
rect 7932 21354 7984 21360
rect 7392 20942 7420 21354
rect 7944 21146 7972 21354
rect 8496 21146 8524 21490
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 19378 7420 20198
rect 7484 19378 7512 20266
rect 7668 19938 7696 20742
rect 7803 20700 8111 20709
rect 7803 20698 7809 20700
rect 7865 20698 7889 20700
rect 7945 20698 7969 20700
rect 8025 20698 8049 20700
rect 8105 20698 8111 20700
rect 7865 20646 7867 20698
rect 8047 20646 8049 20698
rect 7803 20644 7809 20646
rect 7865 20644 7889 20646
rect 7945 20644 7969 20646
rect 8025 20644 8049 20646
rect 8105 20644 8111 20646
rect 7803 20635 8111 20644
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8128 20058 8156 20334
rect 8220 20262 8248 20878
rect 8312 20777 8340 20878
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8298 20768 8354 20777
rect 8298 20703 8354 20712
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8220 19990 8248 20198
rect 8208 19984 8260 19990
rect 7668 19910 8156 19938
rect 8208 19926 8260 19932
rect 8128 19802 8156 19910
rect 8392 19848 8444 19854
rect 7656 19780 7708 19786
rect 8128 19774 8248 19802
rect 8392 19790 8444 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 7656 19722 7708 19728
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7576 19310 7604 19654
rect 7668 19514 7696 19722
rect 7803 19612 8111 19621
rect 7803 19610 7809 19612
rect 7865 19610 7889 19612
rect 7945 19610 7969 19612
rect 8025 19610 8049 19612
rect 8105 19610 8111 19612
rect 7865 19558 7867 19610
rect 8047 19558 8049 19610
rect 7803 19556 7809 19558
rect 7865 19556 7889 19558
rect 7945 19556 7969 19558
rect 8025 19556 8049 19558
rect 8105 19556 8111 19558
rect 7803 19547 8111 19556
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7300 18788 7420 18816
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18358 7236 18566
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7300 18154 7328 18634
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6932 17338 6960 17614
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6920 16992 6972 16998
rect 7024 16980 7052 17478
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 6972 16952 7052 16980
rect 6920 16934 6972 16940
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6052 16408 6408 16436
rect 6000 16390 6052 16396
rect 6012 15638 6040 16390
rect 6748 16250 6776 16526
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 6656 15706 6684 15982
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6932 14958 6960 16934
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15706 7052 15846
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7116 15450 7144 17206
rect 7208 16998 7236 17478
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7024 15422 7144 15450
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6644 14816 6696 14822
rect 6564 14776 6644 14804
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6472 12434 6500 13874
rect 5828 12406 6224 12434
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11898 5120 12038
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5092 11082 5120 11562
rect 5920 11558 5948 12174
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 9625 5120 11018
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9178 5028 9318
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5092 9058 5120 9454
rect 5000 9030 5120 9058
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8634 4200 8774
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4724 8634 4752 8910
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4172 7410 4200 8570
rect 4436 7812 4488 7818
rect 4264 7772 4436 7800
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4264 7206 4292 7772
rect 4436 7754 4488 7760
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4172 5778 4200 7142
rect 4264 7002 4292 7142
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4250 6352 4306 6361
rect 4250 6287 4306 6296
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5364 4120 5370
rect 4264 5352 4292 6287
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4816 5370 4844 8910
rect 5000 8906 5028 9030
rect 5184 8922 5212 9862
rect 5276 9382 5304 10406
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5276 8974 5304 9046
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5092 8894 5212 8922
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5000 8430 5028 8842
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7886 4936 8230
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7546 4936 7686
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5092 6882 5120 8894
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4908 6854 5120 6882
rect 4068 5306 4120 5312
rect 4172 5324 4292 5352
rect 4804 5364 4856 5370
rect 4172 5250 4200 5324
rect 4804 5306 4856 5312
rect 4080 5222 4200 5250
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 4080 4570 4108 5222
rect 4908 5030 4936 6854
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 6118 5028 6598
rect 5092 6458 5120 6734
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5184 6338 5212 8774
rect 5276 8090 5304 8910
rect 5368 8498 5396 10474
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10266 5488 10406
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5276 6866 5304 8026
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5354 6760 5410 6769
rect 5354 6695 5410 6704
rect 5092 6310 5212 6338
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4988 5296 5040 5302
rect 4986 5264 4988 5273
rect 5040 5264 5042 5273
rect 4986 5199 5042 5208
rect 4620 5024 4672 5030
rect 4250 4992 4306 5001
rect 3988 4542 4108 4570
rect 4172 4950 4250 4978
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 3670 4016 4542
rect 4172 4146 4200 4950
rect 4620 4966 4672 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4250 4927 4306 4936
rect 4632 4622 4660 4966
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4080 3058 4108 3975
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3194 4200 3538
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4264 3126 4292 4422
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4724 4214 4752 4694
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4214 4844 4490
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4436 3664 4488 3670
rect 4488 3612 4844 3618
rect 4436 3606 4844 3612
rect 4448 3590 4844 3606
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 3528 2746 3648 2774
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2780 2032 2832 2038
rect 2780 1974 2832 1980
rect 2056 1142 2268 1170
rect 2056 800 2084 1142
rect 2792 800 2820 1974
rect 3528 800 3556 2746
rect 4264 800 4292 2790
rect 4724 2650 4752 3402
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4540 2394 4568 2518
rect 4816 2446 4844 3590
rect 4908 3466 4936 4558
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 5000 3058 5028 3402
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5092 2774 5120 6310
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5184 4593 5212 5238
rect 5170 4584 5226 4593
rect 5170 4519 5226 4528
rect 5276 4162 5304 5850
rect 5368 5370 5396 6695
rect 5460 6662 5488 9522
rect 5552 8090 5580 11086
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10810 5764 11018
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5644 9518 5672 9998
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9178 5672 9454
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5736 8634 5764 9590
rect 5920 9586 5948 10610
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8566 5856 9318
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5552 6322 5580 8026
rect 5644 7274 5672 8366
rect 5828 7410 5856 8502
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5816 7404 5868 7410
rect 5736 7364 5816 7392
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5778 5580 6258
rect 5644 5914 5672 6938
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5460 5370 5488 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4758 5396 4966
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5276 4134 5396 4162
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 2990 5212 3878
rect 5276 3641 5304 4014
rect 5262 3632 5318 3641
rect 5262 3567 5318 3576
rect 5368 3210 5396 4134
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5276 3182 5396 3210
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4908 2746 5120 2774
rect 4804 2440 4856 2446
rect 4540 2366 4752 2394
rect 4804 2382 4856 2388
rect 4724 2258 4752 2366
rect 4908 2258 4936 2746
rect 5184 2650 5212 2926
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4724 2230 4936 2258
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 5000 800 5028 2314
rect 5276 2038 5304 3182
rect 5356 3120 5408 3126
rect 5354 3088 5356 3097
rect 5408 3088 5410 3097
rect 5354 3023 5410 3032
rect 5460 2990 5488 4082
rect 5552 3602 5580 5714
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5030 5672 5646
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4706 5672 4966
rect 5736 4826 5764 7364
rect 5816 7346 5868 7352
rect 5920 7002 5948 8434
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5828 6458 5856 6734
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5828 5370 5856 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5920 5234 5948 6734
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6012 5080 6040 12106
rect 6104 11762 6132 12242
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6196 11540 6224 12406
rect 6288 12406 6500 12434
rect 6288 11762 6316 12406
rect 6460 12232 6512 12238
rect 6564 12220 6592 14776
rect 6644 14758 6696 14764
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6748 13530 6776 13806
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6512 12192 6592 12220
rect 6460 12174 6512 12180
rect 6656 11830 6684 13466
rect 6840 12986 6868 13806
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6932 12866 6960 14894
rect 7024 13870 7052 15422
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7024 13326 7052 13398
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7116 12986 7144 14214
rect 7208 13870 7236 16934
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7300 13682 7328 18090
rect 7392 16794 7420 18788
rect 7852 18766 7880 19178
rect 7944 18902 7972 19178
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 8114 18864 8170 18873
rect 8114 18799 8116 18808
rect 8168 18799 8170 18808
rect 8116 18770 8168 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7576 16998 7604 18702
rect 7668 17882 7696 18702
rect 7803 18524 8111 18533
rect 7803 18522 7809 18524
rect 7865 18522 7889 18524
rect 7945 18522 7969 18524
rect 8025 18522 8049 18524
rect 8105 18522 8111 18524
rect 7865 18470 7867 18522
rect 8047 18470 8049 18522
rect 7803 18468 7809 18470
rect 7865 18468 7889 18470
rect 7945 18468 7969 18470
rect 8025 18468 8049 18470
rect 8105 18468 8111 18470
rect 7803 18459 8111 18468
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 8036 17678 8064 18022
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8128 17524 8156 18090
rect 8220 17864 8248 19774
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19446 8340 19654
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8404 19258 8432 19790
rect 8496 19514 8524 19790
rect 8680 19786 8708 20810
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 19854 8800 20198
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8668 19780 8720 19786
rect 8668 19722 8720 19728
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8312 19230 8432 19258
rect 8312 19174 8340 19230
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8312 18426 8340 19110
rect 8404 18970 8432 19110
rect 8588 19009 8616 19382
rect 8574 19000 8630 19009
rect 8392 18964 8444 18970
rect 8574 18935 8630 18944
rect 8392 18906 8444 18912
rect 8588 18902 8616 18935
rect 8576 18896 8628 18902
rect 8482 18864 8538 18873
rect 8576 18838 8628 18844
rect 8482 18799 8538 18808
rect 8496 18630 8524 18799
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8576 17876 8628 17882
rect 8220 17836 8432 17864
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8128 17496 8248 17524
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 8036 16658 8064 17070
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16250 7420 16390
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 13954 7420 15438
rect 7484 14618 7512 16594
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15026 7604 15982
rect 7668 15706 7696 16390
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14482 7604 14962
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14618 7880 14894
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 14074 7512 14350
rect 7576 14074 7604 14418
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7392 13926 7604 13954
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7208 13654 7328 13682
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7116 12889 7144 12922
rect 6840 12838 6960 12866
rect 7102 12880 7158 12889
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6748 12170 6776 12718
rect 6840 12458 6868 12838
rect 7102 12815 7158 12824
rect 7208 12628 7236 13654
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7300 12986 7328 13330
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7392 12866 7420 13806
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7484 12986 7512 13194
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7288 12844 7340 12850
rect 7392 12838 7512 12866
rect 7288 12786 7340 12792
rect 7116 12600 7236 12628
rect 6840 12430 6960 12458
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6196 11512 6776 11540
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6472 9722 6500 9998
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6472 9178 6500 9318
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6182 8936 6238 8945
rect 6104 8566 6132 8910
rect 6182 8871 6238 8880
rect 6196 8634 6224 8871
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6472 7886 6500 8774
rect 6564 8634 6592 9522
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6460 7336 6512 7342
rect 6564 7324 6592 7822
rect 6512 7296 6592 7324
rect 6460 7278 6512 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6472 6866 6500 7142
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6472 5710 6500 6326
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5234 6500 5646
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 5920 5052 6040 5080
rect 5920 4842 5948 5052
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 5724 4820 5776 4826
rect 5920 4814 6040 4842
rect 5724 4762 5776 4768
rect 5644 4690 5948 4706
rect 5644 4684 5960 4690
rect 5644 4678 5908 4684
rect 5908 4626 5960 4632
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5552 3194 5580 3538
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5736 800 5764 3878
rect 5920 3670 5948 4490
rect 6012 4078 6040 4814
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6104 4282 6132 4762
rect 6472 4690 6500 4966
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6104 3924 6132 4218
rect 6458 4176 6514 4185
rect 6564 4146 6592 7296
rect 6656 6866 6684 9998
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6656 5914 6684 6122
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6644 5228 6696 5234
rect 6748 5216 6776 11512
rect 6932 11098 6960 12430
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 11286 7052 11630
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7024 11150 7052 11222
rect 6840 11070 6960 11098
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6840 10452 6868 11070
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10606 6960 10950
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6840 10424 6960 10452
rect 6932 8634 6960 10424
rect 7024 9586 7052 11086
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6840 7857 6868 8434
rect 6826 7848 6882 7857
rect 6826 7783 6882 7792
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 6662 6868 7482
rect 6932 7410 6960 8570
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6338 6868 6598
rect 6840 6310 6960 6338
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5914 6868 6190
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6932 5778 6960 6310
rect 7024 5794 7052 7890
rect 7116 6866 7144 12600
rect 7300 11898 7328 12786
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12306 7420 12582
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7484 12186 7512 12838
rect 7392 12158 7512 12186
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7208 9994 7236 11562
rect 7300 11014 7328 11834
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7392 10130 7420 12158
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7484 9722 7512 10678
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 9110 7328 9318
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7546 7328 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7208 6254 7236 7346
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7300 5914 7328 6734
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5772 6972 5778
rect 7024 5766 7144 5794
rect 6920 5714 6972 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6696 5188 6868 5216
rect 6644 5170 6696 5176
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6656 4214 6684 4966
rect 6748 4826 6776 4966
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4690 6868 5188
rect 7024 5166 7052 5646
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6932 4826 6960 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 7024 4282 7052 5102
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6458 4111 6460 4120
rect 6512 4111 6514 4120
rect 6552 4140 6604 4146
rect 6460 4082 6512 4088
rect 6552 4082 6604 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6644 4072 6696 4078
rect 6012 3896 6132 3924
rect 6472 4020 6644 4026
rect 6472 4014 6696 4020
rect 6472 3998 6684 4014
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3058 5948 3606
rect 6012 3534 6040 3896
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 3194 6408 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6472 2446 6500 3998
rect 6644 3732 6696 3738
rect 6748 3720 6776 4082
rect 7116 3942 7144 5766
rect 7194 5400 7250 5409
rect 7194 5335 7250 5344
rect 7208 5234 7236 5335
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7392 4049 7420 7958
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7546 7512 7686
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7576 4298 7604 13926
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7760 13530 7788 13874
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 8220 13326 8248 17496
rect 8312 17134 8340 17682
rect 8404 17320 8432 17836
rect 8772 17864 8800 19790
rect 8628 17836 8800 17864
rect 8576 17818 8628 17824
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8404 17292 8616 17320
rect 8300 17128 8352 17134
rect 8352 17088 8524 17116
rect 8300 17070 8352 17076
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 14618 8340 15982
rect 8404 15706 8432 16050
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8404 15162 8432 15642
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8496 13530 8524 17088
rect 8588 15706 8616 17292
rect 8680 16454 8708 17478
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 11898 7696 13194
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 8300 12912 8352 12918
rect 7838 12880 7894 12889
rect 8300 12854 8352 12860
rect 7838 12815 7894 12824
rect 7852 12374 7880 12815
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 8312 11626 8340 12854
rect 8496 12306 8524 13466
rect 8588 13190 8616 14894
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8680 12434 8708 16390
rect 8772 15910 8800 16526
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8864 14260 8892 20878
rect 9036 20596 9088 20602
rect 9036 20538 9088 20544
rect 9048 20466 9076 20538
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8956 18902 8984 19110
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8956 18358 8984 18702
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 9048 16522 9076 20402
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 17338 9168 20198
rect 9232 19378 9260 21898
rect 9784 21690 9812 23200
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9517 21244 9825 21253
rect 9517 21242 9523 21244
rect 9579 21242 9603 21244
rect 9659 21242 9683 21244
rect 9739 21242 9763 21244
rect 9819 21242 9825 21244
rect 9579 21190 9581 21242
rect 9761 21190 9763 21242
rect 9517 21188 9523 21190
rect 9579 21188 9603 21190
rect 9659 21188 9683 21190
rect 9739 21188 9763 21190
rect 9819 21188 9825 21190
rect 9517 21179 9825 21188
rect 9876 20754 9904 22102
rect 10796 21690 10824 23310
rect 11242 23200 11298 24000
rect 11978 23200 12034 24000
rect 12714 23200 12770 24000
rect 13450 23200 13506 24000
rect 13910 23216 13966 23225
rect 11256 22094 11284 23200
rect 11428 22160 11480 22166
rect 11164 22066 11284 22094
rect 11426 22128 11428 22137
rect 11480 22128 11482 22137
rect 11164 21690 11192 22066
rect 11426 22063 11482 22072
rect 11230 21788 11538 21797
rect 11230 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11396 21788
rect 11452 21786 11476 21788
rect 11532 21786 11538 21788
rect 11292 21734 11294 21786
rect 11474 21734 11476 21786
rect 11230 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11396 21734
rect 11452 21732 11476 21734
rect 11532 21732 11538 21734
rect 11230 21723 11538 21732
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 9968 21146 9996 21490
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9692 20726 9904 20754
rect 9692 20330 9720 20726
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9517 20156 9825 20165
rect 9517 20154 9523 20156
rect 9579 20154 9603 20156
rect 9659 20154 9683 20156
rect 9739 20154 9763 20156
rect 9819 20154 9825 20156
rect 9579 20102 9581 20154
rect 9761 20102 9763 20154
rect 9517 20100 9523 20102
rect 9579 20100 9603 20102
rect 9659 20100 9683 20102
rect 9739 20100 9763 20102
rect 9819 20100 9825 20102
rect 9517 20091 9825 20100
rect 9876 20058 9904 20198
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9232 18290 9260 19314
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9324 17882 9352 19926
rect 9784 19514 9812 19994
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9416 19417 9444 19450
rect 9692 19417 9720 19450
rect 9864 19440 9916 19446
rect 9402 19408 9458 19417
rect 9402 19343 9458 19352
rect 9678 19408 9734 19417
rect 9864 19382 9916 19388
rect 9678 19343 9734 19352
rect 9517 19068 9825 19077
rect 9517 19066 9523 19068
rect 9579 19066 9603 19068
rect 9659 19066 9683 19068
rect 9739 19066 9763 19068
rect 9819 19066 9825 19068
rect 9579 19014 9581 19066
rect 9761 19014 9763 19066
rect 9517 19012 9523 19014
rect 9579 19012 9603 19014
rect 9659 19012 9683 19014
rect 9739 19012 9763 19014
rect 9819 19012 9825 19014
rect 9517 19003 9825 19012
rect 9876 18970 9904 19382
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9140 16794 9168 17274
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 15502 9260 15846
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14414 8984 15302
rect 9048 14618 9076 15438
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8864 14232 9076 14260
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8772 13394 8800 14010
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12850 8984 13126
rect 9048 13002 9076 14232
rect 9140 13938 9168 15302
rect 9324 15026 9352 16186
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9416 14958 9444 18158
rect 9692 18154 9720 18702
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9517 17980 9825 17989
rect 9517 17978 9523 17980
rect 9579 17978 9603 17980
rect 9659 17978 9683 17980
rect 9739 17978 9763 17980
rect 9819 17978 9825 17980
rect 9579 17926 9581 17978
rect 9761 17926 9763 17978
rect 9517 17924 9523 17926
rect 9579 17924 9603 17926
rect 9659 17924 9683 17926
rect 9739 17924 9763 17926
rect 9819 17924 9825 17926
rect 9517 17915 9825 17924
rect 9876 17678 9904 18022
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9692 17524 9720 17614
rect 9692 17496 9904 17524
rect 9876 17241 9904 17496
rect 9862 17232 9918 17241
rect 9862 17167 9918 17176
rect 9876 17134 9904 17167
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9968 16590 9996 20878
rect 10152 19446 10180 21422
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20602 10364 20742
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10060 17882 10088 19246
rect 10152 18834 10180 19246
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10152 17882 10180 18158
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10244 17814 10272 19654
rect 10336 18834 10364 20538
rect 10612 20466 10640 20878
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10612 19938 10640 20402
rect 10704 20058 10732 21490
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10428 19718 10456 19926
rect 10612 19910 10732 19938
rect 10796 19922 10824 20198
rect 10888 20058 10916 21082
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10980 20602 11008 20878
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10980 20346 11008 20538
rect 11072 20466 11100 21286
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11164 20466 11192 20742
rect 11230 20700 11538 20709
rect 11230 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11396 20700
rect 11452 20698 11476 20700
rect 11532 20698 11538 20700
rect 11292 20646 11294 20698
rect 11474 20646 11476 20698
rect 11230 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11396 20646
rect 11452 20644 11476 20646
rect 11532 20644 11538 20646
rect 11230 20635 11538 20644
rect 11624 20534 11652 21014
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 10980 20318 11100 20346
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10428 18290 10456 19246
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 17808 10284 17814
rect 10138 17776 10194 17785
rect 10232 17750 10284 17756
rect 10138 17711 10194 17720
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 17513 10088 17614
rect 10152 17610 10180 17711
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10232 17536 10284 17542
rect 10046 17504 10102 17513
rect 10232 17478 10284 17484
rect 10046 17439 10102 17448
rect 10244 16794 10272 17478
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16250 9628 16390
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9968 16182 9996 16526
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9692 15162 9720 15370
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9876 14618 9904 14894
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 13938 9352 14214
rect 9968 13938 9996 16118
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 14550 10088 15302
rect 10152 15162 10180 16458
rect 10336 16114 10364 18158
rect 10414 17776 10470 17785
rect 10414 17711 10470 17720
rect 10428 17270 10456 17711
rect 10520 17270 10548 19790
rect 10612 19417 10640 19790
rect 10704 19514 10732 19910
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10598 19408 10654 19417
rect 10598 19343 10654 19352
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 18834 10732 19110
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18290 10640 18702
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10598 18184 10654 18193
rect 10598 18119 10654 18128
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10612 17202 10640 18119
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10060 14074 10088 14350
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9126 13288 9182 13297
rect 9126 13223 9182 13232
rect 9140 13190 9168 13223
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9048 12974 9168 13002
rect 9232 12986 9260 13874
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 10060 13462 10088 14010
rect 10152 13530 10180 14962
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8680 12406 8800 12434
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8576 12300 8628 12306
rect 8772 12288 8800 12406
rect 8956 12356 8984 12786
rect 8956 12328 9076 12356
rect 8772 12260 8984 12288
rect 8576 12242 8628 12248
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 8220 10792 8248 10950
rect 8128 10764 8248 10792
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 8128 10062 8156 10764
rect 8312 10724 8340 11562
rect 8588 10792 8616 12242
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8220 10696 8340 10724
rect 8496 10764 8616 10792
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9450 7696 9930
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 7886 7696 8910
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 7886 7880 8434
rect 8220 7886 8248 10696
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9042 8340 9998
rect 8404 9586 8432 10406
rect 8496 10130 8524 10764
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8680 10266 8708 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 11354 8800 11698
rect 8864 11694 8892 12038
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8772 10810 8800 11290
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8496 9586 8524 10066
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8392 8968 8444 8974
rect 8312 8916 8392 8922
rect 8312 8910 8444 8916
rect 8312 8894 8432 8910
rect 8312 8634 8340 8894
rect 8588 8838 8616 9318
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8404 8634 8432 8774
rect 8588 8634 8616 8774
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7886 8432 8230
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 7668 7002 7696 7822
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 8220 7478 8248 7822
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 8312 6866 8340 7142
rect 8496 6934 8524 7686
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 5370 7696 6598
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 8312 6225 8340 6695
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6254 8432 6598
rect 8392 6248 8444 6254
rect 8298 6216 8354 6225
rect 8392 6190 8444 6196
rect 8298 6151 8354 6160
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7852 5710 7880 5782
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 7484 4270 7604 4298
rect 7378 4040 7434 4049
rect 7196 4004 7248 4010
rect 7378 3975 7434 3984
rect 7196 3946 7248 3952
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6696 3692 6776 3720
rect 6644 3674 6696 3680
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 2514 6684 3334
rect 7208 3194 7236 3946
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3194 7420 3878
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2514 6960 2790
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6184 2100 6236 2106
rect 6184 2042 6236 2048
rect 6196 1850 6224 2042
rect 7024 1850 7052 3062
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2446 7236 2790
rect 7484 2774 7512 4270
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7300 2746 7512 2774
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7300 2378 7328 2746
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 6196 1822 6500 1850
rect 7024 1822 7236 1850
rect 6472 800 6500 1822
rect 7208 800 7236 1822
rect 570 0 626 800
rect 1306 0 1362 800
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7576 762 7604 4082
rect 8220 4078 8248 5306
rect 8312 5234 8340 5714
rect 8680 5642 8708 9862
rect 8772 9722 8800 10542
rect 8864 10062 8892 11630
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8772 9178 8800 9658
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8956 7834 8984 12260
rect 8864 7806 8984 7834
rect 8760 6792 8812 6798
rect 8758 6760 8760 6769
rect 8812 6760 8814 6769
rect 8758 6695 8814 6704
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4758 8340 5170
rect 8496 4826 8524 5510
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8484 4616 8536 4622
rect 8536 4576 8616 4604
rect 8484 4558 8536 4564
rect 8312 4457 8340 4558
rect 8298 4448 8354 4457
rect 8298 4383 8354 4392
rect 8588 4146 8616 4576
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7852 3738 7880 4014
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 2514 7696 3606
rect 8128 3602 8156 3878
rect 8588 3738 8616 4082
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8864 3670 8892 7806
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 6322 8984 7686
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8956 4826 8984 5238
rect 9048 4826 9076 12328
rect 9140 8906 9168 12974
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9232 12306 9260 12922
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9232 11626 9260 12106
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9722 9260 9998
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7886 9168 8230
rect 9232 7886 9260 8978
rect 9324 7936 9352 13330
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12986 9720 13126
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 10244 12850 10272 15506
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14074 10364 14758
rect 10428 14482 10456 15506
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10324 13320 10376 13326
rect 10376 13280 10456 13308
rect 10324 13262 10376 13268
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9876 12238 9904 12582
rect 10336 12374 10364 12718
rect 10428 12374 10456 13280
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 10606 9444 12038
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 10244 11150 10272 11494
rect 10336 11354 10364 11494
rect 10428 11354 10456 12310
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10146 9996 10610
rect 10520 10282 10548 17070
rect 9876 10118 9996 10146
rect 10336 10254 10548 10282
rect 9876 10062 9904 10118
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9876 9654 9904 9998
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9876 8634 9904 9590
rect 10152 9586 10180 9862
rect 10244 9722 10272 9998
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10336 9110 10364 10254
rect 10704 9674 10732 17478
rect 10796 17082 10824 19722
rect 11072 19378 11100 20318
rect 11992 20058 12020 23200
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12070 21040 12126 21049
rect 12070 20975 12126 20984
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12084 19938 12112 20975
rect 12176 20942 12204 21082
rect 12268 20942 12296 21286
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12438 20360 12494 20369
rect 12438 20295 12494 20304
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11992 19910 12112 19938
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10980 18426 11008 18702
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11072 18358 11100 18702
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10888 17882 10916 18158
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17513 10916 17546
rect 10874 17504 10930 17513
rect 10874 17439 10930 17448
rect 10980 17270 11008 18090
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10796 17066 10916 17082
rect 11072 17066 11100 18158
rect 11164 17921 11192 19722
rect 11230 19612 11538 19621
rect 11230 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11396 19612
rect 11452 19610 11476 19612
rect 11532 19610 11538 19612
rect 11292 19558 11294 19610
rect 11474 19558 11476 19610
rect 11230 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11396 19558
rect 11452 19556 11476 19558
rect 11532 19556 11538 19558
rect 11230 19547 11538 19556
rect 11716 19514 11744 19790
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11532 18850 11560 19450
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11624 18970 11652 19382
rect 11702 19272 11758 19281
rect 11702 19207 11758 19216
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11716 18850 11744 19207
rect 11532 18822 11744 18850
rect 11230 18524 11538 18533
rect 11230 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11396 18524
rect 11452 18522 11476 18524
rect 11532 18522 11538 18524
rect 11292 18470 11294 18522
rect 11474 18470 11476 18522
rect 11230 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11396 18470
rect 11452 18468 11476 18470
rect 11532 18468 11538 18470
rect 11230 18459 11538 18468
rect 11716 18290 11744 18822
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11150 17912 11206 17921
rect 11150 17847 11206 17856
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 11624 17320 11652 18158
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11532 17292 11652 17320
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11440 17105 11468 17206
rect 11532 17202 11560 17292
rect 11716 17252 11744 18022
rect 11624 17224 11744 17252
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11426 17096 11482 17105
rect 10796 17060 10928 17066
rect 10796 17054 10876 17060
rect 10876 17002 10928 17008
rect 11060 17060 11112 17066
rect 11426 17031 11482 17040
rect 11060 17002 11112 17008
rect 11532 16726 11560 17138
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10796 15094 10824 15574
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10888 14482 10916 16050
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15502 11008 15982
rect 11164 15638 11192 16050
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11624 15570 11652 17224
rect 11808 16538 11836 19858
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11900 18154 11928 19246
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 17134 11928 17614
rect 11992 17610 12020 19910
rect 12176 19468 12388 19496
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12084 18630 12112 19382
rect 12176 19281 12204 19468
rect 12360 19378 12388 19468
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12162 19272 12218 19281
rect 12162 19207 12218 19216
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18970 12204 19110
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12176 18426 12204 18702
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17746 12112 18022
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12176 17610 12204 18226
rect 12268 18154 12296 19314
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12360 18222 12388 18906
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11992 17241 12020 17274
rect 11978 17232 12034 17241
rect 11978 17167 12034 17176
rect 12360 17134 12388 17614
rect 12452 17338 12480 20295
rect 12544 19854 12572 20742
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12636 19514 12664 21422
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 11716 16510 11836 16538
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 14074 10916 14418
rect 10980 14074 11008 14894
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10796 13462 10824 13806
rect 10980 13530 11008 14010
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10796 12986 10824 13398
rect 11072 12986 11100 15370
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11164 14006 11192 15030
rect 11624 14482 11652 15302
rect 11716 15162 11744 16510
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16114 11836 16390
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11900 15722 11928 17070
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11808 15694 11928 15722
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11716 15065 11744 15098
rect 11702 15056 11758 15065
rect 11702 14991 11758 15000
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 14618 11744 14758
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 11624 14074 11652 14214
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 11898 11008 12718
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11072 11626 11100 12174
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10612 9646 10732 9674
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9178 10456 9454
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10060 8566 10088 8910
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9324 7908 9444 7936
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5914 9168 6190
rect 9232 5914 9260 6258
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9324 5234 9352 6054
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 4282 9260 4558
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9218 4040 9274 4049
rect 9416 4026 9444 7908
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9876 6866 9904 8298
rect 9968 7750 9996 8366
rect 10060 8090 10088 8502
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7002 9996 7686
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10612 6882 10640 9646
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 8838 10732 9318
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 10980 8634 11008 8842
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7410 10916 7686
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11072 7018 11100 11562
rect 11164 11218 11192 13806
rect 11256 13394 11284 13874
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11354 11560 11494
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11428 11144 11480 11150
rect 11426 11112 11428 11121
rect 11480 11112 11482 11121
rect 11624 11098 11652 12271
rect 11716 12238 11744 13126
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11808 11370 11836 15694
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11900 13870 11928 15506
rect 11992 14278 12020 17002
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12084 15026 12112 16594
rect 12176 16522 12204 17070
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12360 16590 12388 16934
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12348 16448 12400 16454
rect 12268 16408 12348 16436
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12986 11928 13262
rect 11992 13190 12020 13806
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11900 12345 11928 12718
rect 11992 12646 12020 13126
rect 12084 12918 12112 13262
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11900 11898 11928 12106
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11808 11354 11928 11370
rect 11808 11348 11940 11354
rect 11808 11342 11888 11348
rect 11624 11070 11744 11098
rect 11426 11047 11482 11056
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11164 10266 11192 10610
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 10266 11468 10542
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11624 10062 11652 10950
rect 11716 10554 11744 11070
rect 11808 10674 11836 11342
rect 11888 11290 11940 11296
rect 11992 11234 12020 12582
rect 12176 11694 12204 14350
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11992 11206 12204 11234
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11716 10526 11836 10554
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 11164 9110 11192 9551
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11624 7886 11652 9998
rect 11808 8922 11836 10526
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12084 9058 12112 11086
rect 12176 10554 12204 11206
rect 12268 10674 12296 16408
rect 12452 16436 12480 16934
rect 12400 16408 12480 16436
rect 12348 16390 12400 16396
rect 12544 16250 12572 18226
rect 12636 17882 12664 19314
rect 12728 18970 12756 23200
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 21026 12848 21422
rect 12944 21244 13252 21253
rect 12944 21242 12950 21244
rect 13006 21242 13030 21244
rect 13086 21242 13110 21244
rect 13166 21242 13190 21244
rect 13246 21242 13252 21244
rect 13006 21190 13008 21242
rect 13188 21190 13190 21242
rect 12944 21188 12950 21190
rect 13006 21188 13030 21190
rect 13086 21188 13110 21190
rect 13166 21188 13190 21190
rect 13246 21188 13252 21190
rect 12944 21179 13252 21188
rect 12820 20998 12940 21026
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12820 17785 12848 20810
rect 12912 20369 12940 20998
rect 12898 20360 12954 20369
rect 12898 20295 12954 20304
rect 12912 20262 12940 20295
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12944 20156 13252 20165
rect 12944 20154 12950 20156
rect 13006 20154 13030 20156
rect 13086 20154 13110 20156
rect 13166 20154 13190 20156
rect 13246 20154 13252 20156
rect 13006 20102 13008 20154
rect 13188 20102 13190 20154
rect 12944 20100 12950 20102
rect 13006 20100 13030 20102
rect 13086 20100 13110 20102
rect 13166 20100 13190 20102
rect 13246 20100 13252 20102
rect 12944 20091 13252 20100
rect 13372 19922 13400 21626
rect 13464 20262 13492 23200
rect 14186 23200 14242 24000
rect 14922 23338 14978 24000
rect 14922 23310 15056 23338
rect 14922 23200 14978 23310
rect 13910 23151 13966 23160
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13556 20534 13584 21286
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13740 19990 13768 20198
rect 13728 19984 13780 19990
rect 13542 19952 13598 19961
rect 13360 19916 13412 19922
rect 13728 19926 13780 19932
rect 13542 19887 13598 19896
rect 13360 19858 13412 19864
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 19514 13308 19722
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13360 19372 13412 19378
rect 13280 19332 13360 19360
rect 12944 19068 13252 19077
rect 12944 19066 12950 19068
rect 13006 19066 13030 19068
rect 13086 19066 13110 19068
rect 13166 19066 13190 19068
rect 13246 19066 13252 19068
rect 13006 19014 13008 19066
rect 13188 19014 13190 19066
rect 12944 19012 12950 19014
rect 13006 19012 13030 19014
rect 13086 19012 13110 19014
rect 13166 19012 13190 19014
rect 13246 19012 13252 19014
rect 12944 19003 13252 19012
rect 12898 18728 12954 18737
rect 12898 18663 12900 18672
rect 12952 18663 12954 18672
rect 12900 18634 12952 18640
rect 12944 17980 13252 17989
rect 12944 17978 12950 17980
rect 13006 17978 13030 17980
rect 13086 17978 13110 17980
rect 13166 17978 13190 17980
rect 13246 17978 13252 17980
rect 13006 17926 13008 17978
rect 13188 17926 13190 17978
rect 12944 17924 12950 17926
rect 13006 17924 13030 17926
rect 13086 17924 13110 17926
rect 13166 17924 13190 17926
rect 13246 17924 13252 17926
rect 12944 17915 13252 17924
rect 12806 17776 12862 17785
rect 12806 17711 12862 17720
rect 13280 17626 13308 19332
rect 13360 19314 13412 19320
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 12636 17598 13308 17626
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12360 12374 12388 15574
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 15162 12480 15438
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12452 14618 12480 15098
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12452 14074 12480 14350
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13326 12572 14962
rect 12636 13954 12664 17598
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 16250 12756 17478
rect 13372 17338 13400 18022
rect 13464 17882 13492 18158
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16794 12848 17070
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 13280 16794 13308 17206
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 13280 16046 13308 16390
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12728 14482 12756 15914
rect 13280 15910 13308 15982
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12820 14618 12848 15574
rect 13280 15434 13308 15846
rect 13372 15706 13400 17274
rect 13464 16522 13492 17478
rect 13556 16590 13584 19887
rect 13740 18766 13768 19926
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13372 14074 13400 14282
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 12636 13926 12756 13954
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 13530 12664 13806
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 13410 12756 13926
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 13280 13530 13308 13806
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12636 13382 12756 13410
rect 13372 13394 13400 13806
rect 13360 13388 13412 13394
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12544 12442 12572 12786
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11762 12480 12038
rect 12544 11898 12572 12242
rect 12636 12238 12664 13382
rect 13360 13330 13412 13336
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12728 11762 12756 12582
rect 12820 12238 12848 12582
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12452 11218 12480 11698
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12636 11234 12664 11630
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12544 11206 12664 11234
rect 12820 11218 12848 12174
rect 13004 11898 13032 12174
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13280 11694 13308 13262
rect 13464 12306 13492 16186
rect 13648 16114 13676 17614
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13648 15094 13676 15846
rect 13740 15162 13768 17478
rect 13832 17134 13860 20742
rect 13924 18970 13952 23151
rect 14200 22094 14228 23200
rect 15028 22094 15056 23310
rect 14200 22066 14596 22094
rect 15028 22066 15148 22094
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 20874 14044 21286
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 19514 14044 20810
rect 14108 19718 14136 20878
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13910 18864 13966 18873
rect 13910 18799 13966 18808
rect 13924 18358 13952 18799
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 14016 18204 14044 19314
rect 14108 18902 14136 19654
rect 14200 19514 14228 20538
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 13924 18176 14044 18204
rect 13820 17128 13872 17134
rect 13924 17105 13952 18176
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14094 17640 14150 17649
rect 13820 17070 13872 17076
rect 13910 17096 13966 17105
rect 13910 17031 13966 17040
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 16250 13952 16390
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13832 15026 13860 16118
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13924 14550 13952 15370
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13556 12850 13584 13194
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13372 11898 13400 12106
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 12808 11212 12860 11218
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12176 10526 12296 10554
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9586 12204 9862
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 11716 8894 11836 8922
rect 11900 9030 12112 9058
rect 12176 9042 12204 9522
rect 12164 9036 12216 9042
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 11624 7410 11652 7822
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 10980 7002 11100 7018
rect 10980 6996 11112 7002
rect 10980 6990 11060 6996
rect 10784 6928 10836 6934
rect 9864 6860 9916 6866
rect 10612 6854 10732 6882
rect 10784 6870 10836 6876
rect 9864 6802 9916 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9864 5704 9916 5710
rect 9916 5664 9996 5692
rect 9864 5646 9916 5652
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5098 9628 5510
rect 9692 5370 9720 5578
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9678 5128 9734 5137
rect 9588 5092 9640 5098
rect 9784 5114 9812 5510
rect 9734 5086 9812 5114
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9678 5063 9734 5072
rect 9588 5034 9640 5040
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9772 4820 9824 4826
rect 9876 4808 9904 5102
rect 9968 5001 9996 5664
rect 9954 4992 10010 5001
rect 9954 4927 10010 4936
rect 9824 4780 9904 4808
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9772 4762 9824 4768
rect 9968 4706 9996 4791
rect 9784 4690 9996 4706
rect 9772 4684 9996 4690
rect 9824 4678 9996 4684
rect 9772 4626 9824 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4214 9628 4558
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9968 4298 9996 4422
rect 9692 4270 9996 4298
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9692 4078 9720 4270
rect 10060 4146 10088 6734
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10152 5234 10180 5782
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9680 4072 9732 4078
rect 9586 4040 9642 4049
rect 9218 3975 9274 3984
rect 9312 4004 9364 4010
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8116 3596 8168 3602
rect 8168 3556 8248 3584
rect 8116 3538 8168 3544
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 8220 2650 8248 3556
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 8404 2446 8432 2790
rect 8496 2650 8524 2994
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8772 2446 8800 3062
rect 9140 3058 9168 3470
rect 9232 3126 9260 3975
rect 9416 3998 9586 4026
rect 9680 4014 9732 4020
rect 9586 3975 9642 3984
rect 9312 3946 9364 3952
rect 9324 3738 9352 3946
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3466 9444 3878
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 9876 3738 9904 4082
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9968 2922 9996 4014
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 8220 2106 8248 2382
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8864 1170 8892 2246
rect 8680 1142 8892 1170
rect 7852 870 7972 898
rect 7852 762 7880 870
rect 7944 800 7972 870
rect 8680 800 8708 1142
rect 9416 800 9444 2790
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 10060 2582 10088 4082
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10152 2514 10180 4966
rect 10244 2582 10272 6598
rect 10336 5574 10364 6598
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4078 10364 4558
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10428 3942 10456 6734
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 5914 10548 6598
rect 10612 6390 10640 6734
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10704 5794 10732 6854
rect 10612 5766 10732 5794
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10520 4826 10548 5102
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3670 10456 3878
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10428 2514 10456 3606
rect 10612 3194 10640 5766
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5370 10732 5646
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10796 5273 10824 6870
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10888 5642 10916 6734
rect 10980 6118 11008 6990
rect 11060 6938 11112 6944
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10968 5568 11020 5574
rect 10888 5516 10968 5522
rect 10888 5510 11020 5516
rect 10888 5494 11008 5510
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10782 2952 10838 2961
rect 10888 2938 10916 5494
rect 10968 4480 11020 4486
rect 10966 4448 10968 4457
rect 11020 4448 11022 4457
rect 10966 4383 11022 4392
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10838 2910 10916 2938
rect 10782 2887 10838 2896
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10428 1170 10456 2314
rect 10152 1142 10456 1170
rect 10152 800 10180 1142
rect 10888 800 10916 2790
rect 10980 2650 11008 2994
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11072 2446 11100 6802
rect 11164 6390 11192 7210
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5556 11284 6326
rect 11624 6322 11652 7346
rect 11716 6905 11744 8894
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11808 7698 11836 8298
rect 11900 7800 11928 9030
rect 12164 8978 12216 8984
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 7868 12112 8434
rect 12176 8090 12204 8842
rect 12268 8362 12296 10526
rect 12544 10266 12572 11206
rect 12808 11154 12860 11160
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12636 9602 12664 11018
rect 13280 10674 13308 11154
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12990 10568 13046 10577
rect 12990 10503 12992 10512
rect 13044 10503 13046 10512
rect 12992 10474 13044 10480
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12452 9586 12664 9602
rect 12452 9580 12676 9586
rect 12452 9574 12624 9580
rect 12452 8922 12480 9574
rect 12624 9522 12676 9528
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12360 8894 12480 8922
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12162 7984 12218 7993
rect 12218 7942 12296 7970
rect 12162 7919 12218 7928
rect 12164 7880 12216 7886
rect 12084 7840 12164 7868
rect 12164 7822 12216 7828
rect 11900 7772 12112 7800
rect 11808 7670 11928 7698
rect 11702 6896 11758 6905
rect 11900 6866 11928 7670
rect 11702 6831 11758 6840
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6390 11744 6734
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11532 5914 11560 6054
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11624 5710 11652 6054
rect 11716 5914 11744 6190
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11164 5528 11284 5556
rect 11164 3942 11192 5528
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11256 5030 11284 5170
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11256 4690 11284 4966
rect 11532 4826 11560 5170
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11624 4826 11652 5102
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11716 4706 11744 5578
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11532 4678 11744 4706
rect 11532 4570 11560 4678
rect 11704 4616 11756 4622
rect 11532 4542 11652 4570
rect 11704 4558 11756 4564
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3466 11560 3878
rect 11624 3754 11652 4542
rect 11716 4214 11744 4558
rect 11808 4434 11836 6802
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11900 4622 11928 5646
rect 11992 5166 12020 6326
rect 12084 6118 12112 7772
rect 12176 7546 12204 7822
rect 12268 7562 12296 7942
rect 12360 7698 12388 8894
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 7818 12480 8774
rect 12544 8090 12572 9454
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 8838 12664 9318
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12624 8628 12676 8634
rect 12728 8616 12756 10202
rect 12820 9042 12848 10406
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13372 9994 13400 10950
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13556 9602 13584 12786
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11898 13676 12038
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13740 11762 13768 14214
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 10266 13676 10406
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13372 9574 13584 9602
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12728 8588 12848 8616
rect 12624 8570 12676 8576
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12360 7670 12572 7698
rect 12164 7540 12216 7546
rect 12268 7534 12388 7562
rect 12164 7482 12216 7488
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5370 12112 5646
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11808 4406 12020 4434
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11624 3726 11836 3754
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11164 3194 11192 3402
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11624 3194 11652 3334
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11808 2666 11836 3726
rect 11900 3398 11928 3975
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11886 2680 11942 2689
rect 11808 2638 11886 2666
rect 11886 2615 11942 2624
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11610 2408 11666 2417
rect 11610 2343 11612 2352
rect 11664 2343 11666 2352
rect 11612 2314 11664 2320
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 11624 870 11744 898
rect 11624 800 11652 870
rect 7576 734 7880 762
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 11716 762 11744 870
rect 11900 762 11928 2246
rect 11716 734 11928 762
rect 11992 354 12020 4406
rect 12084 3670 12112 4966
rect 12176 4690 12204 6190
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12084 3534 12112 3606
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12176 2650 12204 2926
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12268 1465 12296 4218
rect 12360 3058 12388 7534
rect 12544 7410 12572 7670
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6866 12480 7142
rect 12636 6934 12664 8570
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 7886 12756 8434
rect 12820 8378 12848 8588
rect 13280 8430 13308 9318
rect 13372 8634 13400 9574
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13464 9178 13492 9454
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 12992 8424 13044 8430
rect 12820 8372 12992 8378
rect 12820 8366 13044 8372
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12820 8350 13032 8366
rect 12820 7954 12848 8350
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 13266 7984 13322 7993
rect 12808 7948 12860 7954
rect 13266 7919 13322 7928
rect 12808 7890 12860 7896
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7546 13032 7822
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12820 6798 12848 7278
rect 13188 7274 13216 7346
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 13280 6798 13308 7919
rect 13372 7546 13400 8230
rect 13464 7886 13492 8910
rect 13556 8294 13584 9454
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7002 13492 7686
rect 13556 7018 13584 8026
rect 13648 7206 13676 10202
rect 13740 8498 13768 11018
rect 13832 10674 13860 13126
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13924 10418 13952 14486
rect 14016 13258 14044 17614
rect 14094 17575 14150 17584
rect 14108 17542 14136 17575
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14200 16114 14228 18566
rect 14292 16590 14320 20878
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 17202 14412 19654
rect 14476 18630 14504 21490
rect 14568 19514 14596 22066
rect 14657 21788 14965 21797
rect 14657 21786 14663 21788
rect 14719 21786 14743 21788
rect 14799 21786 14823 21788
rect 14879 21786 14903 21788
rect 14959 21786 14965 21788
rect 14719 21734 14721 21786
rect 14901 21734 14903 21786
rect 14657 21732 14663 21734
rect 14719 21732 14743 21734
rect 14799 21732 14823 21734
rect 14879 21732 14903 21734
rect 14959 21732 14965 21734
rect 14657 21723 14965 21732
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14657 20700 14965 20709
rect 14657 20698 14663 20700
rect 14719 20698 14743 20700
rect 14799 20698 14823 20700
rect 14879 20698 14903 20700
rect 14959 20698 14965 20700
rect 14719 20646 14721 20698
rect 14901 20646 14903 20698
rect 14657 20644 14663 20646
rect 14719 20644 14743 20646
rect 14799 20644 14823 20646
rect 14879 20644 14903 20646
rect 14959 20644 14965 20646
rect 14657 20635 14965 20644
rect 14657 19612 14965 19621
rect 14657 19610 14663 19612
rect 14719 19610 14743 19612
rect 14799 19610 14823 19612
rect 14879 19610 14903 19612
rect 14959 19610 14965 19612
rect 14719 19558 14721 19610
rect 14901 19558 14903 19610
rect 14657 19556 14663 19558
rect 14719 19556 14743 19558
rect 14799 19556 14823 19558
rect 14879 19556 14903 19558
rect 14959 19556 14965 19558
rect 14657 19547 14965 19556
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17785 14504 18022
rect 14462 17776 14518 17785
rect 14462 17711 14518 17720
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16697 14412 16934
rect 14370 16688 14426 16697
rect 14370 16623 14426 16632
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15609 14412 15846
rect 14370 15600 14426 15609
rect 14370 15535 14426 15544
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 14890 14320 15438
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14292 14414 14320 14826
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14521 14412 14758
rect 14370 14512 14426 14521
rect 14370 14447 14426 14456
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 14074 14136 14214
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14108 12442 14136 13874
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13433 14504 13670
rect 14462 13424 14518 13433
rect 14462 13359 14518 13368
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14016 10810 14044 11494
rect 14370 11248 14426 11257
rect 14370 11183 14372 11192
rect 14424 11183 14426 11192
rect 14372 11154 14424 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13832 10390 13952 10418
rect 13832 8566 13860 10390
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9722 13952 9998
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14016 9586 14044 10746
rect 14108 10266 14136 11086
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 9081 13952 9454
rect 14200 9178 14228 11086
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 13910 9072 13966 9081
rect 13910 9007 13966 9016
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 14016 7206 14044 9114
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 7886 14136 8230
rect 14200 7970 14228 8910
rect 14292 8634 14320 10610
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 10169 14412 10406
rect 14370 10160 14426 10169
rect 14370 10095 14426 10104
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14476 8090 14504 11018
rect 14568 10742 14596 19314
rect 14657 18524 14965 18533
rect 14657 18522 14663 18524
rect 14719 18522 14743 18524
rect 14799 18522 14823 18524
rect 14879 18522 14903 18524
rect 14959 18522 14965 18524
rect 14719 18470 14721 18522
rect 14901 18470 14903 18522
rect 14657 18468 14663 18470
rect 14719 18468 14743 18470
rect 14799 18468 14823 18470
rect 14879 18468 14903 18470
rect 14959 18468 14965 18470
rect 14657 18459 14965 18468
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 15028 16590 15056 21082
rect 15120 18193 15148 22066
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15106 18184 15162 18193
rect 15106 18119 15162 18128
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 15212 12850 15240 18702
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15304 12714 15332 19790
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12345 14964 12582
rect 14922 12336 14978 12345
rect 14922 12271 14978 12280
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14200 7942 14320 7970
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7546 14136 7686
rect 14200 7546 14228 7754
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13452 6996 13504 7002
rect 13556 6990 13676 7018
rect 13452 6938 13504 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5846 12572 6598
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5030 12480 5578
rect 12544 5370 12572 5782
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12636 5234 12664 6122
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12728 5098 12756 6326
rect 12820 5710 12848 6734
rect 13464 6458 13492 6938
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13450 6352 13506 6361
rect 13450 6287 13452 6296
rect 13504 6287 13506 6296
rect 13452 6258 13504 6264
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 13372 5914 13400 6190
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 4146 12940 4422
rect 12624 4140 12676 4146
rect 12900 4140 12952 4146
rect 12624 4082 12676 4088
rect 12820 4100 12900 4128
rect 12636 3738 12664 4082
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12820 3602 12848 4100
rect 12900 4082 12952 4088
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12820 3126 12848 3538
rect 13280 3126 13308 5714
rect 13648 5710 13676 6990
rect 13740 6905 13768 7142
rect 13726 6896 13782 6905
rect 13726 6831 13782 6840
rect 13832 6718 14044 6746
rect 13832 6662 13860 6718
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 13372 2650 13400 5102
rect 13556 4826 13584 5646
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12438 2544 12494 2553
rect 12438 2479 12494 2488
rect 12452 2446 12480 2479
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12254 1456 12310 1465
rect 12254 1391 12310 1400
rect 12360 800 12388 2246
rect 12728 2009 12756 2314
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12714 2000 12770 2009
rect 12714 1935 12770 1944
rect 13096 800 13124 2246
rect 13832 800 13860 6054
rect 13924 5234 13952 6598
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 14016 2446 14044 6718
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14108 6225 14136 6258
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 14292 5914 14320 7942
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 6798 14412 7278
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 4729 14136 5510
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14094 4720 14150 4729
rect 14094 4655 14150 4664
rect 14200 4593 14228 5034
rect 14292 4622 14320 5646
rect 14280 4616 14332 4622
rect 14186 4584 14242 4593
rect 14280 4558 14332 4564
rect 14186 4519 14242 4528
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3738 14136 4082
rect 14292 3754 14320 4558
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14200 3726 14320 3754
rect 14384 3738 14412 6734
rect 14462 5808 14518 5817
rect 14462 5743 14518 5752
rect 14372 3732 14424 3738
rect 14200 3534 14228 3726
rect 14372 3674 14424 3680
rect 14280 3664 14332 3670
rect 14278 3632 14280 3641
rect 14332 3632 14334 3641
rect 14278 3567 14334 3576
rect 14188 3528 14240 3534
rect 14108 3488 14188 3516
rect 14108 2650 14136 3488
rect 14188 3470 14240 3476
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 3058 14228 3334
rect 14476 3058 14504 5743
rect 14568 3534 14596 8774
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 15028 6769 15056 12174
rect 15014 6760 15070 6769
rect 15014 6695 15070 6704
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4729 14872 5170
rect 14830 4720 14886 4729
rect 14830 4655 14886 4664
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 2106 14228 2246
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14568 800 14596 2790
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 12070 368 12126 377
rect 11992 326 12070 354
rect 12070 303 12126 312
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
<< via2 >>
rect 938 20984 994 21040
rect 938 19896 994 19952
rect 938 18808 994 18864
rect 938 17720 994 17776
rect 938 16632 994 16688
rect 938 15544 994 15600
rect 1490 22072 1546 22128
rect 938 14456 994 14512
rect 1766 20712 1822 20768
rect 2134 20712 2190 20768
rect 2778 23160 2834 23216
rect 2669 21242 2725 21244
rect 2749 21242 2805 21244
rect 2829 21242 2885 21244
rect 2909 21242 2965 21244
rect 2669 21190 2715 21242
rect 2715 21190 2725 21242
rect 2749 21190 2779 21242
rect 2779 21190 2791 21242
rect 2791 21190 2805 21242
rect 2829 21190 2843 21242
rect 2843 21190 2855 21242
rect 2855 21190 2885 21242
rect 2909 21190 2919 21242
rect 2919 21190 2965 21242
rect 2669 21188 2725 21190
rect 2749 21188 2805 21190
rect 2829 21188 2885 21190
rect 2909 21188 2965 21190
rect 2669 20154 2725 20156
rect 2749 20154 2805 20156
rect 2829 20154 2885 20156
rect 2909 20154 2965 20156
rect 2669 20102 2715 20154
rect 2715 20102 2725 20154
rect 2749 20102 2779 20154
rect 2779 20102 2791 20154
rect 2791 20102 2805 20154
rect 2829 20102 2843 20154
rect 2843 20102 2855 20154
rect 2855 20102 2885 20154
rect 2909 20102 2919 20154
rect 2919 20102 2965 20154
rect 2669 20100 2725 20102
rect 2749 20100 2805 20102
rect 2829 20100 2885 20102
rect 2909 20100 2965 20102
rect 2502 19352 2558 19408
rect 1766 17604 1822 17640
rect 1766 17584 1768 17604
rect 1768 17584 1820 17604
rect 1820 17584 1822 17604
rect 938 12280 994 12336
rect 1398 11056 1454 11112
rect 1306 10104 1362 10160
rect 938 9016 994 9072
rect 1398 8200 1454 8256
rect 2669 19066 2725 19068
rect 2749 19066 2805 19068
rect 2829 19066 2885 19068
rect 2909 19066 2965 19068
rect 2669 19014 2715 19066
rect 2715 19014 2725 19066
rect 2749 19014 2779 19066
rect 2779 19014 2791 19066
rect 2791 19014 2805 19066
rect 2829 19014 2843 19066
rect 2843 19014 2855 19066
rect 2855 19014 2885 19066
rect 2909 19014 2919 19066
rect 2919 19014 2965 19066
rect 2669 19012 2725 19014
rect 2749 19012 2805 19014
rect 2829 19012 2885 19014
rect 2909 19012 2965 19014
rect 2669 17978 2725 17980
rect 2749 17978 2805 17980
rect 2829 17978 2885 17980
rect 2909 17978 2965 17980
rect 2669 17926 2715 17978
rect 2715 17926 2725 17978
rect 2749 17926 2779 17978
rect 2779 17926 2791 17978
rect 2791 17926 2805 17978
rect 2829 17926 2843 17978
rect 2843 17926 2855 17978
rect 2855 17926 2885 17978
rect 2909 17926 2919 17978
rect 2919 17926 2965 17978
rect 2669 17924 2725 17926
rect 2749 17924 2805 17926
rect 2829 17924 2885 17926
rect 2909 17924 2965 17926
rect 3422 20712 3478 20768
rect 4382 21786 4438 21788
rect 4462 21786 4518 21788
rect 4542 21786 4598 21788
rect 4622 21786 4678 21788
rect 4382 21734 4428 21786
rect 4428 21734 4438 21786
rect 4462 21734 4492 21786
rect 4492 21734 4504 21786
rect 4504 21734 4518 21786
rect 4542 21734 4556 21786
rect 4556 21734 4568 21786
rect 4568 21734 4598 21786
rect 4622 21734 4632 21786
rect 4632 21734 4678 21786
rect 4382 21732 4438 21734
rect 4462 21732 4518 21734
rect 4542 21732 4598 21734
rect 4622 21732 4678 21734
rect 4382 20698 4438 20700
rect 4462 20698 4518 20700
rect 4542 20698 4598 20700
rect 4622 20698 4678 20700
rect 4382 20646 4428 20698
rect 4428 20646 4438 20698
rect 4462 20646 4492 20698
rect 4492 20646 4504 20698
rect 4504 20646 4518 20698
rect 4542 20646 4556 20698
rect 4556 20646 4568 20698
rect 4568 20646 4598 20698
rect 4622 20646 4632 20698
rect 4632 20646 4678 20698
rect 4382 20644 4438 20646
rect 4462 20644 4518 20646
rect 4542 20644 4598 20646
rect 4622 20644 4678 20646
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 2410 14356 2412 14376
rect 2412 14356 2464 14376
rect 2464 14356 2466 14376
rect 2410 14320 2466 14356
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 938 6860 994 6896
rect 938 6840 940 6860
rect 940 6840 992 6860
rect 992 6840 994 6860
rect 1306 5752 1362 5808
rect 1674 6860 1730 6896
rect 1674 6840 1676 6860
rect 1676 6840 1728 6860
rect 1728 6840 1730 6860
rect 1674 6160 1730 6216
rect 938 4664 994 4720
rect 1950 7792 2006 7848
rect 938 3576 994 3632
rect 1674 3052 1730 3088
rect 1674 3032 1676 3052
rect 1676 3032 1728 3052
rect 1728 3032 1730 3052
rect 1398 2624 1454 2680
rect 1674 1808 1730 1864
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 3606 17176 3662 17232
rect 4382 19610 4438 19612
rect 4462 19610 4518 19612
rect 4542 19610 4598 19612
rect 4622 19610 4678 19612
rect 4382 19558 4428 19610
rect 4428 19558 4438 19610
rect 4462 19558 4492 19610
rect 4492 19558 4504 19610
rect 4504 19558 4518 19610
rect 4542 19558 4556 19610
rect 4556 19558 4568 19610
rect 4568 19558 4598 19610
rect 4622 19558 4632 19610
rect 4632 19558 4678 19610
rect 4382 19556 4438 19558
rect 4462 19556 4518 19558
rect 4542 19556 4598 19558
rect 4622 19556 4678 19558
rect 7809 21786 7865 21788
rect 7889 21786 7945 21788
rect 7969 21786 8025 21788
rect 8049 21786 8105 21788
rect 7809 21734 7855 21786
rect 7855 21734 7865 21786
rect 7889 21734 7919 21786
rect 7919 21734 7931 21786
rect 7931 21734 7945 21786
rect 7969 21734 7983 21786
rect 7983 21734 7995 21786
rect 7995 21734 8025 21786
rect 8049 21734 8059 21786
rect 8059 21734 8105 21786
rect 7809 21732 7865 21734
rect 7889 21732 7945 21734
rect 7969 21732 8025 21734
rect 8049 21732 8105 21734
rect 6096 21242 6152 21244
rect 6176 21242 6232 21244
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6096 21190 6142 21242
rect 6142 21190 6152 21242
rect 6176 21190 6206 21242
rect 6206 21190 6218 21242
rect 6218 21190 6232 21242
rect 6256 21190 6270 21242
rect 6270 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6096 21188 6152 21190
rect 6176 21188 6232 21190
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 4434 18808 4490 18864
rect 4710 18672 4766 18728
rect 4382 18522 4438 18524
rect 4462 18522 4518 18524
rect 4542 18522 4598 18524
rect 4622 18522 4678 18524
rect 4382 18470 4428 18522
rect 4428 18470 4438 18522
rect 4462 18470 4492 18522
rect 4492 18470 4504 18522
rect 4504 18470 4518 18522
rect 4542 18470 4556 18522
rect 4556 18470 4568 18522
rect 4568 18470 4598 18522
rect 4622 18470 4632 18522
rect 4632 18470 4678 18522
rect 4382 18468 4438 18470
rect 4462 18468 4518 18470
rect 4542 18468 4598 18470
rect 4622 18468 4678 18470
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 3422 9560 3478 9616
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2318 5752 2374 5808
rect 2042 4120 2098 4176
rect 2042 2524 2044 2544
rect 2044 2524 2096 2544
rect 2096 2524 2098 2544
rect 2042 2488 2098 2524
rect 1950 1400 2006 1456
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 3422 5072 3478 5128
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2778 3576 2834 3632
rect 2778 3440 2834 3496
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 3514 3032 3570 3088
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 5354 20712 5410 20768
rect 5722 20712 5778 20768
rect 6096 20154 6152 20156
rect 6176 20154 6232 20156
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6096 20102 6142 20154
rect 6142 20102 6152 20154
rect 6176 20102 6206 20154
rect 6206 20102 6218 20154
rect 6218 20102 6232 20154
rect 6256 20102 6270 20154
rect 6270 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6096 20100 6152 20102
rect 6176 20100 6232 20102
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 6096 19066 6152 19068
rect 6176 19066 6232 19068
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6096 19014 6142 19066
rect 6142 19014 6152 19066
rect 6176 19014 6206 19066
rect 6206 19014 6218 19066
rect 6218 19014 6232 19066
rect 6256 19014 6270 19066
rect 6270 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6096 19012 6152 19014
rect 6176 19012 6232 19014
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6096 17978 6152 17980
rect 6176 17978 6232 17980
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6096 17926 6142 17978
rect 6142 17926 6152 17978
rect 6176 17926 6206 17978
rect 6206 17926 6218 17978
rect 6218 17926 6232 17978
rect 6256 17926 6270 17978
rect 6270 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6096 17924 6152 17926
rect 6176 17924 6232 17926
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 5630 16652 5686 16688
rect 5630 16632 5632 16652
rect 5632 16632 5684 16652
rect 5684 16632 5686 16652
rect 4066 13404 4068 13424
rect 4068 13404 4120 13424
rect 4120 13404 4122 13424
rect 4066 13368 4122 13404
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 4710 12824 4766 12880
rect 4066 12588 4068 12608
rect 4068 12588 4120 12608
rect 4120 12588 4122 12608
rect 4066 12552 4122 12588
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4066 9632 4122 9688
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4066 9424 4122 9480
rect 3974 8916 3976 8936
rect 3976 8916 4028 8936
rect 4028 8916 4030 8936
rect 3974 8880 4030 8916
rect 3790 8200 3846 8256
rect 3790 4664 3846 4720
rect 4434 9288 4490 9344
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 7809 20698 7865 20700
rect 7889 20698 7945 20700
rect 7969 20698 8025 20700
rect 8049 20698 8105 20700
rect 7809 20646 7855 20698
rect 7855 20646 7865 20698
rect 7889 20646 7919 20698
rect 7919 20646 7931 20698
rect 7931 20646 7945 20698
rect 7969 20646 7983 20698
rect 7983 20646 7995 20698
rect 7995 20646 8025 20698
rect 8049 20646 8059 20698
rect 8059 20646 8105 20698
rect 7809 20644 7865 20646
rect 7889 20644 7945 20646
rect 7969 20644 8025 20646
rect 8049 20644 8105 20646
rect 8298 20712 8354 20768
rect 7809 19610 7865 19612
rect 7889 19610 7945 19612
rect 7969 19610 8025 19612
rect 8049 19610 8105 19612
rect 7809 19558 7855 19610
rect 7855 19558 7865 19610
rect 7889 19558 7919 19610
rect 7919 19558 7931 19610
rect 7931 19558 7945 19610
rect 7969 19558 7983 19610
rect 7983 19558 7995 19610
rect 7995 19558 8025 19610
rect 8049 19558 8059 19610
rect 8059 19558 8105 19610
rect 7809 19556 7865 19558
rect 7889 19556 7945 19558
rect 7969 19556 8025 19558
rect 8049 19556 8105 19558
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 5078 9560 5134 9616
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 4250 6296 4306 6352
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 5354 6704 5410 6760
rect 4986 5244 4988 5264
rect 4988 5244 5040 5264
rect 5040 5244 5042 5264
rect 4986 5208 5042 5244
rect 4250 4936 4306 4992
rect 4066 3984 4122 4040
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 5170 4528 5226 4584
rect 5262 3576 5318 3632
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 5354 3068 5356 3088
rect 5356 3068 5408 3088
rect 5408 3068 5410 3088
rect 5354 3032 5410 3068
rect 8114 18828 8170 18864
rect 8114 18808 8116 18828
rect 8116 18808 8168 18828
rect 8168 18808 8170 18828
rect 7809 18522 7865 18524
rect 7889 18522 7945 18524
rect 7969 18522 8025 18524
rect 8049 18522 8105 18524
rect 7809 18470 7855 18522
rect 7855 18470 7865 18522
rect 7889 18470 7919 18522
rect 7919 18470 7931 18522
rect 7931 18470 7945 18522
rect 7969 18470 7983 18522
rect 7983 18470 7995 18522
rect 7995 18470 8025 18522
rect 8049 18470 8059 18522
rect 8059 18470 8105 18522
rect 7809 18468 7865 18470
rect 7889 18468 7945 18470
rect 7969 18468 8025 18470
rect 8049 18468 8105 18470
rect 8574 18944 8630 19000
rect 8482 18808 8538 18864
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7102 12824 7158 12880
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6182 8880 6238 8936
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6458 4140 6514 4176
rect 6826 7792 6882 7848
rect 6458 4120 6460 4140
rect 6460 4120 6512 4140
rect 6512 4120 6514 4140
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 7194 5344 7250 5400
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 7838 12824 7894 12880
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 9523 21242 9579 21244
rect 9603 21242 9659 21244
rect 9683 21242 9739 21244
rect 9763 21242 9819 21244
rect 9523 21190 9569 21242
rect 9569 21190 9579 21242
rect 9603 21190 9633 21242
rect 9633 21190 9645 21242
rect 9645 21190 9659 21242
rect 9683 21190 9697 21242
rect 9697 21190 9709 21242
rect 9709 21190 9739 21242
rect 9763 21190 9773 21242
rect 9773 21190 9819 21242
rect 9523 21188 9579 21190
rect 9603 21188 9659 21190
rect 9683 21188 9739 21190
rect 9763 21188 9819 21190
rect 11426 22108 11428 22128
rect 11428 22108 11480 22128
rect 11480 22108 11482 22128
rect 11426 22072 11482 22108
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11396 21786 11452 21788
rect 11476 21786 11532 21788
rect 11236 21734 11282 21786
rect 11282 21734 11292 21786
rect 11316 21734 11346 21786
rect 11346 21734 11358 21786
rect 11358 21734 11372 21786
rect 11396 21734 11410 21786
rect 11410 21734 11422 21786
rect 11422 21734 11452 21786
rect 11476 21734 11486 21786
rect 11486 21734 11532 21786
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11396 21732 11452 21734
rect 11476 21732 11532 21734
rect 9523 20154 9579 20156
rect 9603 20154 9659 20156
rect 9683 20154 9739 20156
rect 9763 20154 9819 20156
rect 9523 20102 9569 20154
rect 9569 20102 9579 20154
rect 9603 20102 9633 20154
rect 9633 20102 9645 20154
rect 9645 20102 9659 20154
rect 9683 20102 9697 20154
rect 9697 20102 9709 20154
rect 9709 20102 9739 20154
rect 9763 20102 9773 20154
rect 9773 20102 9819 20154
rect 9523 20100 9579 20102
rect 9603 20100 9659 20102
rect 9683 20100 9739 20102
rect 9763 20100 9819 20102
rect 9402 19352 9458 19408
rect 9678 19352 9734 19408
rect 9523 19066 9579 19068
rect 9603 19066 9659 19068
rect 9683 19066 9739 19068
rect 9763 19066 9819 19068
rect 9523 19014 9569 19066
rect 9569 19014 9579 19066
rect 9603 19014 9633 19066
rect 9633 19014 9645 19066
rect 9645 19014 9659 19066
rect 9683 19014 9697 19066
rect 9697 19014 9709 19066
rect 9709 19014 9739 19066
rect 9763 19014 9773 19066
rect 9773 19014 9819 19066
rect 9523 19012 9579 19014
rect 9603 19012 9659 19014
rect 9683 19012 9739 19014
rect 9763 19012 9819 19014
rect 9523 17978 9579 17980
rect 9603 17978 9659 17980
rect 9683 17978 9739 17980
rect 9763 17978 9819 17980
rect 9523 17926 9569 17978
rect 9569 17926 9579 17978
rect 9603 17926 9633 17978
rect 9633 17926 9645 17978
rect 9645 17926 9659 17978
rect 9683 17926 9697 17978
rect 9697 17926 9709 17978
rect 9709 17926 9739 17978
rect 9763 17926 9773 17978
rect 9773 17926 9819 17978
rect 9523 17924 9579 17926
rect 9603 17924 9659 17926
rect 9683 17924 9739 17926
rect 9763 17924 9819 17926
rect 9862 17176 9918 17232
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11396 20698 11452 20700
rect 11476 20698 11532 20700
rect 11236 20646 11282 20698
rect 11282 20646 11292 20698
rect 11316 20646 11346 20698
rect 11346 20646 11358 20698
rect 11358 20646 11372 20698
rect 11396 20646 11410 20698
rect 11410 20646 11422 20698
rect 11422 20646 11452 20698
rect 11476 20646 11486 20698
rect 11486 20646 11532 20698
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11396 20644 11452 20646
rect 11476 20644 11532 20646
rect 10138 17720 10194 17776
rect 10046 17448 10102 17504
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 10414 17720 10470 17776
rect 10598 19352 10654 19408
rect 10598 18128 10654 18184
rect 9126 13232 9182 13288
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 8298 6704 8354 6760
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 8298 6160 8354 6216
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7378 3984 7434 4040
rect 8758 6740 8760 6760
rect 8760 6740 8812 6760
rect 8812 6740 8814 6760
rect 8758 6704 8814 6740
rect 8298 4392 8354 4448
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 12070 20984 12126 21040
rect 12438 20304 12494 20360
rect 10874 17448 10930 17504
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11396 19610 11452 19612
rect 11476 19610 11532 19612
rect 11236 19558 11282 19610
rect 11282 19558 11292 19610
rect 11316 19558 11346 19610
rect 11346 19558 11358 19610
rect 11358 19558 11372 19610
rect 11396 19558 11410 19610
rect 11410 19558 11422 19610
rect 11422 19558 11452 19610
rect 11476 19558 11486 19610
rect 11486 19558 11532 19610
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 11396 19556 11452 19558
rect 11476 19556 11532 19558
rect 11702 19216 11758 19272
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11396 18522 11452 18524
rect 11476 18522 11532 18524
rect 11236 18470 11282 18522
rect 11282 18470 11292 18522
rect 11316 18470 11346 18522
rect 11346 18470 11358 18522
rect 11358 18470 11372 18522
rect 11396 18470 11410 18522
rect 11410 18470 11422 18522
rect 11422 18470 11452 18522
rect 11476 18470 11486 18522
rect 11486 18470 11532 18522
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11396 18468 11452 18470
rect 11476 18468 11532 18470
rect 11150 17856 11206 17912
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 11426 17040 11482 17096
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 12162 19216 12218 19272
rect 11978 17176 12034 17232
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11702 15000 11758 15056
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 9218 3984 9274 4040
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 11610 12280 11666 12336
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 11426 11092 11428 11112
rect 11428 11092 11480 11112
rect 11480 11092 11482 11112
rect 11426 11056 11482 11092
rect 11886 12280 11942 12336
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 11150 9560 11206 9616
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 12950 21242 13006 21244
rect 13030 21242 13086 21244
rect 13110 21242 13166 21244
rect 13190 21242 13246 21244
rect 12950 21190 12996 21242
rect 12996 21190 13006 21242
rect 13030 21190 13060 21242
rect 13060 21190 13072 21242
rect 13072 21190 13086 21242
rect 13110 21190 13124 21242
rect 13124 21190 13136 21242
rect 13136 21190 13166 21242
rect 13190 21190 13200 21242
rect 13200 21190 13246 21242
rect 12950 21188 13006 21190
rect 13030 21188 13086 21190
rect 13110 21188 13166 21190
rect 13190 21188 13246 21190
rect 12898 20304 12954 20360
rect 12950 20154 13006 20156
rect 13030 20154 13086 20156
rect 13110 20154 13166 20156
rect 13190 20154 13246 20156
rect 12950 20102 12996 20154
rect 12996 20102 13006 20154
rect 13030 20102 13060 20154
rect 13060 20102 13072 20154
rect 13072 20102 13086 20154
rect 13110 20102 13124 20154
rect 13124 20102 13136 20154
rect 13136 20102 13166 20154
rect 13190 20102 13200 20154
rect 13200 20102 13246 20154
rect 12950 20100 13006 20102
rect 13030 20100 13086 20102
rect 13110 20100 13166 20102
rect 13190 20100 13246 20102
rect 13910 23160 13966 23216
rect 13542 19896 13598 19952
rect 12950 19066 13006 19068
rect 13030 19066 13086 19068
rect 13110 19066 13166 19068
rect 13190 19066 13246 19068
rect 12950 19014 12996 19066
rect 12996 19014 13006 19066
rect 13030 19014 13060 19066
rect 13060 19014 13072 19066
rect 13072 19014 13086 19066
rect 13110 19014 13124 19066
rect 13124 19014 13136 19066
rect 13136 19014 13166 19066
rect 13190 19014 13200 19066
rect 13200 19014 13246 19066
rect 12950 19012 13006 19014
rect 13030 19012 13086 19014
rect 13110 19012 13166 19014
rect 13190 19012 13246 19014
rect 12898 18692 12954 18728
rect 12898 18672 12900 18692
rect 12900 18672 12952 18692
rect 12952 18672 12954 18692
rect 12950 17978 13006 17980
rect 13030 17978 13086 17980
rect 13110 17978 13166 17980
rect 13190 17978 13246 17980
rect 12950 17926 12996 17978
rect 12996 17926 13006 17978
rect 13030 17926 13060 17978
rect 13060 17926 13072 17978
rect 13072 17926 13086 17978
rect 13110 17926 13124 17978
rect 13124 17926 13136 17978
rect 13136 17926 13166 17978
rect 13190 17926 13200 17978
rect 13200 17926 13246 17978
rect 12950 17924 13006 17926
rect 13030 17924 13086 17926
rect 13110 17924 13166 17926
rect 13190 17924 13246 17926
rect 12806 17720 12862 17776
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 13910 18808 13966 18864
rect 13910 17040 13966 17096
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9678 5072 9734 5128
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9954 4936 10010 4992
rect 9954 4800 10010 4856
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9586 3984 9642 4040
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 10782 5208 10838 5264
rect 10782 2896 10838 2952
rect 10966 4428 10968 4448
rect 10968 4428 11020 4448
rect 11020 4428 11022 4448
rect 10966 4392 11022 4428
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 12990 10532 13046 10568
rect 12990 10512 12992 10532
rect 12992 10512 13044 10532
rect 13044 10512 13046 10532
rect 12162 7928 12218 7984
rect 11702 6840 11758 6896
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 11886 3984 11942 4040
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 11886 2624 11942 2680
rect 11610 2372 11666 2408
rect 11610 2352 11612 2372
rect 11612 2352 11664 2372
rect 11664 2352 11666 2372
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 13266 7928 13322 7984
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 14094 17584 14150 17640
rect 14663 21786 14719 21788
rect 14743 21786 14799 21788
rect 14823 21786 14879 21788
rect 14903 21786 14959 21788
rect 14663 21734 14709 21786
rect 14709 21734 14719 21786
rect 14743 21734 14773 21786
rect 14773 21734 14785 21786
rect 14785 21734 14799 21786
rect 14823 21734 14837 21786
rect 14837 21734 14849 21786
rect 14849 21734 14879 21786
rect 14903 21734 14913 21786
rect 14913 21734 14959 21786
rect 14663 21732 14719 21734
rect 14743 21732 14799 21734
rect 14823 21732 14879 21734
rect 14903 21732 14959 21734
rect 14663 20698 14719 20700
rect 14743 20698 14799 20700
rect 14823 20698 14879 20700
rect 14903 20698 14959 20700
rect 14663 20646 14709 20698
rect 14709 20646 14719 20698
rect 14743 20646 14773 20698
rect 14773 20646 14785 20698
rect 14785 20646 14799 20698
rect 14823 20646 14837 20698
rect 14837 20646 14849 20698
rect 14849 20646 14879 20698
rect 14903 20646 14913 20698
rect 14913 20646 14959 20698
rect 14663 20644 14719 20646
rect 14743 20644 14799 20646
rect 14823 20644 14879 20646
rect 14903 20644 14959 20646
rect 14663 19610 14719 19612
rect 14743 19610 14799 19612
rect 14823 19610 14879 19612
rect 14903 19610 14959 19612
rect 14663 19558 14709 19610
rect 14709 19558 14719 19610
rect 14743 19558 14773 19610
rect 14773 19558 14785 19610
rect 14785 19558 14799 19610
rect 14823 19558 14837 19610
rect 14837 19558 14849 19610
rect 14849 19558 14879 19610
rect 14903 19558 14913 19610
rect 14913 19558 14959 19610
rect 14663 19556 14719 19558
rect 14743 19556 14799 19558
rect 14823 19556 14879 19558
rect 14903 19556 14959 19558
rect 14462 17720 14518 17776
rect 14370 16632 14426 16688
rect 14370 15544 14426 15600
rect 14370 14456 14426 14512
rect 14462 13368 14518 13424
rect 14370 11212 14426 11248
rect 14370 11192 14372 11212
rect 14372 11192 14424 11212
rect 14424 11192 14426 11212
rect 13910 9016 13966 9072
rect 14370 10104 14426 10160
rect 14663 18522 14719 18524
rect 14743 18522 14799 18524
rect 14823 18522 14879 18524
rect 14903 18522 14959 18524
rect 14663 18470 14709 18522
rect 14709 18470 14719 18522
rect 14743 18470 14773 18522
rect 14773 18470 14785 18522
rect 14785 18470 14799 18522
rect 14823 18470 14837 18522
rect 14837 18470 14849 18522
rect 14849 18470 14879 18522
rect 14903 18470 14913 18522
rect 14913 18470 14959 18522
rect 14663 18468 14719 18470
rect 14743 18468 14799 18470
rect 14823 18468 14879 18470
rect 14903 18468 14959 18470
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 15106 18128 15162 18184
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14922 12280 14978 12336
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 13450 6316 13506 6352
rect 13450 6296 13452 6316
rect 13452 6296 13504 6316
rect 13504 6296 13506 6316
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 13726 6840 13782 6896
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 12438 2488 12494 2544
rect 12254 1400 12310 1456
rect 12714 1944 12770 2000
rect 14094 6160 14150 6216
rect 14094 4664 14150 4720
rect 14186 4528 14242 4584
rect 14462 5752 14518 5808
rect 14278 3612 14280 3632
rect 14280 3612 14332 3632
rect 14332 3612 14334 3632
rect 14278 3576 14334 3612
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 15014 6704 15070 6760
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14830 4664 14886 4720
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 12070 312 12126 368
<< metal3 >>
rect 0 23218 800 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 800 23158
rect 2773 23155 2839 23158
rect 13905 23218 13971 23221
rect 15200 23218 16000 23248
rect 13905 23216 16000 23218
rect 13905 23160 13910 23216
rect 13966 23160 16000 23216
rect 13905 23158 16000 23160
rect 13905 23155 13971 23158
rect 15200 23128 16000 23158
rect 0 22130 800 22160
rect 1485 22130 1551 22133
rect 0 22128 1551 22130
rect 0 22072 1490 22128
rect 1546 22072 1551 22128
rect 0 22070 1551 22072
rect 0 22040 800 22070
rect 1485 22067 1551 22070
rect 11421 22130 11487 22133
rect 15200 22130 16000 22160
rect 11421 22128 16000 22130
rect 11421 22072 11426 22128
rect 11482 22072 16000 22128
rect 11421 22070 16000 22072
rect 11421 22067 11487 22070
rect 15200 22040 16000 22070
rect 4372 21792 4688 21793
rect 4372 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4688 21792
rect 4372 21727 4688 21728
rect 7799 21792 8115 21793
rect 7799 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8115 21792
rect 7799 21727 8115 21728
rect 11226 21792 11542 21793
rect 11226 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11542 21792
rect 11226 21727 11542 21728
rect 14653 21792 14969 21793
rect 14653 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14969 21792
rect 14653 21727 14969 21728
rect 2659 21248 2975 21249
rect 2659 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2975 21248
rect 2659 21183 2975 21184
rect 6086 21248 6402 21249
rect 6086 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6402 21248
rect 6086 21183 6402 21184
rect 9513 21248 9829 21249
rect 9513 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9829 21248
rect 9513 21183 9829 21184
rect 12940 21248 13256 21249
rect 12940 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13256 21248
rect 12940 21183 13256 21184
rect 0 21042 800 21072
rect 933 21042 999 21045
rect 0 21040 999 21042
rect 0 20984 938 21040
rect 994 20984 999 21040
rect 0 20982 999 20984
rect 0 20952 800 20982
rect 933 20979 999 20982
rect 12065 21042 12131 21045
rect 15200 21042 16000 21072
rect 12065 21040 16000 21042
rect 12065 20984 12070 21040
rect 12126 20984 16000 21040
rect 12065 20982 16000 20984
rect 12065 20979 12131 20982
rect 15200 20952 16000 20982
rect 1761 20770 1827 20773
rect 2129 20772 2195 20773
rect 1894 20770 1900 20772
rect 1761 20768 1900 20770
rect 1761 20712 1766 20768
rect 1822 20712 1900 20768
rect 1761 20710 1900 20712
rect 1761 20707 1827 20710
rect 1894 20708 1900 20710
rect 1964 20708 1970 20772
rect 2078 20770 2084 20772
rect 2038 20710 2084 20770
rect 2148 20768 2195 20772
rect 2190 20712 2195 20768
rect 2078 20708 2084 20710
rect 2148 20708 2195 20712
rect 2129 20707 2195 20708
rect 3417 20770 3483 20773
rect 5349 20772 5415 20773
rect 5717 20772 5783 20773
rect 8293 20772 8359 20773
rect 3550 20770 3556 20772
rect 3417 20768 3556 20770
rect 3417 20712 3422 20768
rect 3478 20712 3556 20768
rect 3417 20710 3556 20712
rect 3417 20707 3483 20710
rect 3550 20708 3556 20710
rect 3620 20708 3626 20772
rect 5349 20768 5396 20772
rect 5460 20770 5466 20772
rect 5349 20712 5354 20768
rect 5349 20708 5396 20712
rect 5460 20710 5506 20770
rect 5717 20768 5764 20772
rect 5828 20770 5834 20772
rect 5717 20712 5722 20768
rect 5460 20708 5466 20710
rect 5717 20708 5764 20712
rect 5828 20710 5874 20770
rect 8293 20768 8340 20772
rect 8404 20770 8410 20772
rect 8293 20712 8298 20768
rect 5828 20708 5834 20710
rect 8293 20708 8340 20712
rect 8404 20710 8450 20770
rect 8404 20708 8410 20710
rect 5349 20707 5415 20708
rect 5717 20707 5783 20708
rect 8293 20707 8359 20708
rect 4372 20704 4688 20705
rect 4372 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4688 20704
rect 4372 20639 4688 20640
rect 7799 20704 8115 20705
rect 7799 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8115 20704
rect 7799 20639 8115 20640
rect 11226 20704 11542 20705
rect 11226 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11542 20704
rect 11226 20639 11542 20640
rect 14653 20704 14969 20705
rect 14653 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14969 20704
rect 14653 20639 14969 20640
rect 12433 20362 12499 20365
rect 12893 20362 12959 20365
rect 12433 20360 12959 20362
rect 12433 20304 12438 20360
rect 12494 20304 12898 20360
rect 12954 20304 12959 20360
rect 12433 20302 12959 20304
rect 12433 20299 12499 20302
rect 12893 20299 12959 20302
rect 2659 20160 2975 20161
rect 2659 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2975 20160
rect 2659 20095 2975 20096
rect 6086 20160 6402 20161
rect 6086 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6402 20160
rect 6086 20095 6402 20096
rect 9513 20160 9829 20161
rect 9513 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9829 20160
rect 9513 20095 9829 20096
rect 12940 20160 13256 20161
rect 12940 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13256 20160
rect 12940 20095 13256 20096
rect 0 19954 800 19984
rect 933 19954 999 19957
rect 0 19952 999 19954
rect 0 19896 938 19952
rect 994 19896 999 19952
rect 0 19894 999 19896
rect 0 19864 800 19894
rect 933 19891 999 19894
rect 13537 19954 13603 19957
rect 15200 19954 16000 19984
rect 13537 19952 16000 19954
rect 13537 19896 13542 19952
rect 13598 19896 16000 19952
rect 13537 19894 16000 19896
rect 13537 19891 13603 19894
rect 15200 19864 16000 19894
rect 4372 19616 4688 19617
rect 4372 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4688 19616
rect 4372 19551 4688 19552
rect 7799 19616 8115 19617
rect 7799 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8115 19616
rect 7799 19551 8115 19552
rect 11226 19616 11542 19617
rect 11226 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11542 19616
rect 11226 19551 11542 19552
rect 14653 19616 14969 19617
rect 14653 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14969 19616
rect 14653 19551 14969 19552
rect 2262 19348 2268 19412
rect 2332 19410 2338 19412
rect 2497 19410 2563 19413
rect 2332 19408 2563 19410
rect 2332 19352 2502 19408
rect 2558 19352 2563 19408
rect 2332 19350 2563 19352
rect 2332 19348 2338 19350
rect 2497 19347 2563 19350
rect 9254 19348 9260 19412
rect 9324 19410 9330 19412
rect 9397 19410 9463 19413
rect 9324 19408 9463 19410
rect 9324 19352 9402 19408
rect 9458 19352 9463 19408
rect 9324 19350 9463 19352
rect 9324 19348 9330 19350
rect 9397 19347 9463 19350
rect 9673 19410 9739 19413
rect 9990 19410 9996 19412
rect 9673 19408 9996 19410
rect 9673 19352 9678 19408
rect 9734 19352 9996 19408
rect 9673 19350 9996 19352
rect 9673 19347 9739 19350
rect 9990 19348 9996 19350
rect 10060 19348 10066 19412
rect 10593 19410 10659 19413
rect 10726 19410 10732 19412
rect 10593 19408 10732 19410
rect 10593 19352 10598 19408
rect 10654 19352 10732 19408
rect 10593 19350 10732 19352
rect 10593 19347 10659 19350
rect 10726 19348 10732 19350
rect 10796 19348 10802 19412
rect 11697 19274 11763 19277
rect 12157 19274 12223 19277
rect 11697 19272 12223 19274
rect 11697 19216 11702 19272
rect 11758 19216 12162 19272
rect 12218 19216 12223 19272
rect 11697 19214 12223 19216
rect 11697 19211 11763 19214
rect 12157 19211 12223 19214
rect 2659 19072 2975 19073
rect 2659 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2975 19072
rect 2659 19007 2975 19008
rect 6086 19072 6402 19073
rect 6086 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6402 19072
rect 6086 19007 6402 19008
rect 9513 19072 9829 19073
rect 9513 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9829 19072
rect 9513 19007 9829 19008
rect 12940 19072 13256 19073
rect 12940 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13256 19072
rect 12940 19007 13256 19008
rect 8569 19002 8635 19005
rect 7974 19000 8635 19002
rect 7974 18944 8574 19000
rect 8630 18944 8635 19000
rect 7974 18942 8635 18944
rect 0 18866 800 18896
rect 933 18866 999 18869
rect 0 18864 999 18866
rect 0 18808 938 18864
rect 994 18808 999 18864
rect 0 18806 999 18808
rect 0 18776 800 18806
rect 933 18803 999 18806
rect 4429 18866 4495 18869
rect 7974 18866 8034 18942
rect 8569 18939 8635 18942
rect 4429 18864 8034 18866
rect 4429 18808 4434 18864
rect 4490 18808 8034 18864
rect 4429 18806 8034 18808
rect 8109 18866 8175 18869
rect 8477 18866 8543 18869
rect 8109 18864 8543 18866
rect 8109 18808 8114 18864
rect 8170 18808 8482 18864
rect 8538 18808 8543 18864
rect 8109 18806 8543 18808
rect 4429 18803 4495 18806
rect 8109 18803 8175 18806
rect 8477 18803 8543 18806
rect 13905 18866 13971 18869
rect 15200 18866 16000 18896
rect 13905 18864 16000 18866
rect 13905 18808 13910 18864
rect 13966 18808 16000 18864
rect 13905 18806 16000 18808
rect 13905 18803 13971 18806
rect 15200 18776 16000 18806
rect 4705 18730 4771 18733
rect 12893 18730 12959 18733
rect 4705 18728 12959 18730
rect 4705 18672 4710 18728
rect 4766 18672 12898 18728
rect 12954 18672 12959 18728
rect 4705 18670 12959 18672
rect 4705 18667 4771 18670
rect 12893 18667 12959 18670
rect 4372 18528 4688 18529
rect 4372 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4688 18528
rect 4372 18463 4688 18464
rect 7799 18528 8115 18529
rect 7799 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8115 18528
rect 7799 18463 8115 18464
rect 11226 18528 11542 18529
rect 11226 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11542 18528
rect 11226 18463 11542 18464
rect 14653 18528 14969 18529
rect 14653 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14969 18528
rect 14653 18463 14969 18464
rect 10593 18186 10659 18189
rect 15101 18186 15167 18189
rect 10593 18184 15167 18186
rect 10593 18128 10598 18184
rect 10654 18128 15106 18184
rect 15162 18128 15167 18184
rect 10593 18126 15167 18128
rect 10593 18123 10659 18126
rect 15101 18123 15167 18126
rect 2659 17984 2975 17985
rect 2659 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2975 17984
rect 2659 17919 2975 17920
rect 6086 17984 6402 17985
rect 6086 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6402 17984
rect 6086 17919 6402 17920
rect 9513 17984 9829 17985
rect 9513 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9829 17984
rect 9513 17919 9829 17920
rect 12940 17984 13256 17985
rect 12940 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13256 17984
rect 12940 17919 13256 17920
rect 11145 17914 11211 17917
rect 10182 17912 11211 17914
rect 10182 17856 11150 17912
rect 11206 17856 11211 17912
rect 10182 17854 11211 17856
rect 0 17778 800 17808
rect 10182 17781 10242 17854
rect 11145 17851 11211 17854
rect 933 17778 999 17781
rect 0 17776 999 17778
rect 0 17720 938 17776
rect 994 17720 999 17776
rect 0 17718 999 17720
rect 0 17688 800 17718
rect 933 17715 999 17718
rect 10133 17776 10242 17781
rect 10133 17720 10138 17776
rect 10194 17720 10242 17776
rect 10133 17718 10242 17720
rect 10409 17778 10475 17781
rect 12801 17778 12867 17781
rect 10409 17776 12867 17778
rect 10409 17720 10414 17776
rect 10470 17720 12806 17776
rect 12862 17720 12867 17776
rect 10409 17718 12867 17720
rect 10133 17715 10199 17718
rect 10409 17715 10475 17718
rect 12801 17715 12867 17718
rect 14457 17778 14523 17781
rect 15200 17778 16000 17808
rect 14457 17776 16000 17778
rect 14457 17720 14462 17776
rect 14518 17720 16000 17776
rect 14457 17718 16000 17720
rect 14457 17715 14523 17718
rect 15200 17688 16000 17718
rect 1761 17642 1827 17645
rect 14089 17642 14155 17645
rect 1761 17640 14155 17642
rect 1761 17584 1766 17640
rect 1822 17584 14094 17640
rect 14150 17584 14155 17640
rect 1761 17582 14155 17584
rect 1761 17579 1827 17582
rect 14089 17579 14155 17582
rect 10041 17506 10107 17509
rect 10869 17506 10935 17509
rect 10041 17504 10935 17506
rect 10041 17448 10046 17504
rect 10102 17448 10874 17504
rect 10930 17448 10935 17504
rect 10041 17446 10935 17448
rect 10041 17443 10107 17446
rect 10869 17443 10935 17446
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 3601 17236 3667 17237
rect 3550 17172 3556 17236
rect 3620 17234 3667 17236
rect 9857 17234 9923 17237
rect 11973 17234 12039 17237
rect 3620 17232 3712 17234
rect 3662 17176 3712 17232
rect 3620 17174 3712 17176
rect 9857 17232 12039 17234
rect 9857 17176 9862 17232
rect 9918 17176 11978 17232
rect 12034 17176 12039 17232
rect 9857 17174 12039 17176
rect 3620 17172 3667 17174
rect 3601 17171 3667 17172
rect 9857 17171 9923 17174
rect 11973 17171 12039 17174
rect 11421 17098 11487 17101
rect 13905 17098 13971 17101
rect 11421 17096 13971 17098
rect 11421 17040 11426 17096
rect 11482 17040 13910 17096
rect 13966 17040 13971 17096
rect 11421 17038 13971 17040
rect 11421 17035 11487 17038
rect 13905 17035 13971 17038
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 12940 16831 13256 16832
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 5625 16692 5691 16693
rect 5574 16690 5580 16692
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 5534 16630 5580 16690
rect 5644 16688 5691 16692
rect 5686 16632 5691 16688
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 5574 16628 5580 16630
rect 5644 16628 5691 16632
rect 5625 16627 5691 16628
rect 14365 16690 14431 16693
rect 15200 16690 16000 16720
rect 14365 16688 16000 16690
rect 14365 16632 14370 16688
rect 14426 16632 16000 16688
rect 14365 16630 16000 16632
rect 14365 16627 14431 16630
rect 15200 16600 16000 16630
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 0 15602 800 15632
rect 933 15602 999 15605
rect 0 15600 999 15602
rect 0 15544 938 15600
rect 994 15544 999 15600
rect 0 15542 999 15544
rect 0 15512 800 15542
rect 933 15539 999 15542
rect 14365 15602 14431 15605
rect 15200 15602 16000 15632
rect 14365 15600 16000 15602
rect 14365 15544 14370 15600
rect 14426 15544 16000 15600
rect 14365 15542 16000 15544
rect 14365 15539 14431 15542
rect 15200 15512 16000 15542
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 14653 15199 14969 15200
rect 11697 15058 11763 15061
rect 11830 15058 11836 15060
rect 11697 15056 11836 15058
rect 11697 15000 11702 15056
rect 11758 15000 11836 15056
rect 11697 14998 11836 15000
rect 11697 14995 11763 14998
rect 11830 14996 11836 14998
rect 11900 14996 11906 15060
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 0 14514 800 14544
rect 933 14514 999 14517
rect 0 14512 999 14514
rect 0 14456 938 14512
rect 994 14456 999 14512
rect 0 14454 999 14456
rect 0 14424 800 14454
rect 933 14451 999 14454
rect 14365 14514 14431 14517
rect 15200 14514 16000 14544
rect 14365 14512 16000 14514
rect 14365 14456 14370 14512
rect 14426 14456 16000 14512
rect 14365 14454 16000 14456
rect 14365 14451 14431 14454
rect 15200 14424 16000 14454
rect 2405 14378 2471 14381
rect 3182 14378 3188 14380
rect 2405 14376 3188 14378
rect 2405 14320 2410 14376
rect 2466 14320 3188 14376
rect 2405 14318 3188 14320
rect 2405 14315 2471 14318
rect 3182 14316 3188 14318
rect 3252 14316 3258 14380
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 0 13426 800 13456
rect 4061 13426 4127 13429
rect 0 13424 4127 13426
rect 0 13368 4066 13424
rect 4122 13368 4127 13424
rect 0 13366 4127 13368
rect 0 13336 800 13366
rect 4061 13363 4127 13366
rect 14457 13426 14523 13429
rect 15200 13426 16000 13456
rect 14457 13424 16000 13426
rect 14457 13368 14462 13424
rect 14518 13368 16000 13424
rect 14457 13366 16000 13368
rect 14457 13363 14523 13366
rect 15200 13336 16000 13366
rect 2078 13228 2084 13292
rect 2148 13290 2154 13292
rect 9121 13290 9187 13293
rect 2148 13288 9187 13290
rect 2148 13232 9126 13288
rect 9182 13232 9187 13288
rect 2148 13230 9187 13232
rect 2148 13228 2154 13230
rect 9121 13227 9187 13230
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 4705 12882 4771 12885
rect 4838 12882 4844 12884
rect 4705 12880 4844 12882
rect 4705 12824 4710 12880
rect 4766 12824 4844 12880
rect 4705 12822 4844 12824
rect 4705 12819 4771 12822
rect 4838 12820 4844 12822
rect 4908 12820 4914 12884
rect 7097 12882 7163 12885
rect 7833 12882 7899 12885
rect 7097 12880 7899 12882
rect 7097 12824 7102 12880
rect 7158 12824 7838 12880
rect 7894 12824 7899 12880
rect 7097 12822 7899 12824
rect 7097 12819 7163 12822
rect 7833 12819 7899 12822
rect 9070 12746 9076 12748
rect 5950 12686 9076 12746
rect 4061 12610 4127 12613
rect 5950 12610 6010 12686
rect 9070 12684 9076 12686
rect 9140 12684 9146 12748
rect 4061 12608 6010 12610
rect 4061 12552 4066 12608
rect 4122 12552 6010 12608
rect 4061 12550 6010 12552
rect 4061 12547 4127 12550
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 0 12338 800 12368
rect 933 12338 999 12341
rect 0 12336 999 12338
rect 0 12280 938 12336
rect 994 12280 999 12336
rect 0 12278 999 12280
rect 0 12248 800 12278
rect 933 12275 999 12278
rect 11605 12338 11671 12341
rect 11881 12338 11947 12341
rect 11605 12336 11947 12338
rect 11605 12280 11610 12336
rect 11666 12280 11886 12336
rect 11942 12280 11947 12336
rect 11605 12278 11947 12280
rect 11605 12275 11671 12278
rect 11881 12275 11947 12278
rect 14917 12338 14983 12341
rect 15200 12338 16000 12368
rect 14917 12336 16000 12338
rect 14917 12280 14922 12336
rect 14978 12280 16000 12336
rect 14917 12278 16000 12280
rect 14917 12275 14983 12278
rect 15200 12248 16000 12278
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 14653 11935 14969 11936
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 0 11250 800 11280
rect 14365 11250 14431 11253
rect 15200 11250 16000 11280
rect 0 11190 1456 11250
rect 0 11160 800 11190
rect 1396 11117 1456 11190
rect 14365 11248 16000 11250
rect 14365 11192 14370 11248
rect 14426 11192 16000 11248
rect 14365 11190 16000 11192
rect 14365 11187 14431 11190
rect 15200 11160 16000 11190
rect 1393 11112 1459 11117
rect 1393 11056 1398 11112
rect 1454 11056 1459 11112
rect 1393 11051 1459 11056
rect 8886 11052 8892 11116
rect 8956 11114 8962 11116
rect 11421 11114 11487 11117
rect 8956 11112 11487 11114
rect 8956 11056 11426 11112
rect 11482 11056 11487 11112
rect 8956 11054 11487 11056
rect 8956 11052 8962 11054
rect 11421 11051 11487 11054
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 1894 10508 1900 10572
rect 1964 10570 1970 10572
rect 12985 10570 13051 10573
rect 1964 10568 13051 10570
rect 1964 10512 12990 10568
rect 13046 10512 13051 10568
rect 1964 10510 13051 10512
rect 1964 10508 1970 10510
rect 12985 10507 13051 10510
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 0 10162 800 10192
rect 1301 10162 1367 10165
rect 0 10160 1367 10162
rect 0 10104 1306 10160
rect 1362 10104 1367 10160
rect 0 10102 1367 10104
rect 0 10072 800 10102
rect 1301 10099 1367 10102
rect 14365 10162 14431 10165
rect 15200 10162 16000 10192
rect 14365 10160 16000 10162
rect 14365 10104 14370 10160
rect 14426 10104 16000 10160
rect 14365 10102 16000 10104
rect 14365 10099 14431 10102
rect 15200 10072 16000 10102
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 4061 9688 4127 9693
rect 4061 9632 4066 9688
rect 4122 9632 4127 9688
rect 4061 9627 4127 9632
rect 3417 9618 3483 9621
rect 3550 9618 3556 9620
rect 3417 9616 3556 9618
rect 3417 9560 3422 9616
rect 3478 9560 3556 9616
rect 3417 9558 3556 9560
rect 3417 9555 3483 9558
rect 3550 9556 3556 9558
rect 3620 9556 3626 9620
rect 4064 9485 4124 9627
rect 5073 9620 5139 9621
rect 5022 9618 5028 9620
rect 4982 9558 5028 9618
rect 5092 9616 5139 9620
rect 5134 9560 5139 9616
rect 5022 9556 5028 9558
rect 5092 9556 5139 9560
rect 10726 9556 10732 9620
rect 10796 9618 10802 9620
rect 11145 9618 11211 9621
rect 10796 9616 11211 9618
rect 10796 9560 11150 9616
rect 11206 9560 11211 9616
rect 10796 9558 11211 9560
rect 10796 9556 10802 9558
rect 5073 9555 5139 9556
rect 11145 9555 11211 9558
rect 4061 9480 4127 9485
rect 4061 9424 4066 9480
rect 4122 9424 4127 9480
rect 4061 9419 4127 9424
rect 3366 9284 3372 9348
rect 3436 9346 3442 9348
rect 4429 9346 4495 9349
rect 3436 9344 4495 9346
rect 3436 9288 4434 9344
rect 4490 9288 4495 9344
rect 3436 9286 4495 9288
rect 3436 9284 3442 9286
rect 4429 9283 4495 9286
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 13905 9074 13971 9077
rect 15200 9074 16000 9104
rect 13905 9072 16000 9074
rect 13905 9016 13910 9072
rect 13966 9016 16000 9072
rect 13905 9014 16000 9016
rect 13905 9011 13971 9014
rect 15200 8984 16000 9014
rect 3969 8938 4035 8941
rect 6177 8938 6243 8941
rect 3969 8936 6243 8938
rect 3969 8880 3974 8936
rect 4030 8880 6182 8936
rect 6238 8880 6243 8936
rect 3969 8878 6243 8880
rect 3969 8875 4035 8878
rect 6177 8875 6243 8878
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 1393 8256 1459 8261
rect 1393 8200 1398 8256
rect 1454 8200 1459 8256
rect 1393 8195 1459 8200
rect 3182 8196 3188 8260
rect 3252 8258 3258 8260
rect 3785 8258 3851 8261
rect 3252 8256 3851 8258
rect 3252 8200 3790 8256
rect 3846 8200 3851 8256
rect 3252 8198 3851 8200
rect 3252 8196 3258 8198
rect 3785 8195 3851 8198
rect 0 7986 800 8016
rect 1396 7986 1456 8195
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 0 7926 1456 7986
rect 0 7896 800 7926
rect 9990 7924 9996 7988
rect 10060 7986 10066 7988
rect 12157 7986 12223 7989
rect 10060 7984 12223 7986
rect 10060 7928 12162 7984
rect 12218 7928 12223 7984
rect 10060 7926 12223 7928
rect 10060 7924 10066 7926
rect 12157 7923 12223 7926
rect 13261 7986 13327 7989
rect 15200 7986 16000 8016
rect 13261 7984 16000 7986
rect 13261 7928 13266 7984
rect 13322 7928 16000 7984
rect 13261 7926 16000 7928
rect 13261 7923 13327 7926
rect 15200 7896 16000 7926
rect 1945 7850 2011 7853
rect 6821 7850 6887 7853
rect 1945 7848 6887 7850
rect 1945 7792 1950 7848
rect 2006 7792 6826 7848
rect 6882 7792 6887 7848
rect 1945 7790 6887 7792
rect 1945 7787 2011 7790
rect 6821 7787 6887 7790
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 12940 7039 13256 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 1669 6898 1735 6901
rect 11697 6898 11763 6901
rect 1669 6896 11763 6898
rect 1669 6840 1674 6896
rect 1730 6840 11702 6896
rect 11758 6840 11763 6896
rect 1669 6838 11763 6840
rect 1669 6835 1735 6838
rect 11697 6835 11763 6838
rect 13721 6898 13787 6901
rect 15200 6898 16000 6928
rect 13721 6896 16000 6898
rect 13721 6840 13726 6896
rect 13782 6840 16000 6896
rect 13721 6838 16000 6840
rect 13721 6835 13787 6838
rect 15200 6808 16000 6838
rect 2262 6700 2268 6764
rect 2332 6762 2338 6764
rect 5349 6762 5415 6765
rect 2332 6760 5415 6762
rect 2332 6704 5354 6760
rect 5410 6704 5415 6760
rect 2332 6702 5415 6704
rect 2332 6700 2338 6702
rect 5349 6699 5415 6702
rect 8293 6762 8359 6765
rect 8753 6762 8819 6765
rect 15009 6762 15075 6765
rect 8293 6760 15075 6762
rect 8293 6704 8298 6760
rect 8354 6704 8758 6760
rect 8814 6704 15014 6760
rect 15070 6704 15075 6760
rect 8293 6702 15075 6704
rect 8293 6699 8359 6702
rect 8753 6699 8819 6702
rect 15009 6699 15075 6702
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 4245 6354 4311 6357
rect 13445 6354 13511 6357
rect 4245 6352 13511 6354
rect 4245 6296 4250 6352
rect 4306 6296 13450 6352
rect 13506 6296 13511 6352
rect 4245 6294 13511 6296
rect 4245 6291 4311 6294
rect 13445 6291 13511 6294
rect 1669 6218 1735 6221
rect 8293 6218 8359 6221
rect 1669 6216 8359 6218
rect 1669 6160 1674 6216
rect 1730 6160 8298 6216
rect 8354 6160 8359 6216
rect 1669 6158 8359 6160
rect 1669 6155 1735 6158
rect 8293 6155 8359 6158
rect 9254 6156 9260 6220
rect 9324 6218 9330 6220
rect 14089 6218 14155 6221
rect 9324 6216 14155 6218
rect 9324 6160 14094 6216
rect 14150 6160 14155 6216
rect 9324 6158 14155 6160
rect 9324 6156 9330 6158
rect 14089 6155 14155 6158
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 0 5810 800 5840
rect 1301 5810 1367 5813
rect 0 5808 1367 5810
rect 0 5752 1306 5808
rect 1362 5752 1367 5808
rect 0 5750 1367 5752
rect 0 5720 800 5750
rect 1301 5747 1367 5750
rect 2313 5810 2379 5813
rect 3366 5810 3372 5812
rect 2313 5808 3372 5810
rect 2313 5752 2318 5808
rect 2374 5752 3372 5808
rect 2313 5750 3372 5752
rect 2313 5747 2379 5750
rect 3366 5748 3372 5750
rect 3436 5748 3442 5812
rect 14457 5810 14523 5813
rect 15200 5810 16000 5840
rect 14457 5808 16000 5810
rect 14457 5752 14462 5808
rect 14518 5752 16000 5808
rect 14457 5750 16000 5752
rect 14457 5747 14523 5750
rect 15200 5720 16000 5750
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 5022 5340 5028 5404
rect 5092 5402 5098 5404
rect 7189 5402 7255 5405
rect 5092 5400 7255 5402
rect 5092 5344 7194 5400
rect 7250 5344 7255 5400
rect 5092 5342 7255 5344
rect 5092 5340 5098 5342
rect 7189 5339 7255 5342
rect 4981 5266 5047 5269
rect 10777 5266 10843 5269
rect 4981 5264 10843 5266
rect 4981 5208 4986 5264
rect 5042 5208 10782 5264
rect 10838 5208 10843 5264
rect 4981 5206 10843 5208
rect 4981 5203 5047 5206
rect 10777 5203 10843 5206
rect 3417 5130 3483 5133
rect 9673 5130 9739 5133
rect 3417 5128 9739 5130
rect 3417 5072 3422 5128
rect 3478 5072 9678 5128
rect 9734 5072 9739 5128
rect 3417 5070 9739 5072
rect 3417 5067 3483 5070
rect 9673 5067 9739 5070
rect 4245 4994 4311 4997
rect 5022 4994 5028 4996
rect 4245 4992 5028 4994
rect 4245 4936 4250 4992
rect 4306 4936 5028 4992
rect 4245 4934 5028 4936
rect 4245 4931 4311 4934
rect 5022 4932 5028 4934
rect 5092 4932 5098 4996
rect 9949 4994 10015 4997
rect 9949 4992 10058 4994
rect 9949 4936 9954 4992
rect 10010 4936 10058 4992
rect 9949 4931 10058 4936
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 9998 4861 10058 4931
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 9949 4856 10058 4861
rect 9949 4800 9954 4856
rect 10010 4800 10058 4856
rect 9949 4798 10058 4800
rect 9949 4795 10015 4798
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 3785 4722 3851 4725
rect 14089 4722 14155 4725
rect 3785 4720 14155 4722
rect 3785 4664 3790 4720
rect 3846 4664 14094 4720
rect 14150 4664 14155 4720
rect 3785 4662 14155 4664
rect 3785 4659 3851 4662
rect 14089 4659 14155 4662
rect 14825 4722 14891 4725
rect 15200 4722 16000 4752
rect 14825 4720 16000 4722
rect 14825 4664 14830 4720
rect 14886 4664 16000 4720
rect 14825 4662 16000 4664
rect 14825 4659 14891 4662
rect 15200 4632 16000 4662
rect 5165 4586 5231 4589
rect 14181 4586 14247 4589
rect 5165 4584 14247 4586
rect 5165 4528 5170 4584
rect 5226 4528 14186 4584
rect 14242 4528 14247 4584
rect 5165 4526 14247 4528
rect 5165 4523 5231 4526
rect 14181 4523 14247 4526
rect 8293 4450 8359 4453
rect 10961 4450 11027 4453
rect 8293 4448 11027 4450
rect 8293 4392 8298 4448
rect 8354 4392 10966 4448
rect 11022 4392 11027 4448
rect 8293 4390 11027 4392
rect 8293 4387 8359 4390
rect 10961 4387 11027 4390
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 2037 4178 2103 4181
rect 6453 4178 6519 4181
rect 2037 4176 6519 4178
rect 2037 4120 2042 4176
rect 2098 4120 6458 4176
rect 6514 4120 6519 4176
rect 2037 4118 6519 4120
rect 2037 4115 2103 4118
rect 6453 4115 6519 4118
rect 4061 4042 4127 4045
rect 7373 4042 7439 4045
rect 4061 4040 7439 4042
rect 4061 3984 4066 4040
rect 4122 3984 7378 4040
rect 7434 3984 7439 4040
rect 4061 3982 7439 3984
rect 4061 3979 4127 3982
rect 7373 3979 7439 3982
rect 9070 3980 9076 4044
rect 9140 4042 9146 4044
rect 9213 4042 9279 4045
rect 9140 4040 9279 4042
rect 9140 3984 9218 4040
rect 9274 3984 9279 4040
rect 9140 3982 9279 3984
rect 9140 3980 9146 3982
rect 9213 3979 9279 3982
rect 9581 4042 9647 4045
rect 11881 4042 11947 4045
rect 9581 4040 11947 4042
rect 9581 3984 9586 4040
rect 9642 3984 11886 4040
rect 11942 3984 11947 4040
rect 9581 3982 11947 3984
rect 9581 3979 9647 3982
rect 11881 3979 11947 3982
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 2773 3634 2839 3637
rect 5257 3634 5323 3637
rect 2773 3632 5323 3634
rect 2773 3576 2778 3632
rect 2834 3576 5262 3632
rect 5318 3576 5323 3632
rect 2773 3574 5323 3576
rect 2773 3571 2839 3574
rect 5257 3571 5323 3574
rect 14273 3634 14339 3637
rect 15200 3634 16000 3664
rect 14273 3632 16000 3634
rect 14273 3576 14278 3632
rect 14334 3576 16000 3632
rect 14273 3574 16000 3576
rect 14273 3571 14339 3574
rect 15200 3544 16000 3574
rect 2773 3498 2839 3501
rect 11830 3498 11836 3500
rect 2773 3496 11836 3498
rect 2773 3440 2778 3496
rect 2834 3440 11836 3496
rect 2773 3438 11836 3440
rect 2773 3435 2839 3438
rect 11830 3436 11836 3438
rect 11900 3436 11906 3500
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 1669 3090 1735 3093
rect 3509 3090 3575 3093
rect 5349 3090 5415 3093
rect 1669 3088 2790 3090
rect 1669 3032 1674 3088
rect 1730 3032 2790 3088
rect 1669 3030 2790 3032
rect 1669 3027 1735 3030
rect 2730 2954 2790 3030
rect 3509 3088 5415 3090
rect 3509 3032 3514 3088
rect 3570 3032 5354 3088
rect 5410 3032 5415 3088
rect 3509 3030 5415 3032
rect 3509 3027 3575 3030
rect 5349 3027 5415 3030
rect 10777 2954 10843 2957
rect 2730 2952 10843 2954
rect 2730 2896 10782 2952
rect 10838 2896 10843 2952
rect 2730 2894 10843 2896
rect 10777 2891 10843 2894
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 1393 2682 1459 2685
rect 798 2680 1459 2682
rect 798 2624 1398 2680
rect 1454 2624 1459 2680
rect 798 2622 1459 2624
rect 798 2576 858 2622
rect 1393 2619 1459 2622
rect 5574 2620 5580 2684
rect 5644 2620 5650 2684
rect 11881 2682 11947 2685
rect 11881 2680 12634 2682
rect 11881 2624 11886 2680
rect 11942 2624 12634 2680
rect 11881 2622 12634 2624
rect 0 2486 858 2576
rect 2037 2546 2103 2549
rect 5582 2546 5642 2620
rect 11881 2619 11947 2622
rect 2037 2544 5642 2546
rect 2037 2488 2042 2544
rect 2098 2488 5642 2544
rect 2037 2486 5642 2488
rect 0 2456 800 2486
rect 2037 2483 2103 2486
rect 5758 2484 5764 2548
rect 5828 2546 5834 2548
rect 12433 2546 12499 2549
rect 5828 2544 12499 2546
rect 5828 2488 12438 2544
rect 12494 2488 12499 2544
rect 5828 2486 12499 2488
rect 12574 2546 12634 2622
rect 15200 2546 16000 2576
rect 12574 2486 16000 2546
rect 5828 2484 5834 2486
rect 12433 2483 12499 2486
rect 15200 2456 16000 2486
rect 5390 2348 5396 2412
rect 5460 2410 5466 2412
rect 11605 2410 11671 2413
rect 5460 2408 11671 2410
rect 5460 2352 11610 2408
rect 11666 2352 11671 2408
rect 5460 2350 11671 2352
rect 5460 2348 5466 2350
rect 11605 2347 11671 2350
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 4838 1940 4844 2004
rect 4908 2002 4914 2004
rect 12709 2002 12775 2005
rect 4908 2000 12775 2002
rect 4908 1944 12714 2000
rect 12770 1944 12775 2000
rect 4908 1942 12775 1944
rect 4908 1940 4914 1942
rect 12709 1939 12775 1942
rect 1669 1866 1735 1869
rect 8886 1866 8892 1868
rect 1669 1864 8892 1866
rect 1669 1808 1674 1864
rect 1730 1808 8892 1864
rect 1669 1806 8892 1808
rect 1669 1803 1735 1806
rect 8886 1804 8892 1806
rect 8956 1804 8962 1868
rect 0 1458 800 1488
rect 1945 1458 2011 1461
rect 0 1456 2011 1458
rect 0 1400 1950 1456
rect 2006 1400 2011 1456
rect 0 1398 2011 1400
rect 0 1368 800 1398
rect 1945 1395 2011 1398
rect 12249 1458 12315 1461
rect 15200 1458 16000 1488
rect 12249 1456 16000 1458
rect 12249 1400 12254 1456
rect 12310 1400 16000 1456
rect 12249 1398 16000 1400
rect 12249 1395 12315 1398
rect 15200 1368 16000 1398
rect 12065 370 12131 373
rect 15200 370 16000 400
rect 12065 368 16000 370
rect 12065 312 12070 368
rect 12126 312 16000 368
rect 12065 310 16000 312
rect 12065 307 12131 310
rect 15200 280 16000 310
<< via3 >>
rect 4378 21788 4442 21792
rect 4378 21732 4382 21788
rect 4382 21732 4438 21788
rect 4438 21732 4442 21788
rect 4378 21728 4442 21732
rect 4458 21788 4522 21792
rect 4458 21732 4462 21788
rect 4462 21732 4518 21788
rect 4518 21732 4522 21788
rect 4458 21728 4522 21732
rect 4538 21788 4602 21792
rect 4538 21732 4542 21788
rect 4542 21732 4598 21788
rect 4598 21732 4602 21788
rect 4538 21728 4602 21732
rect 4618 21788 4682 21792
rect 4618 21732 4622 21788
rect 4622 21732 4678 21788
rect 4678 21732 4682 21788
rect 4618 21728 4682 21732
rect 7805 21788 7869 21792
rect 7805 21732 7809 21788
rect 7809 21732 7865 21788
rect 7865 21732 7869 21788
rect 7805 21728 7869 21732
rect 7885 21788 7949 21792
rect 7885 21732 7889 21788
rect 7889 21732 7945 21788
rect 7945 21732 7949 21788
rect 7885 21728 7949 21732
rect 7965 21788 8029 21792
rect 7965 21732 7969 21788
rect 7969 21732 8025 21788
rect 8025 21732 8029 21788
rect 7965 21728 8029 21732
rect 8045 21788 8109 21792
rect 8045 21732 8049 21788
rect 8049 21732 8105 21788
rect 8105 21732 8109 21788
rect 8045 21728 8109 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 11392 21788 11456 21792
rect 11392 21732 11396 21788
rect 11396 21732 11452 21788
rect 11452 21732 11456 21788
rect 11392 21728 11456 21732
rect 11472 21788 11536 21792
rect 11472 21732 11476 21788
rect 11476 21732 11532 21788
rect 11532 21732 11536 21788
rect 11472 21728 11536 21732
rect 14659 21788 14723 21792
rect 14659 21732 14663 21788
rect 14663 21732 14719 21788
rect 14719 21732 14723 21788
rect 14659 21728 14723 21732
rect 14739 21788 14803 21792
rect 14739 21732 14743 21788
rect 14743 21732 14799 21788
rect 14799 21732 14803 21788
rect 14739 21728 14803 21732
rect 14819 21788 14883 21792
rect 14819 21732 14823 21788
rect 14823 21732 14879 21788
rect 14879 21732 14883 21788
rect 14819 21728 14883 21732
rect 14899 21788 14963 21792
rect 14899 21732 14903 21788
rect 14903 21732 14959 21788
rect 14959 21732 14963 21788
rect 14899 21728 14963 21732
rect 2665 21244 2729 21248
rect 2665 21188 2669 21244
rect 2669 21188 2725 21244
rect 2725 21188 2729 21244
rect 2665 21184 2729 21188
rect 2745 21244 2809 21248
rect 2745 21188 2749 21244
rect 2749 21188 2805 21244
rect 2805 21188 2809 21244
rect 2745 21184 2809 21188
rect 2825 21244 2889 21248
rect 2825 21188 2829 21244
rect 2829 21188 2885 21244
rect 2885 21188 2889 21244
rect 2825 21184 2889 21188
rect 2905 21244 2969 21248
rect 2905 21188 2909 21244
rect 2909 21188 2965 21244
rect 2965 21188 2969 21244
rect 2905 21184 2969 21188
rect 6092 21244 6156 21248
rect 6092 21188 6096 21244
rect 6096 21188 6152 21244
rect 6152 21188 6156 21244
rect 6092 21184 6156 21188
rect 6172 21244 6236 21248
rect 6172 21188 6176 21244
rect 6176 21188 6232 21244
rect 6232 21188 6236 21244
rect 6172 21184 6236 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 9519 21244 9583 21248
rect 9519 21188 9523 21244
rect 9523 21188 9579 21244
rect 9579 21188 9583 21244
rect 9519 21184 9583 21188
rect 9599 21244 9663 21248
rect 9599 21188 9603 21244
rect 9603 21188 9659 21244
rect 9659 21188 9663 21244
rect 9599 21184 9663 21188
rect 9679 21244 9743 21248
rect 9679 21188 9683 21244
rect 9683 21188 9739 21244
rect 9739 21188 9743 21244
rect 9679 21184 9743 21188
rect 9759 21244 9823 21248
rect 9759 21188 9763 21244
rect 9763 21188 9819 21244
rect 9819 21188 9823 21244
rect 9759 21184 9823 21188
rect 12946 21244 13010 21248
rect 12946 21188 12950 21244
rect 12950 21188 13006 21244
rect 13006 21188 13010 21244
rect 12946 21184 13010 21188
rect 13026 21244 13090 21248
rect 13026 21188 13030 21244
rect 13030 21188 13086 21244
rect 13086 21188 13090 21244
rect 13026 21184 13090 21188
rect 13106 21244 13170 21248
rect 13106 21188 13110 21244
rect 13110 21188 13166 21244
rect 13166 21188 13170 21244
rect 13106 21184 13170 21188
rect 13186 21244 13250 21248
rect 13186 21188 13190 21244
rect 13190 21188 13246 21244
rect 13246 21188 13250 21244
rect 13186 21184 13250 21188
rect 1900 20708 1964 20772
rect 2084 20768 2148 20772
rect 2084 20712 2134 20768
rect 2134 20712 2148 20768
rect 2084 20708 2148 20712
rect 3556 20708 3620 20772
rect 5396 20768 5460 20772
rect 5396 20712 5410 20768
rect 5410 20712 5460 20768
rect 5396 20708 5460 20712
rect 5764 20768 5828 20772
rect 5764 20712 5778 20768
rect 5778 20712 5828 20768
rect 5764 20708 5828 20712
rect 8340 20768 8404 20772
rect 8340 20712 8354 20768
rect 8354 20712 8404 20768
rect 8340 20708 8404 20712
rect 4378 20700 4442 20704
rect 4378 20644 4382 20700
rect 4382 20644 4438 20700
rect 4438 20644 4442 20700
rect 4378 20640 4442 20644
rect 4458 20700 4522 20704
rect 4458 20644 4462 20700
rect 4462 20644 4518 20700
rect 4518 20644 4522 20700
rect 4458 20640 4522 20644
rect 4538 20700 4602 20704
rect 4538 20644 4542 20700
rect 4542 20644 4598 20700
rect 4598 20644 4602 20700
rect 4538 20640 4602 20644
rect 4618 20700 4682 20704
rect 4618 20644 4622 20700
rect 4622 20644 4678 20700
rect 4678 20644 4682 20700
rect 4618 20640 4682 20644
rect 7805 20700 7869 20704
rect 7805 20644 7809 20700
rect 7809 20644 7865 20700
rect 7865 20644 7869 20700
rect 7805 20640 7869 20644
rect 7885 20700 7949 20704
rect 7885 20644 7889 20700
rect 7889 20644 7945 20700
rect 7945 20644 7949 20700
rect 7885 20640 7949 20644
rect 7965 20700 8029 20704
rect 7965 20644 7969 20700
rect 7969 20644 8025 20700
rect 8025 20644 8029 20700
rect 7965 20640 8029 20644
rect 8045 20700 8109 20704
rect 8045 20644 8049 20700
rect 8049 20644 8105 20700
rect 8105 20644 8109 20700
rect 8045 20640 8109 20644
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 11392 20700 11456 20704
rect 11392 20644 11396 20700
rect 11396 20644 11452 20700
rect 11452 20644 11456 20700
rect 11392 20640 11456 20644
rect 11472 20700 11536 20704
rect 11472 20644 11476 20700
rect 11476 20644 11532 20700
rect 11532 20644 11536 20700
rect 11472 20640 11536 20644
rect 14659 20700 14723 20704
rect 14659 20644 14663 20700
rect 14663 20644 14719 20700
rect 14719 20644 14723 20700
rect 14659 20640 14723 20644
rect 14739 20700 14803 20704
rect 14739 20644 14743 20700
rect 14743 20644 14799 20700
rect 14799 20644 14803 20700
rect 14739 20640 14803 20644
rect 14819 20700 14883 20704
rect 14819 20644 14823 20700
rect 14823 20644 14879 20700
rect 14879 20644 14883 20700
rect 14819 20640 14883 20644
rect 14899 20700 14963 20704
rect 14899 20644 14903 20700
rect 14903 20644 14959 20700
rect 14959 20644 14963 20700
rect 14899 20640 14963 20644
rect 2665 20156 2729 20160
rect 2665 20100 2669 20156
rect 2669 20100 2725 20156
rect 2725 20100 2729 20156
rect 2665 20096 2729 20100
rect 2745 20156 2809 20160
rect 2745 20100 2749 20156
rect 2749 20100 2805 20156
rect 2805 20100 2809 20156
rect 2745 20096 2809 20100
rect 2825 20156 2889 20160
rect 2825 20100 2829 20156
rect 2829 20100 2885 20156
rect 2885 20100 2889 20156
rect 2825 20096 2889 20100
rect 2905 20156 2969 20160
rect 2905 20100 2909 20156
rect 2909 20100 2965 20156
rect 2965 20100 2969 20156
rect 2905 20096 2969 20100
rect 6092 20156 6156 20160
rect 6092 20100 6096 20156
rect 6096 20100 6152 20156
rect 6152 20100 6156 20156
rect 6092 20096 6156 20100
rect 6172 20156 6236 20160
rect 6172 20100 6176 20156
rect 6176 20100 6232 20156
rect 6232 20100 6236 20156
rect 6172 20096 6236 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 9519 20156 9583 20160
rect 9519 20100 9523 20156
rect 9523 20100 9579 20156
rect 9579 20100 9583 20156
rect 9519 20096 9583 20100
rect 9599 20156 9663 20160
rect 9599 20100 9603 20156
rect 9603 20100 9659 20156
rect 9659 20100 9663 20156
rect 9599 20096 9663 20100
rect 9679 20156 9743 20160
rect 9679 20100 9683 20156
rect 9683 20100 9739 20156
rect 9739 20100 9743 20156
rect 9679 20096 9743 20100
rect 9759 20156 9823 20160
rect 9759 20100 9763 20156
rect 9763 20100 9819 20156
rect 9819 20100 9823 20156
rect 9759 20096 9823 20100
rect 12946 20156 13010 20160
rect 12946 20100 12950 20156
rect 12950 20100 13006 20156
rect 13006 20100 13010 20156
rect 12946 20096 13010 20100
rect 13026 20156 13090 20160
rect 13026 20100 13030 20156
rect 13030 20100 13086 20156
rect 13086 20100 13090 20156
rect 13026 20096 13090 20100
rect 13106 20156 13170 20160
rect 13106 20100 13110 20156
rect 13110 20100 13166 20156
rect 13166 20100 13170 20156
rect 13106 20096 13170 20100
rect 13186 20156 13250 20160
rect 13186 20100 13190 20156
rect 13190 20100 13246 20156
rect 13246 20100 13250 20156
rect 13186 20096 13250 20100
rect 4378 19612 4442 19616
rect 4378 19556 4382 19612
rect 4382 19556 4438 19612
rect 4438 19556 4442 19612
rect 4378 19552 4442 19556
rect 4458 19612 4522 19616
rect 4458 19556 4462 19612
rect 4462 19556 4518 19612
rect 4518 19556 4522 19612
rect 4458 19552 4522 19556
rect 4538 19612 4602 19616
rect 4538 19556 4542 19612
rect 4542 19556 4598 19612
rect 4598 19556 4602 19612
rect 4538 19552 4602 19556
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 7805 19612 7869 19616
rect 7805 19556 7809 19612
rect 7809 19556 7865 19612
rect 7865 19556 7869 19612
rect 7805 19552 7869 19556
rect 7885 19612 7949 19616
rect 7885 19556 7889 19612
rect 7889 19556 7945 19612
rect 7945 19556 7949 19612
rect 7885 19552 7949 19556
rect 7965 19612 8029 19616
rect 7965 19556 7969 19612
rect 7969 19556 8025 19612
rect 8025 19556 8029 19612
rect 7965 19552 8029 19556
rect 8045 19612 8109 19616
rect 8045 19556 8049 19612
rect 8049 19556 8105 19612
rect 8105 19556 8109 19612
rect 8045 19552 8109 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 11392 19612 11456 19616
rect 11392 19556 11396 19612
rect 11396 19556 11452 19612
rect 11452 19556 11456 19612
rect 11392 19552 11456 19556
rect 11472 19612 11536 19616
rect 11472 19556 11476 19612
rect 11476 19556 11532 19612
rect 11532 19556 11536 19612
rect 11472 19552 11536 19556
rect 14659 19612 14723 19616
rect 14659 19556 14663 19612
rect 14663 19556 14719 19612
rect 14719 19556 14723 19612
rect 14659 19552 14723 19556
rect 14739 19612 14803 19616
rect 14739 19556 14743 19612
rect 14743 19556 14799 19612
rect 14799 19556 14803 19612
rect 14739 19552 14803 19556
rect 14819 19612 14883 19616
rect 14819 19556 14823 19612
rect 14823 19556 14879 19612
rect 14879 19556 14883 19612
rect 14819 19552 14883 19556
rect 14899 19612 14963 19616
rect 14899 19556 14903 19612
rect 14903 19556 14959 19612
rect 14959 19556 14963 19612
rect 14899 19552 14963 19556
rect 2268 19348 2332 19412
rect 9260 19348 9324 19412
rect 9996 19348 10060 19412
rect 10732 19348 10796 19412
rect 2665 19068 2729 19072
rect 2665 19012 2669 19068
rect 2669 19012 2725 19068
rect 2725 19012 2729 19068
rect 2665 19008 2729 19012
rect 2745 19068 2809 19072
rect 2745 19012 2749 19068
rect 2749 19012 2805 19068
rect 2805 19012 2809 19068
rect 2745 19008 2809 19012
rect 2825 19068 2889 19072
rect 2825 19012 2829 19068
rect 2829 19012 2885 19068
rect 2885 19012 2889 19068
rect 2825 19008 2889 19012
rect 2905 19068 2969 19072
rect 2905 19012 2909 19068
rect 2909 19012 2965 19068
rect 2965 19012 2969 19068
rect 2905 19008 2969 19012
rect 6092 19068 6156 19072
rect 6092 19012 6096 19068
rect 6096 19012 6152 19068
rect 6152 19012 6156 19068
rect 6092 19008 6156 19012
rect 6172 19068 6236 19072
rect 6172 19012 6176 19068
rect 6176 19012 6232 19068
rect 6232 19012 6236 19068
rect 6172 19008 6236 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 9519 19068 9583 19072
rect 9519 19012 9523 19068
rect 9523 19012 9579 19068
rect 9579 19012 9583 19068
rect 9519 19008 9583 19012
rect 9599 19068 9663 19072
rect 9599 19012 9603 19068
rect 9603 19012 9659 19068
rect 9659 19012 9663 19068
rect 9599 19008 9663 19012
rect 9679 19068 9743 19072
rect 9679 19012 9683 19068
rect 9683 19012 9739 19068
rect 9739 19012 9743 19068
rect 9679 19008 9743 19012
rect 9759 19068 9823 19072
rect 9759 19012 9763 19068
rect 9763 19012 9819 19068
rect 9819 19012 9823 19068
rect 9759 19008 9823 19012
rect 12946 19068 13010 19072
rect 12946 19012 12950 19068
rect 12950 19012 13006 19068
rect 13006 19012 13010 19068
rect 12946 19008 13010 19012
rect 13026 19068 13090 19072
rect 13026 19012 13030 19068
rect 13030 19012 13086 19068
rect 13086 19012 13090 19068
rect 13026 19008 13090 19012
rect 13106 19068 13170 19072
rect 13106 19012 13110 19068
rect 13110 19012 13166 19068
rect 13166 19012 13170 19068
rect 13106 19008 13170 19012
rect 13186 19068 13250 19072
rect 13186 19012 13190 19068
rect 13190 19012 13246 19068
rect 13246 19012 13250 19068
rect 13186 19008 13250 19012
rect 4378 18524 4442 18528
rect 4378 18468 4382 18524
rect 4382 18468 4438 18524
rect 4438 18468 4442 18524
rect 4378 18464 4442 18468
rect 4458 18524 4522 18528
rect 4458 18468 4462 18524
rect 4462 18468 4518 18524
rect 4518 18468 4522 18524
rect 4458 18464 4522 18468
rect 4538 18524 4602 18528
rect 4538 18468 4542 18524
rect 4542 18468 4598 18524
rect 4598 18468 4602 18524
rect 4538 18464 4602 18468
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 7805 18524 7869 18528
rect 7805 18468 7809 18524
rect 7809 18468 7865 18524
rect 7865 18468 7869 18524
rect 7805 18464 7869 18468
rect 7885 18524 7949 18528
rect 7885 18468 7889 18524
rect 7889 18468 7945 18524
rect 7945 18468 7949 18524
rect 7885 18464 7949 18468
rect 7965 18524 8029 18528
rect 7965 18468 7969 18524
rect 7969 18468 8025 18524
rect 8025 18468 8029 18524
rect 7965 18464 8029 18468
rect 8045 18524 8109 18528
rect 8045 18468 8049 18524
rect 8049 18468 8105 18524
rect 8105 18468 8109 18524
rect 8045 18464 8109 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 11392 18524 11456 18528
rect 11392 18468 11396 18524
rect 11396 18468 11452 18524
rect 11452 18468 11456 18524
rect 11392 18464 11456 18468
rect 11472 18524 11536 18528
rect 11472 18468 11476 18524
rect 11476 18468 11532 18524
rect 11532 18468 11536 18524
rect 11472 18464 11536 18468
rect 14659 18524 14723 18528
rect 14659 18468 14663 18524
rect 14663 18468 14719 18524
rect 14719 18468 14723 18524
rect 14659 18464 14723 18468
rect 14739 18524 14803 18528
rect 14739 18468 14743 18524
rect 14743 18468 14799 18524
rect 14799 18468 14803 18524
rect 14739 18464 14803 18468
rect 14819 18524 14883 18528
rect 14819 18468 14823 18524
rect 14823 18468 14879 18524
rect 14879 18468 14883 18524
rect 14819 18464 14883 18468
rect 14899 18524 14963 18528
rect 14899 18468 14903 18524
rect 14903 18468 14959 18524
rect 14959 18468 14963 18524
rect 14899 18464 14963 18468
rect 2665 17980 2729 17984
rect 2665 17924 2669 17980
rect 2669 17924 2725 17980
rect 2725 17924 2729 17980
rect 2665 17920 2729 17924
rect 2745 17980 2809 17984
rect 2745 17924 2749 17980
rect 2749 17924 2805 17980
rect 2805 17924 2809 17980
rect 2745 17920 2809 17924
rect 2825 17980 2889 17984
rect 2825 17924 2829 17980
rect 2829 17924 2885 17980
rect 2885 17924 2889 17980
rect 2825 17920 2889 17924
rect 2905 17980 2969 17984
rect 2905 17924 2909 17980
rect 2909 17924 2965 17980
rect 2965 17924 2969 17980
rect 2905 17920 2969 17924
rect 6092 17980 6156 17984
rect 6092 17924 6096 17980
rect 6096 17924 6152 17980
rect 6152 17924 6156 17980
rect 6092 17920 6156 17924
rect 6172 17980 6236 17984
rect 6172 17924 6176 17980
rect 6176 17924 6232 17980
rect 6232 17924 6236 17980
rect 6172 17920 6236 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 9519 17980 9583 17984
rect 9519 17924 9523 17980
rect 9523 17924 9579 17980
rect 9579 17924 9583 17980
rect 9519 17920 9583 17924
rect 9599 17980 9663 17984
rect 9599 17924 9603 17980
rect 9603 17924 9659 17980
rect 9659 17924 9663 17980
rect 9599 17920 9663 17924
rect 9679 17980 9743 17984
rect 9679 17924 9683 17980
rect 9683 17924 9739 17980
rect 9739 17924 9743 17980
rect 9679 17920 9743 17924
rect 9759 17980 9823 17984
rect 9759 17924 9763 17980
rect 9763 17924 9819 17980
rect 9819 17924 9823 17980
rect 9759 17920 9823 17924
rect 12946 17980 13010 17984
rect 12946 17924 12950 17980
rect 12950 17924 13006 17980
rect 13006 17924 13010 17980
rect 12946 17920 13010 17924
rect 13026 17980 13090 17984
rect 13026 17924 13030 17980
rect 13030 17924 13086 17980
rect 13086 17924 13090 17980
rect 13026 17920 13090 17924
rect 13106 17980 13170 17984
rect 13106 17924 13110 17980
rect 13110 17924 13166 17980
rect 13166 17924 13170 17980
rect 13106 17920 13170 17924
rect 13186 17980 13250 17984
rect 13186 17924 13190 17980
rect 13190 17924 13246 17980
rect 13246 17924 13250 17980
rect 13186 17920 13250 17924
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 3556 17232 3620 17236
rect 3556 17176 3606 17232
rect 3606 17176 3620 17232
rect 3556 17172 3620 17176
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 5580 16688 5644 16692
rect 5580 16632 5630 16688
rect 5630 16632 5644 16688
rect 5580 16628 5644 16632
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 11836 14996 11900 15060
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 3188 14316 3252 14380
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 2084 13228 2148 13292
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 4844 12820 4908 12884
rect 9076 12684 9140 12748
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 8892 11052 8956 11116
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 1900 10508 1964 10572
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 3556 9556 3620 9620
rect 5028 9616 5092 9620
rect 5028 9560 5078 9616
rect 5078 9560 5092 9616
rect 5028 9556 5092 9560
rect 10732 9556 10796 9620
rect 3372 9284 3436 9348
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 3188 8196 3252 8260
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 9996 7924 10060 7988
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 2268 6700 2332 6764
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 9260 6156 9324 6220
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 3372 5748 3436 5812
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 5028 5340 5092 5404
rect 5028 4932 5092 4996
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 9076 3980 9140 4044
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 11836 3436 11900 3500
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 5580 2620 5644 2684
rect 5764 2484 5828 2548
rect 5396 2348 5460 2412
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
rect 4844 1940 4908 2004
rect 8892 1804 8956 1868
<< metal4 >>
rect 2657 21248 2977 21808
rect 2657 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2977 21248
rect 1899 20772 1965 20773
rect 1899 20708 1900 20772
rect 1964 20708 1965 20772
rect 1899 20707 1965 20708
rect 2083 20772 2149 20773
rect 2083 20708 2084 20772
rect 2148 20708 2149 20772
rect 2083 20707 2149 20708
rect 1902 10573 1962 20707
rect 2086 13293 2146 20707
rect 2657 20160 2977 21184
rect 4370 21792 4690 21808
rect 4370 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4690 21792
rect 3555 20772 3621 20773
rect 3555 20708 3556 20772
rect 3620 20708 3621 20772
rect 3555 20707 3621 20708
rect 2657 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2977 20160
rect 2267 19412 2333 19413
rect 2267 19348 2268 19412
rect 2332 19348 2333 19412
rect 2267 19347 2333 19348
rect 2083 13292 2149 13293
rect 2083 13228 2084 13292
rect 2148 13228 2149 13292
rect 2083 13227 2149 13228
rect 1899 10572 1965 10573
rect 1899 10508 1900 10572
rect 1964 10508 1965 10572
rect 1899 10507 1965 10508
rect 2270 6765 2330 19347
rect 2657 19072 2977 20096
rect 2657 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2977 19072
rect 2657 17984 2977 19008
rect 2657 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2977 17984
rect 2657 16896 2977 17920
rect 3558 17237 3618 20707
rect 4370 20704 4690 21728
rect 6084 21248 6404 21808
rect 6084 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6404 21248
rect 5395 20772 5461 20773
rect 5395 20708 5396 20772
rect 5460 20708 5461 20772
rect 5395 20707 5461 20708
rect 5763 20772 5829 20773
rect 5763 20708 5764 20772
rect 5828 20708 5829 20772
rect 5763 20707 5829 20708
rect 4370 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4690 20704
rect 4370 19616 4690 20640
rect 4370 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4690 19616
rect 4370 18528 4690 19552
rect 4370 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4690 18528
rect 4370 17440 4690 18464
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 3555 17236 3621 17237
rect 3555 17172 3556 17236
rect 3620 17172 3621 17236
rect 3555 17171 3621 17172
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 3187 14380 3253 14381
rect 3187 14316 3188 14380
rect 3252 14316 3253 14380
rect 3187 14315 3253 14316
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 3190 8261 3250 14315
rect 3558 9621 3618 17171
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4843 12884 4909 12885
rect 4843 12820 4844 12884
rect 4908 12820 4909 12884
rect 4843 12819 4909 12820
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 3555 9620 3621 9621
rect 3555 9556 3556 9620
rect 3620 9556 3621 9620
rect 3555 9555 3621 9556
rect 3371 9348 3437 9349
rect 3371 9284 3372 9348
rect 3436 9284 3437 9348
rect 3371 9283 3437 9284
rect 3187 8260 3253 8261
rect 3187 8196 3188 8260
rect 3252 8196 3253 8260
rect 3187 8195 3253 8196
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2267 6764 2333 6765
rect 2267 6700 2268 6764
rect 2332 6700 2333 6764
rect 2267 6699 2333 6700
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 3374 5813 3434 9283
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 3371 5812 3437 5813
rect 3371 5748 3372 5812
rect 3436 5748 3437 5812
rect 3371 5747 3437 5748
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 4846 2005 4906 12819
rect 5027 9620 5093 9621
rect 5027 9556 5028 9620
rect 5092 9556 5093 9620
rect 5027 9555 5093 9556
rect 5030 5405 5090 9555
rect 5027 5404 5093 5405
rect 5027 5340 5028 5404
rect 5092 5340 5093 5404
rect 5027 5339 5093 5340
rect 5030 4997 5090 5339
rect 5027 4996 5093 4997
rect 5027 4932 5028 4996
rect 5092 4932 5093 4996
rect 5027 4931 5093 4932
rect 5398 2413 5458 20707
rect 5579 16692 5645 16693
rect 5579 16628 5580 16692
rect 5644 16628 5645 16692
rect 5579 16627 5645 16628
rect 5582 2685 5642 16627
rect 5579 2684 5645 2685
rect 5579 2620 5580 2684
rect 5644 2620 5645 2684
rect 5579 2619 5645 2620
rect 5766 2549 5826 20707
rect 6084 20160 6404 21184
rect 6084 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6404 20160
rect 6084 19072 6404 20096
rect 6084 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6404 19072
rect 6084 17984 6404 19008
rect 6084 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6404 17984
rect 6084 16896 6404 17920
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 5763 2548 5829 2549
rect 5763 2484 5764 2548
rect 5828 2484 5829 2548
rect 5763 2483 5829 2484
rect 5395 2412 5461 2413
rect 5395 2348 5396 2412
rect 5460 2348 5461 2412
rect 5395 2347 5461 2348
rect 6084 2128 6404 2688
rect 7797 21792 8117 21808
rect 7797 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8117 21792
rect 7797 20704 8117 21728
rect 9511 21248 9831 21808
rect 9511 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9831 21248
rect 8339 20772 8405 20773
rect 8339 20708 8340 20772
rect 8404 20708 8405 20772
rect 8339 20707 8405 20708
rect 7797 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8117 20704
rect 7797 19616 8117 20640
rect 7797 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8117 19616
rect 7797 18528 8117 19552
rect 7797 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8117 18528
rect 7797 17440 8117 18464
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 8342 12450 8402 20707
rect 9511 20160 9831 21184
rect 9511 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9831 20160
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 9075 12748 9141 12749
rect 9075 12684 9076 12748
rect 9140 12684 9141 12748
rect 9075 12683 9141 12684
rect 8342 12390 8954 12450
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 8894 11117 8954 12390
rect 8891 11116 8957 11117
rect 8891 11052 8892 11116
rect 8956 11052 8957 11116
rect 8891 11051 8957 11052
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 4843 2004 4909 2005
rect 4843 1940 4844 2004
rect 4908 1940 4909 2004
rect 4843 1939 4909 1940
rect 8894 1869 8954 11051
rect 9078 4045 9138 12683
rect 9262 6221 9322 19347
rect 9511 19072 9831 20096
rect 11224 21792 11544 21808
rect 11224 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11544 21792
rect 11224 20704 11544 21728
rect 11224 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11544 20704
rect 11224 19616 11544 20640
rect 11224 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11544 19616
rect 9995 19412 10061 19413
rect 9995 19348 9996 19412
rect 10060 19348 10061 19412
rect 9995 19347 10061 19348
rect 10731 19412 10797 19413
rect 10731 19348 10732 19412
rect 10796 19348 10797 19412
rect 10731 19347 10797 19348
rect 9511 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9831 19072
rect 9511 17984 9831 19008
rect 9511 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9831 17984
rect 9511 16896 9831 17920
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9998 7989 10058 19347
rect 10734 9621 10794 19347
rect 11224 18528 11544 19552
rect 11224 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11544 18528
rect 11224 17440 11544 18464
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 12938 21248 13258 21808
rect 12938 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13258 21248
rect 12938 20160 13258 21184
rect 12938 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13258 20160
rect 12938 19072 13258 20096
rect 12938 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13258 19072
rect 12938 17984 13258 19008
rect 12938 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13258 17984
rect 12938 16896 13258 17920
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 11835 15060 11901 15061
rect 11835 14996 11836 15060
rect 11900 14996 11901 15060
rect 11835 14995 11901 14996
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 10731 9620 10797 9621
rect 10731 9556 10732 9620
rect 10796 9556 10797 9620
rect 10731 9555 10797 9556
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 9995 7988 10061 7989
rect 9995 7924 9996 7988
rect 10060 7924 10061 7988
rect 9995 7923 10061 7924
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9259 6220 9325 6221
rect 9259 6156 9260 6220
rect 9324 6156 9325 6220
rect 9259 6155 9325 6156
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9075 4044 9141 4045
rect 9075 3980 9076 4044
rect 9140 3980 9141 4044
rect 9075 3979 9141 3980
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11838 3501 11898 14995
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 11835 3500 11901 3501
rect 11835 3436 11836 3500
rect 11900 3436 11901 3500
rect 11835 3435 11901 3436
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 21792 14971 21808
rect 14651 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14971 21792
rect 14651 20704 14971 21728
rect 14651 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14971 20704
rect 14651 19616 14971 20640
rect 14651 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14971 19616
rect 14651 18528 14971 19552
rect 14651 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14971 18528
rect 14651 17440 14971 18464
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
rect 8891 1868 8957 1869
rect 8891 1804 8892 1868
rect 8956 1804 8957 1868
rect 8891 1803 8957 1804
use sky130_fd_sc_hd__clkbuf_1  _324_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1688980957
transform -1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1688980957
transform -1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1688980957
transform -1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1688980957
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1688980957
transform -1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1688980957
transform -1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform -1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1688980957
transform -1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1688980957
transform -1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1688980957
transform 1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1688980957
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform -1 0 4508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _351_
timestamp 1688980957
transform -1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1688980957
transform -1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1688980957
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1688980957
transform -1 0 4784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1688980957
transform -1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1688980957
transform -1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1688980957
transform -1 0 4140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1688980957
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp 1688980957
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1688980957
transform 1 0 4784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1688980957
transform -1 0 3680 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1688980957
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1688980957
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1688980957
transform -1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1688980957
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1688980957
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1688980957
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1688980957
transform -1 0 13616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1688980957
transform 1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1688980957
transform -1 0 9844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1688980957
transform -1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1688980957
transform -1 0 11224 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1688980957
transform -1 0 11408 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1688980957
transform -1 0 12328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1688980957
transform 1 0 12696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1688980957
transform -1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1688980957
transform 1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1688980957
transform -1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1688980957
transform -1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _391_
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1688980957
transform -1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1688980957
transform -1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _394_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1688980957
transform -1 0 11500 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1688980957
transform -1 0 13892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1688980957
transform 1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1688980957
transform -1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1688980957
transform -1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1688980957
transform -1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1688980957
transform 1 0 12144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1688980957
transform -1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1688980957
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1688980957
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1688980957
transform -1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1688980957
transform -1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1688980957
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _417_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1688980957
transform 1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1688980957
transform -1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1688980957
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1688980957
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1688980957
transform -1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1688980957
transform -1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1688980957
transform -1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _427_
timestamp 1688980957
transform -1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1688980957
transform -1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1688980957
transform -1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1688980957
transform 1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1688980957
transform -1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1688980957
transform -1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1688980957
transform 1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _441_
timestamp 1688980957
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _443_
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1688980957
transform 1 0 9016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1688980957
transform -1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _447_
timestamp 1688980957
transform -1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1688980957
transform -1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _449_
timestamp 1688980957
transform -1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1688980957
transform -1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _452_
timestamp 1688980957
transform -1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1688980957
transform -1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1688980957
transform -1 0 10120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1688980957
transform -1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1688980957
transform 1 0 13064 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1688980957
transform 1 0 13616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1688980957
transform -1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1688980957
transform 1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1688980957
transform 1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1688980957
transform -1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1688980957
transform -1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1688980957
transform -1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1688980957
transform -1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1688980957
transform -1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1688980957
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1688980957
transform -1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1688980957
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _478_
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1688980957
transform -1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1688980957
transform 1 0 6440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1688980957
transform 1 0 4968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1688980957
transform -1 0 1748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1688980957
transform -1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1688980957
transform -1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1688980957
transform 1 0 3864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _489_
timestamp 1688980957
transform -1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1688980957
transform 1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _493_
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1688980957
transform -1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1688980957
transform 1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1688980957
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1688980957
transform -1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _500_
timestamp 1688980957
transform -1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp 1688980957
transform 1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1688980957
transform -1 0 4784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1688980957
transform -1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1688980957
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _511_
timestamp 1688980957
transform -1 0 8280 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _512_
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _513_
timestamp 1688980957
transform -1 0 11316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _514_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _515_
timestamp 1688980957
transform 1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _516_
timestamp 1688980957
transform -1 0 5428 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1688980957
transform -1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _520_
timestamp 1688980957
transform -1 0 8004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _521_
timestamp 1688980957
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _522_
timestamp 1688980957
transform -1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1688980957
transform -1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _524_
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _525_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1688980957
transform -1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _528_
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1688980957
transform -1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1688980957
transform -1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _531_
timestamp 1688980957
transform 1 0 14076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1688980957
transform -1 0 12512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _533_
timestamp 1688980957
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1688980957
transform -1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1688980957
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1688980957
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _537_
timestamp 1688980957
transform -1 0 12420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _538_
timestamp 1688980957
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp 1688980957
transform -1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1688980957
transform 1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1688980957
transform -1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1688980957
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _545_
timestamp 1688980957
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1688980957
transform -1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1688980957
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _550_
timestamp 1688980957
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _551_
timestamp 1688980957
transform -1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1688980957
transform -1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1688980957
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _556_
timestamp 1688980957
transform -1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1688980957
transform -1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1688980957
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _559_
timestamp 1688980957
transform -1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1688980957
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _561_
timestamp 1688980957
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1688980957
transform -1 0 5060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1688980957
transform -1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1688980957
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _566_
timestamp 1688980957
transform -1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1688980957
transform 1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1688980957
transform -1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1688980957
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1688980957
transform -1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1688980957
transform -1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1688980957
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1688980957
transform -1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1688980957
transform -1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _579_
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _581_
timestamp 1688980957
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1688980957
transform -1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1688980957
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1688980957
transform -1 0 6072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _587_
timestamp 1688980957
transform -1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _589_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 1688980957
transform -1 0 6256 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _591_
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1688980957
transform -1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _594_
timestamp 1688980957
transform -1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1688980957
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _597_
timestamp 1688980957
transform -1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1688980957
transform -1 0 3680 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1688980957
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _600_
timestamp 1688980957
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _601_
timestamp 1688980957
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _602_
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _603_
timestamp 1688980957
transform -1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _604_
timestamp 1688980957
transform -1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _605_
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _606_
timestamp 1688980957
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1688980957
transform -1 0 3680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1688980957
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1688980957
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _610_
timestamp 1688980957
transform 1 0 8648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _611_
timestamp 1688980957
transform -1 0 8280 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _612_
timestamp 1688980957
transform -1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _613_
timestamp 1688980957
transform -1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _614_
timestamp 1688980957
transform -1 0 8740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1688980957
transform -1 0 8464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _616_
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _617_
timestamp 1688980957
transform 1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _618_
timestamp 1688980957
transform -1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _619_
timestamp 1688980957
transform -1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _621_
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _622_
timestamp 1688980957
transform -1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _623_
timestamp 1688980957
transform 1 0 3864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _624_
timestamp 1688980957
transform -1 0 2944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1688980957
transform 1 0 2576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1688980957
transform -1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _627_
timestamp 1688980957
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _628_
timestamp 1688980957
transform -1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1688980957
transform -1 0 2576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _630_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1688980957
transform -1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _632_
timestamp 1688980957
transform -1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _633_
timestamp 1688980957
transform 1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1688980957
transform -1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _638_
timestamp 1688980957
transform -1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _639_
timestamp 1688980957
transform -1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _640_
timestamp 1688980957
transform -1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _641_
timestamp 1688980957
transform -1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1688980957
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _643_
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _644_
timestamp 1688980957
transform -1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _645_
timestamp 1688980957
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _646_
timestamp 1688980957
transform -1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _648_
timestamp 1688980957
transform -1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _649_
timestamp 1688980957
transform -1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _650_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _651_
timestamp 1688980957
transform -1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1688980957
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _653_
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _654_
timestamp 1688980957
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _655_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _656_
timestamp 1688980957
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _657_
timestamp 1688980957
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1688980957
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _660_
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1688980957
transform -1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1688980957
transform -1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _665_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _666_
timestamp 1688980957
transform -1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _667_
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _668_
timestamp 1688980957
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1688980957
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _671_
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _673_
timestamp 1688980957
transform 1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1688980957
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _675_
timestamp 1688980957
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _677_
timestamp 1688980957
transform -1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _678_
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _679_
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _680_
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _681_
timestamp 1688980957
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _682_
timestamp 1688980957
transform -1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _683_
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _684_
timestamp 1688980957
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _686_
timestamp 1688980957
transform -1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _687_
timestamp 1688980957
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1688980957
transform -1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1688980957
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _690_
timestamp 1688980957
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1688980957
transform 1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _692_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _693_
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _694_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10672 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _695_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _696_
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _697_
timestamp 1688980957
transform -1 0 11500 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _698_
timestamp 1688980957
transform -1 0 13892 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _699_
timestamp 1688980957
transform 1 0 10948 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _700_
timestamp 1688980957
transform -1 0 13984 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _701_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _702_
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _703_
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _704_
timestamp 1688980957
transform 1 0 2668 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _705_
timestamp 1688980957
transform -1 0 2852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _706_
timestamp 1688980957
transform -1 0 4324 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _707_
timestamp 1688980957
transform -1 0 6992 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _708_
timestamp 1688980957
transform -1 0 4692 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _709_
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _710_
timestamp 1688980957
transform -1 0 6164 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _711_
timestamp 1688980957
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _712_
timestamp 1688980957
transform 1 0 9108 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _713_
timestamp 1688980957
transform -1 0 9200 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _714_
timestamp 1688980957
transform 1 0 6256 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _715_
timestamp 1688980957
transform 1 0 4416 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _716_
timestamp 1688980957
transform -1 0 3128 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _717_
timestamp 1688980957
transform -1 0 2852 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _718_
timestamp 1688980957
transform -1 0 5336 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _719_
timestamp 1688980957
transform 1 0 12420 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _720_
timestamp 1688980957
transform 1 0 2576 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _721_
timestamp 1688980957
transform -1 0 3220 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _722_
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1688980957
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _724_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _725_
timestamp 1688980957
transform 1 0 2208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _726_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _727_
timestamp 1688980957
transform -1 0 11408 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _728_
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _729_
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _730_
timestamp 1688980957
transform 1 0 5152 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _731_
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _732_
timestamp 1688980957
transform -1 0 14444 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _733_
timestamp 1688980957
transform -1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _734_
timestamp 1688980957
transform 1 0 10672 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _735_
timestamp 1688980957
transform -1 0 11316 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _736_
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _737_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _738_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _739_
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _752_
timestamp 1688980957
transform -1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _753_
timestamp 1688980957
transform -1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _754_
timestamp 1688980957
transform 1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _755_
timestamp 1688980957
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _756_
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _757_
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _758_
timestamp 1688980957
transform -1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _759_
timestamp 1688980957
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp 1688980957
transform -1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _761_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _762_
timestamp 1688980957
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp 1688980957
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _764_
timestamp 1688980957
transform 1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _765_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _766_
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _767_
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _768_
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _769_
timestamp 1688980957
transform 1 0 2668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _770_
timestamp 1688980957
transform 1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _771_
timestamp 1688980957
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _772_
timestamp 1688980957
transform -1 0 3128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _773_
timestamp 1688980957
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _774_
timestamp 1688980957
transform -1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _775_
timestamp 1688980957
transform -1 0 7636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11408 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _777_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _778_
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _779_
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _779__83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _780_
timestamp 1688980957
transform -1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _781_
timestamp 1688980957
transform 1 0 6440 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _782_
timestamp 1688980957
transform 1 0 8096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _783_
timestamp 1688980957
transform 1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _784_
timestamp 1688980957
transform 1 0 8188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _785_
timestamp 1688980957
transform 1 0 10120 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _786_
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _787_
timestamp 1688980957
transform 1 0 9292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _788_
timestamp 1688980957
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _789_
timestamp 1688980957
transform -1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _790_
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _791_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _792_
timestamp 1688980957
transform 1 0 7636 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _793_
timestamp 1688980957
transform -1 0 9844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _794_
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _795_
timestamp 1688980957
transform 1 0 10212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _796_
timestamp 1688980957
transform 1 0 13156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _797_
timestamp 1688980957
transform 1 0 10212 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _797__84
timestamp 1688980957
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _798_
timestamp 1688980957
transform 1 0 9200 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _799_
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _800_
timestamp 1688980957
transform -1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _801_
timestamp 1688980957
transform -1 0 14076 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _802_
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _803_
timestamp 1688980957
transform -1 0 12420 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _804_
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _805_
timestamp 1688980957
transform -1 0 12512 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _806_
timestamp 1688980957
transform 1 0 9476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _807_
timestamp 1688980957
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _808_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _809_
timestamp 1688980957
transform -1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _810_
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _811_
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _812_
timestamp 1688980957
transform 1 0 13156 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _813_
timestamp 1688980957
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _814_
timestamp 1688980957
transform -1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _815_
timestamp 1688980957
transform -1 0 13432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _815__85
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _816_
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _817_
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _818_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _819_
timestamp 1688980957
transform -1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _820_
timestamp 1688980957
transform 1 0 9844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _821_
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _822_
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _823_
timestamp 1688980957
transform 1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _824_
timestamp 1688980957
transform 1 0 11960 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _825_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _826_
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _827_
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _828_
timestamp 1688980957
transform 1 0 9844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _829_
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _830_
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _831_
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _832_
timestamp 1688980957
transform 1 0 4140 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _833__86
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _833_
timestamp 1688980957
transform 1 0 1748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _834_
timestamp 1688980957
transform 1 0 2024 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _835_
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _836_
timestamp 1688980957
transform -1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _837_
timestamp 1688980957
transform -1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _838_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _839_
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _840_
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _841_
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _842_
timestamp 1688980957
transform 1 0 1840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _843_
timestamp 1688980957
transform -1 0 2668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _844_
timestamp 1688980957
transform -1 0 4784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _845_
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _846_
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _847_
timestamp 1688980957
transform 1 0 3496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _848_
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _849_
timestamp 1688980957
transform 1 0 3220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _850_
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _851__87
timestamp 1688980957
transform -1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _851_
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _852_
timestamp 1688980957
transform 1 0 2024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _853_
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _854_
timestamp 1688980957
transform -1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _855_
timestamp 1688980957
transform -1 0 7728 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _856_
timestamp 1688980957
transform -1 0 5060 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _857_
timestamp 1688980957
transform 1 0 5060 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _858_
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _859_
timestamp 1688980957
transform -1 0 5888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _860_
timestamp 1688980957
transform 1 0 2116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _861_
timestamp 1688980957
transform 1 0 2116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _862_
timestamp 1688980957
transform -1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _863_
timestamp 1688980957
transform 1 0 5060 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _864_
timestamp 1688980957
transform -1 0 8556 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _865_
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _866_
timestamp 1688980957
transform -1 0 10304 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _867_
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _868_
timestamp 1688980957
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _869_
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _869__88
timestamp 1688980957
transform -1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _870_
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _871_
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _872_
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _873_
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _874_
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _875_
timestamp 1688980957
transform -1 0 10948 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _876_
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _877_
timestamp 1688980957
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _878_
timestamp 1688980957
transform 1 0 9016 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _879_
timestamp 1688980957
transform -1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _880_
timestamp 1688980957
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _881_
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _882_
timestamp 1688980957
transform 1 0 6072 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _883_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _884_
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _885_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _886_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _887__89
timestamp 1688980957
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _887_
timestamp 1688980957
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _888_
timestamp 1688980957
transform -1 0 5980 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _889_
timestamp 1688980957
transform -1 0 5336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _890_
timestamp 1688980957
transform -1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _891_
timestamp 1688980957
transform -1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _892_
timestamp 1688980957
transform 1 0 3312 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _893_
timestamp 1688980957
transform -1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _894_
timestamp 1688980957
transform -1 0 3312 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _895_
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _896_
timestamp 1688980957
transform -1 0 3128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _897_
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _898_
timestamp 1688980957
transform -1 0 6072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _899_
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _900_
timestamp 1688980957
transform -1 0 5060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _901_
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _902_
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _903_
timestamp 1688980957
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _904_
timestamp 1688980957
transform -1 0 5796 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _905__90
timestamp 1688980957
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _905_
timestamp 1688980957
transform 1 0 1840 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _906_
timestamp 1688980957
transform 1 0 2392 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _907_
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _908_
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _909_
timestamp 1688980957
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _910_
timestamp 1688980957
transform 1 0 9016 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _911_
timestamp 1688980957
transform -1 0 5060 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _912_
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _913_
timestamp 1688980957
transform -1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _914_
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _915_
timestamp 1688980957
transform -1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _916_
timestamp 1688980957
transform -1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _917_
timestamp 1688980957
transform -1 0 9016 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _918_
timestamp 1688980957
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _919_
timestamp 1688980957
transform -1 0 11224 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _920_
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _921_
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _922_
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _923__91
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _923_
timestamp 1688980957
transform -1 0 2576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _924_
timestamp 1688980957
transform 1 0 2024 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _925_
timestamp 1688980957
transform 1 0 5152 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _926_
timestamp 1688980957
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _927_
timestamp 1688980957
transform -1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _928_
timestamp 1688980957
transform 1 0 7544 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _929_
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _930_
timestamp 1688980957
transform -1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _931_
timestamp 1688980957
transform 1 0 2300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _932_
timestamp 1688980957
transform 1 0 2024 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _933_
timestamp 1688980957
transform 1 0 5152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _934_
timestamp 1688980957
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _935_
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _936_
timestamp 1688980957
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _937_
timestamp 1688980957
transform -1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _938_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _939__92
timestamp 1688980957
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _939_
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _940_
timestamp 1688980957
transform -1 0 8556 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _941_
timestamp 1688980957
transform 1 0 6164 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _942_
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _943_
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _944_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _945_
timestamp 1688980957
transform 1 0 7636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _946_
timestamp 1688980957
transform -1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _947_
timestamp 1688980957
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _948_
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _949_
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _950_
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _951_
timestamp 1688980957
transform 1 0 7176 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _952_
timestamp 1688980957
transform -1 0 12604 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _953_
timestamp 1688980957
transform -1 0 14076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _954_
timestamp 1688980957
transform 1 0 13248 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _955_
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _955__93
timestamp 1688980957
transform -1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _956_
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _957_
timestamp 1688980957
transform -1 0 13892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _958_
timestamp 1688980957
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _959_
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _960_
timestamp 1688980957
transform -1 0 13248 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _961_
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _962_
timestamp 1688980957
transform -1 0 13800 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _963_
timestamp 1688980957
transform 1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _964_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _965_
timestamp 1688980957
transform 1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _966_
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _967_
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _968_
timestamp 1688980957
transform 1 0 13156 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _969_
timestamp 1688980957
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _970_
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _971__94
timestamp 1688980957
transform -1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _971_
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _972_
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _973_
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _974_
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _975_
timestamp 1688980957
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _976_
timestamp 1688980957
transform 1 0 13156 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _977_
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _978_
timestamp 1688980957
transform 1 0 12420 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _979_
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _980_
timestamp 1688980957
transform 1 0 11868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _981_
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _982_
timestamp 1688980957
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _983_
timestamp 1688980957
transform 1 0 5888 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1688980957
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1688980957
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_108
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_13
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_52
timestamp 1688980957
transform 1 0 5888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_65
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_88
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 1688980957
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_103
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_13
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_34
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_64
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_10
timestamp 1688980957
transform 1 0 2024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_68
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_72
timestamp 1688980957
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_80
timestamp 1688980957
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_104
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_144
timestamp 1688980957
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_13
timestamp 1688980957
transform 1 0 2300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_22
timestamp 1688980957
transform 1 0 3128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_50
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_60
timestamp 1688980957
transform 1 0 6624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_14
timestamp 1688980957
transform 1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_24
timestamp 1688980957
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_102
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_128
timestamp 1688980957
transform 1 0 12880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_26
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_83
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_13
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_22
timestamp 1688980957
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_54
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_63
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_110
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_144
timestamp 1688980957
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_44
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_68
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_144
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_96
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_144
timestamp 1688980957
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_13
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_63
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_82 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_88
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_95
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_130
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_32
timestamp 1688980957
transform 1 0 4048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_96
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_103
timestamp 1688980957
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_144
timestamp 1688980957
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_24
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_34
timestamp 1688980957
transform 1 0 4232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_60
timestamp 1688980957
transform 1 0 6624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_77
timestamp 1688980957
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_90
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_98
timestamp 1688980957
transform 1 0 10120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_118
timestamp 1688980957
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_40
timestamp 1688980957
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_107
timestamp 1688980957
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_112
timestamp 1688980957
transform 1 0 11408 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_116
timestamp 1688980957
transform 1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_144
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_8
timestamp 1688980957
transform 1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_24
timestamp 1688980957
transform 1 0 3312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_37
timestamp 1688980957
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_50
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_104
timestamp 1688980957
transform 1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_132
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_10
timestamp 1688980957
transform 1 0 2024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_46
timestamp 1688980957
transform 1 0 5336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_66
timestamp 1688980957
transform 1 0 7176 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_123
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_60
timestamp 1688980957
transform 1 0 6624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_119
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_127
timestamp 1688980957
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_145
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_6
timestamp 1688980957
transform 1 0 1656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_18
timestamp 1688980957
transform 1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_52
timestamp 1688980957
transform 1 0 5888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_56
timestamp 1688980957
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_94
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_98
timestamp 1688980957
transform 1 0 10120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_126
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_144
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_14
timestamp 1688980957
transform 1 0 2392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_42
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_123
timestamp 1688980957
transform 1 0 12420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_127
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_139
timestamp 1688980957
transform 1 0 13892 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_8
timestamp 1688980957
transform 1 0 1840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_18
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_40
timestamp 1688980957
transform 1 0 4784 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_136
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_144
timestamp 1688980957
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_16
timestamp 1688980957
transform 1 0 2576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_35
timestamp 1688980957
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_68
timestamp 1688980957
transform 1 0 7360 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_116
timestamp 1688980957
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_20
timestamp 1688980957
transform 1 0 2944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_111
timestamp 1688980957
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_144
timestamp 1688980957
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_35
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_68
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_79
timestamp 1688980957
transform 1 0 8372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_101
timestamp 1688980957
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_140
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_43
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_47
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_88
timestamp 1688980957
transform 1 0 9200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_113
timestamp 1688980957
transform 1 0 11500 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_119
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_144
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_17
timestamp 1688980957
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_74
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_84
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_107
timestamp 1688980957
transform 1 0 10948 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_140
timestamp 1688980957
transform 1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_70
timestamp 1688980957
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_80
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_112
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_144
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_49
timestamp 1688980957
transform 1 0 5612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_73
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_88
timestamp 1688980957
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_116
timestamp 1688980957
transform 1 0 11776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_9
timestamp 1688980957
transform 1 0 1932 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_33
timestamp 1688980957
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_42
timestamp 1688980957
transform 1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_61
timestamp 1688980957
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1688980957
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_115
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_44
timestamp 1688980957
transform 1 0 5152 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_80
timestamp 1688980957
transform 1 0 8464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_85
timestamp 1688980957
transform 1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_95
timestamp 1688980957
transform 1 0 9844 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_116
timestamp 1688980957
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_124
timestamp 1688980957
transform 1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_6
timestamp 1688980957
transform 1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_16
timestamp 1688980957
transform 1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_126
timestamp 1688980957
transform 1 0 12696 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_144
timestamp 1688980957
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_12
timestamp 1688980957
transform 1 0 2208 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_36
timestamp 1688980957
transform 1 0 4416 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_86
timestamp 1688980957
transform 1 0 9016 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_94
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_106
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_124
timestamp 1688980957
transform 1 0 12512 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_144
timestamp 1688980957
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_23
timestamp 1688980957
transform 1 0 3220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_51
timestamp 1688980957
transform 1 0 5796 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_144
timestamp 1688980957
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_82
timestamp 1688980957
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_16
timestamp 1688980957
transform 1 0 2576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_129
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_144
timestamp 1688980957
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_60
timestamp 1688980957
transform 1 0 6624 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_77
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_85
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_101
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_122
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_139
timestamp 1688980957
transform 1 0 13892 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_144
timestamp 1688980957
transform 1 0 14352 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 6992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 4140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 4968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 11040 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 11684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 8188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 5520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 11040 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 3588 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 2392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 3680 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 12236 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 13156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 10488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 5980 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 7360 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform -1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform -1 0 14536 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 12420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1688980957
transform -1 0 3496 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform -1 0 4048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 2668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform -1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform -1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform -1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform -1 0 10304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 1688980957
transform -1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1688980957
transform -1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output49
timestamp 1688980957
transform -1 0 1932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 1688980957
transform -1 0 1932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 1688980957
transform -1 0 1932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 1688980957
transform -1 0 1932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output53
timestamp 1688980957
transform -1 0 2300 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1688980957
transform -1 0 1932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform -1 0 2852 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1688980957
transform 1 0 14168 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1688980957
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 13984 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform 1 0 13432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 7636 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform -1 0 11408 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
<< labels >>
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 0 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
flabel metal3 s 15200 22040 16000 22160 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 15200 23128 16000 23248 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 5 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 6 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 7 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 8 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 9 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 10 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 11 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 12 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 13 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 14 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 15 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 16 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 17 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 18 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 19 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 20 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 21 nsew signal tristate
flabel metal3 s 15200 280 16000 400 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 22 nsew signal input
flabel metal3 s 15200 1368 16000 1488 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 23 nsew signal input
flabel metal3 s 15200 2456 16000 2576 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 24 nsew signal input
flabel metal3 s 15200 3544 16000 3664 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 25 nsew signal input
flabel metal3 s 15200 4632 16000 4752 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 26 nsew signal input
flabel metal3 s 15200 5720 16000 5840 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 27 nsew signal input
flabel metal3 s 15200 6808 16000 6928 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 28 nsew signal input
flabel metal3 s 15200 7896 16000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 29 nsew signal input
flabel metal3 s 15200 8984 16000 9104 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 30 nsew signal input
flabel metal3 s 15200 10072 16000 10192 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal3 s 15200 11160 16000 11280 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 32 nsew signal tristate
flabel metal3 s 15200 12248 16000 12368 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 33 nsew signal tristate
flabel metal3 s 15200 13336 16000 13456 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 34 nsew signal tristate
flabel metal3 s 15200 14424 16000 14544 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 35 nsew signal tristate
flabel metal3 s 15200 15512 16000 15632 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 36 nsew signal tristate
flabel metal3 s 15200 16600 16000 16720 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 37 nsew signal tristate
flabel metal3 s 15200 17688 16000 17808 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 38 nsew signal tristate
flabel metal3 s 15200 18776 16000 18896 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 39 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 40 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 41 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 42 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 43 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 44 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 45 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 46 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 47 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 48 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 49 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 50 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 51 nsew signal tristate
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 52 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 53 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 54 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 55 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 56 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 57 nsew signal tristate
flabel metal2 s 938 23200 994 24000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 58 nsew signal input
flabel metal2 s 1674 23200 1730 24000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 59 nsew signal input
flabel metal2 s 2410 23200 2466 24000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 60 nsew signal input
flabel metal2 s 3146 23200 3202 24000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 61 nsew signal input
flabel metal2 s 3882 23200 3938 24000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 62 nsew signal input
flabel metal2 s 4618 23200 4674 24000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 63 nsew signal input
flabel metal2 s 5354 23200 5410 24000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 64 nsew signal input
flabel metal2 s 6090 23200 6146 24000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 65 nsew signal input
flabel metal2 s 6826 23200 6882 24000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 66 nsew signal input
flabel metal2 s 7562 23200 7618 24000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 67 nsew signal tristate
flabel metal2 s 8298 23200 8354 24000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 68 nsew signal tristate
flabel metal2 s 9034 23200 9090 24000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 69 nsew signal tristate
flabel metal2 s 9770 23200 9826 24000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 70 nsew signal tristate
flabel metal2 s 10506 23200 10562 24000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 71 nsew signal tristate
flabel metal2 s 11242 23200 11298 24000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 72 nsew signal tristate
flabel metal2 s 11978 23200 12034 24000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 73 nsew signal tristate
flabel metal2 s 12714 23200 12770 24000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 74 nsew signal tristate
flabel metal2 s 13450 23200 13506 24000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 75 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 76 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 77 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 prog_clk
port 78 nsew signal input
flabel metal3 s 15200 19864 16000 19984 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 79 nsew signal input
flabel metal3 s 15200 20952 16000 21072 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 80 nsew signal input
flabel metal2 s 14186 23200 14242 24000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 81 nsew signal input
flabel metal2 s 14922 23200 14978 24000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 82 nsew signal input
flabel metal4 s 2657 2128 2977 21808 0 FreeSans 1920 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 6084 2128 6404 21808 0 FreeSans 1920 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 9511 2128 9831 21808 0 FreeSans 1920 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 12938 2128 13258 21808 0 FreeSans 1920 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 4370 2128 4690 21808 0 FreeSans 1920 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 21808 0 FreeSans 1920 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 21808 0 FreeSans 1920 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 21808 0 FreeSans 1920 90 0 0 vss
port 84 nsew ground bidirectional
rlabel metal1 7958 21216 7958 21216 0 vdd
rlabel via1 8037 21760 8037 21760 0 vss
rlabel metal1 11684 13906 11684 13906 0 _000_
rlabel metal1 5336 20910 5336 20910 0 _001_
rlabel metal1 7222 19448 7222 19448 0 _002_
rlabel metal1 8602 17782 8602 17782 0 _003_
rlabel metal1 12604 12410 12604 12410 0 _004_
rlabel metal1 9430 17646 9430 17646 0 _005_
rlabel metal1 11316 17646 11316 17646 0 _006_
rlabel metal1 13386 18632 13386 18632 0 _007_
rlabel metal1 10718 19856 10718 19856 0 _008_
rlabel metal1 11086 17680 11086 17680 0 _009_
rlabel metal1 12926 9656 12926 9656 0 _010_
rlabel metal2 14122 5117 14122 5117 0 _011_
rlabel metal1 13110 7480 13110 7480 0 _012_
rlabel metal1 8878 4590 8878 4590 0 _013_
rlabel metal1 10902 5338 10902 5338 0 _014_
rlabel metal1 14306 6732 14306 6732 0 _015_
rlabel metal1 11454 4794 11454 4794 0 _016_
rlabel metal1 5060 18734 5060 18734 0 _017_
rlabel metal1 7268 17306 7268 17306 0 _018_
rlabel metal1 8556 10234 8556 10234 0 _019_
rlabel metal2 6578 9078 6578 9078 0 _020_
rlabel metal1 10626 10608 10626 10608 0 _021_
rlabel metal1 7498 7446 7498 7446 0 _022_
rlabel metal1 9338 9588 9338 9588 0 _023_
rlabel metal1 7360 8466 7360 8466 0 _024_
rlabel metal1 8234 5678 8234 5678 0 _025_
rlabel metal1 6210 7378 6210 7378 0 _026_
rlabel metal1 5014 10132 5014 10132 0 _027_
rlabel metal1 4600 9554 4600 9554 0 _028_
rlabel metal1 6486 10574 6486 10574 0 _029_
rlabel metal1 1656 10234 1656 10234 0 _030_
rlabel metal1 3726 9486 3726 9486 0 _031_
rlabel metal1 2806 8976 2806 8976 0 _032_
rlabel viali 8326 18735 8326 18735 0 _033_
rlabel metal1 8234 19482 8234 19482 0 _034_
rlabel metal1 8188 18258 8188 18258 0 _035_
rlabel metal2 4186 19380 4186 19380 0 _036_
rlabel metal1 5566 16524 5566 16524 0 _037_
rlabel metal1 2714 20944 2714 20944 0 _038_
rlabel metal1 1794 18938 1794 18938 0 _039_
rlabel metal2 4002 17476 4002 17476 0 _040_
rlabel metal2 2254 20740 2254 20740 0 _041_
rlabel metal1 3036 11730 3036 11730 0 _042_
rlabel metal1 4140 8466 4140 8466 0 _043_
rlabel metal1 3956 4250 3956 4250 0 _044_
rlabel metal1 2254 6426 2254 6426 0 _045_
rlabel metal1 3864 6290 3864 6290 0 _046_
rlabel metal2 2438 8262 2438 8262 0 _047_
rlabel metal1 4968 6154 4968 6154 0 _048_
rlabel metal1 1702 4590 1702 4590 0 _049_
rlabel metal1 4324 10166 4324 10166 0 _050_
rlabel metal1 5336 17306 5336 17306 0 _051_
rlabel metal1 7682 4556 7682 4556 0 _052_
rlabel metal1 7084 4590 7084 4590 0 _053_
rlabel metal1 9844 2618 9844 2618 0 _054_
rlabel metal1 6624 3026 6624 3026 0 _055_
rlabel metal1 11224 2414 11224 2414 0 _056_
rlabel metal1 7912 5678 7912 5678 0 _057_
rlabel metal1 9940 4586 9940 4586 0 _058_
rlabel metal1 8556 5202 8556 5202 0 _059_
rlabel metal1 4968 12818 4968 12818 0 _060_
rlabel metal1 5566 12818 5566 12818 0 _061_
rlabel metal1 6808 13906 6808 13906 0 _062_
rlabel metal2 1886 3978 1886 3978 0 _063_
rlabel metal1 2576 3026 2576 3026 0 _064_
rlabel metal1 4600 3366 4600 3366 0 _065_
rlabel metal1 1794 11152 1794 11152 0 _066_
rlabel metal1 5750 4624 5750 4624 0 _067_
rlabel metal1 6118 8602 6118 8602 0 _068_
rlabel metal1 3312 12818 3312 12818 0 _069_
rlabel metal1 4278 14246 4278 14246 0 _070_
rlabel metal1 6026 12886 6026 12886 0 _071_
rlabel metal1 3588 16218 3588 16218 0 _072_
rlabel metal1 1702 17306 1702 17306 0 _073_
rlabel metal1 5106 15470 5106 15470 0 _074_
rlabel metal1 2162 12682 2162 12682 0 _075_
rlabel metal1 1978 15538 1978 15538 0 _076_
rlabel metal1 1518 14042 1518 14042 0 _077_
rlabel metal1 9844 17646 9844 17646 0 _078_
rlabel metal2 12282 18734 12282 18734 0 _079_
rlabel metal2 12282 21114 12282 21114 0 _080_
rlabel metal1 14306 16490 14306 16490 0 _081_
rlabel metal2 12374 16762 12374 16762 0 _082_
rlabel metal1 13938 13940 13938 13940 0 _083_
rlabel metal1 11316 12954 11316 12954 0 _084_
rlabel metal1 13938 16150 13938 16150 0 _085_
rlabel metal1 13110 13260 13110 13260 0 _086_
rlabel metal1 13800 13294 13800 13294 0 _087_
rlabel metal1 14260 7378 14260 7378 0 _088_
rlabel metal1 14214 7854 14214 7854 0 _089_
rlabel metal2 12558 8772 12558 8772 0 _090_
rlabel metal2 11178 10438 11178 10438 0 _091_
rlabel metal1 11408 8466 11408 8466 0 _092_
rlabel metal1 9062 7854 9062 7854 0 _093_
rlabel metal1 10304 8942 10304 8942 0 _094_
rlabel metal1 9430 9690 9430 9690 0 _095_
rlabel metal1 8648 17170 8648 17170 0 _096_
rlabel metal1 8786 14382 8786 14382 0 _097_
rlabel metal1 8188 16558 8188 16558 0 _098_
rlabel metal1 11500 11730 11500 11730 0 _099_
rlabel metal1 9246 14416 9246 14416 0 _100_
rlabel metal1 5566 15436 5566 15436 0 _101_
rlabel metal1 10074 13498 10074 13498 0 _102_
rlabel metal2 9890 12410 9890 12410 0 _103_
rlabel metal1 11546 14008 11546 14008 0 _104_
rlabel metal1 10626 13906 10626 13906 0 _105_
rlabel metal2 9062 15028 9062 15028 0 _106_
rlabel metal1 10212 12342 10212 12342 0 _107_
rlabel metal1 10902 11220 10902 11220 0 _108_
rlabel metal1 6210 15674 6210 15674 0 _109_
rlabel metal1 8372 14586 8372 14586 0 _110_
rlabel metal1 7636 15538 7636 15538 0 _111_
rlabel metal1 8694 17102 8694 17102 0 _112_
rlabel metal1 10672 15402 10672 15402 0 _113_
rlabel metal1 10350 13362 10350 13362 0 _114_
rlabel metal1 10028 14586 10028 14586 0 _115_
rlabel metal1 11316 12886 11316 12886 0 _116_
rlabel metal2 11914 12002 11914 12002 0 _117_
rlabel metal1 6256 15538 6256 15538 0 _118_
rlabel metal1 8924 16626 8924 16626 0 _119_
rlabel metal1 7958 14586 7958 14586 0 _120_
rlabel metal1 9292 20366 9292 20366 0 _121_
rlabel metal1 11040 8602 11040 8602 0 _122_
rlabel metal1 10488 9146 10488 9146 0 _123_
rlabel metal1 13386 9078 13386 9078 0 _124_
rlabel metal1 10442 9996 10442 9996 0 _125_
rlabel metal1 9292 7922 9292 7922 0 _126_
rlabel metal1 12466 10540 12466 10540 0 _127_
rlabel metal1 14076 7174 14076 7174 0 _128_
rlabel metal1 13984 7378 13984 7378 0 _129_
rlabel metal1 13984 13158 13984 13158 0 _130_
rlabel metal1 12282 8058 12282 8058 0 _131_
rlabel metal1 10580 8398 10580 8398 0 _132_
rlabel metal1 12466 8466 12466 8466 0 _133_
rlabel metal1 9798 10098 9798 10098 0 _134_
rlabel metal1 9614 6834 9614 6834 0 _135_
rlabel metal1 11546 10234 11546 10234 0 _136_
rlabel metal1 14214 9452 14214 9452 0 _137_
rlabel metal1 13156 8466 13156 8466 0 _138_
rlabel metal1 13938 11764 13938 11764 0 _139_
rlabel metal1 13570 14042 13570 14042 0 _140_
rlabel metal1 12696 14450 12696 14450 0 _141_
rlabel metal2 13846 18938 13846 18938 0 _142_
rlabel metal2 13294 13668 13294 13668 0 _143_
rlabel metal1 11684 14450 11684 14450 0 _144_
rlabel metal1 12788 16762 12788 16762 0 _145_
rlabel metal1 11730 19244 11730 19244 0 _146_
rlabel metal1 11730 20876 11730 20876 0 _147_
rlabel metal1 10028 17850 10028 17850 0 _148_
rlabel metal1 13386 15368 13386 15368 0 _149_
rlabel metal1 12466 15538 12466 15538 0 _150_
rlabel metal2 13478 18020 13478 18020 0 _151_
rlabel metal1 12788 13498 12788 13498 0 _152_
rlabel metal1 12052 14926 12052 14926 0 _153_
rlabel metal2 12190 16796 12190 16796 0 _154_
rlabel metal1 11914 18394 11914 18394 0 _155_
rlabel metal1 10580 20366 10580 20366 0 _156_
rlabel metal1 11086 18802 11086 18802 0 _157_
rlabel metal2 4830 15912 4830 15912 0 _158_
rlabel metal1 2323 15606 2323 15606 0 _159_
rlabel metal1 4370 16558 4370 16558 0 _160_
rlabel metal1 1794 14926 1794 14926 0 _161_
rlabel metal1 2346 13362 2346 13362 0 _162_
rlabel metal1 3082 16524 3082 16524 0 _163_
rlabel metal1 5014 13906 5014 13906 0 _164_
rlabel metal1 6532 12954 6532 12954 0 _165_
rlabel metal1 3726 12954 3726 12954 0 _166_
rlabel metal1 5658 16184 5658 16184 0 _167_
rlabel metal1 3036 14994 3036 14994 0 _168_
rlabel metal1 3772 16014 3772 16014 0 _169_
rlabel metal1 1886 13498 1886 13498 0 _170_
rlabel metal1 2438 15980 2438 15980 0 _171_
rlabel metal1 4140 15538 4140 15538 0 _172_
rlabel metal1 4278 14518 4278 14518 0 _173_
rlabel metal1 5750 13940 5750 13940 0 _174_
rlabel metal1 3680 12750 3680 12750 0 _175_
rlabel metal1 4646 4182 4646 4182 0 _176_
rlabel metal1 3496 4046 3496 4046 0 _177_
rlabel metal1 3864 2414 3864 2414 0 _178_
rlabel metal1 3128 4658 3128 4658 0 _179_
rlabel metal1 2116 11322 2116 11322 0 _180_
rlabel metal1 6026 2346 6026 2346 0 _181_
rlabel metal1 6624 12886 6624 12886 0 _182_
rlabel metal1 7406 14042 7406 14042 0 _183_
rlabel metal1 5014 12274 5014 12274 0 _184_
rlabel metal1 5014 3094 5014 3094 0 _185_
rlabel metal2 4140 10268 4140 10268 0 _186_
rlabel metal1 5658 4148 5658 4148 0 _187_
rlabel metal1 4324 10438 4324 10438 0 _188_
rlabel metal1 2116 11186 2116 11186 0 _189_
rlabel metal1 6762 2482 6762 2482 0 _190_
rlabel metal1 5198 13158 5198 13158 0 _191_
rlabel metal1 7866 12274 7866 12274 0 _192_
rlabel metal1 4324 12342 4324 12342 0 _193_
rlabel metal1 10074 2312 10074 2312 0 _194_
rlabel metal1 10304 4794 10304 4794 0 _195_
rlabel metal1 12972 2890 12972 2890 0 _196_
rlabel metal1 9246 5338 9246 5338 0 _197_
rlabel metal1 8648 5882 8648 5882 0 _198_
rlabel metal1 7130 2482 7130 2482 0 _199_
rlabel metal1 7590 4794 7590 4794 0 _200_
rlabel metal1 6900 4794 6900 4794 0 _201_
rlabel metal1 5106 18360 5106 18360 0 _202_
rlabel metal1 10902 4182 10902 4182 0 _203_
rlabel metal1 9752 4794 9752 4794 0 _204_
rlabel metal2 9706 4165 9706 4165 0 _205_
rlabel metal1 8970 5746 8970 5746 0 _206_
rlabel metal1 7774 6188 7774 6188 0 _207_
rlabel metal1 7912 3706 7912 3706 0 _208_
rlabel metal1 7406 5882 7406 5882 0 _209_
rlabel metal1 6394 4658 6394 4658 0 _210_
rlabel metal1 6348 17306 6348 17306 0 _211_
rlabel metal2 2530 7888 2530 7888 0 _212_
rlabel metal1 2116 4794 2116 4794 0 _213_
rlabel metal1 4002 6732 4002 6732 0 _214_
rlabel metal1 3634 5304 3634 5304 0 _215_
rlabel metal1 5750 7276 5750 7276 0 _216_
rlabel metal1 4600 6426 4600 6426 0 _217_
rlabel metal1 4692 8602 4692 8602 0 _218_
rlabel metal1 4738 5134 4738 5134 0 _219_
rlabel metal1 3542 11628 3542 11628 0 _220_
rlabel metal1 4370 7752 4370 7752 0 _221_
rlabel metal1 1886 5848 1886 5848 0 _222_
rlabel metal1 4646 7412 4646 7412 0 _223_
rlabel metal1 3220 5134 3220 5134 0 _224_
rlabel metal1 5014 8466 5014 8466 0 _225_
rlabel metal1 4738 6358 4738 6358 0 _226_
rlabel metal1 3726 8058 3726 8058 0 _227_
rlabel metal1 5014 11118 5014 11118 0 _228_
rlabel metal1 3680 11866 3680 11866 0 _229_
rlabel metal1 3588 19414 3588 19414 0 _230_
rlabel metal2 3818 17204 3818 17204 0 _231_
rlabel metal1 5566 19754 5566 19754 0 _232_
rlabel metal1 2208 18802 2208 18802 0 _233_
rlabel metal1 2392 18258 2392 18258 0 _234_
rlabel metal1 6578 16660 6578 16660 0 _235_
rlabel metal1 9154 19924 9154 19924 0 _236_
rlabel metal1 8096 17646 8096 17646 0 _237_
rlabel metal1 9062 18802 9062 18802 0 _238_
rlabel metal2 4830 20043 4830 20043 0 _239_
rlabel metal1 2898 19346 2898 19346 0 _240_
rlabel metal1 5014 19312 5014 19312 0 _241_
rlabel metal1 1748 18258 1748 18258 0 _242_
rlabel metal2 3266 17884 3266 17884 0 _243_
rlabel metal1 7544 16082 7544 16082 0 _244_
rlabel metal1 8786 19312 8786 19312 0 _245_
rlabel metal1 8234 20026 8234 20026 0 _246_
rlabel metal1 9890 18394 9890 18394 0 _247_
rlabel metal1 6808 10710 6808 10710 0 _248_
rlabel metal1 3956 9690 3956 9690 0 _249_
rlabel metal1 5474 10132 5474 10132 0 _250_
rlabel metal1 2484 8942 2484 8942 0 _251_
rlabel metal1 1932 10778 1932 10778 0 _252_
rlabel metal1 5382 9452 5382 9452 0 _253_
rlabel metal1 6440 6834 6440 6834 0 _254_
rlabel metal1 6854 5746 6854 5746 0 _255_
rlabel metal1 7314 9690 7314 9690 0 _256_
rlabel metal1 3358 10778 3358 10778 0 _257_
rlabel metal1 6256 9690 6256 9690 0 _258_
rlabel metal1 2852 9486 2852 9486 0 _259_
rlabel metal1 2208 10574 2208 10574 0 _260_
rlabel metal1 5198 9010 5198 9010 0 _261_
rlabel metal1 7038 5882 7038 5882 0 _262_
rlabel metal1 5888 5338 5888 5338 0 _263_
rlabel metal1 9798 10710 9798 10710 0 _264_
rlabel metal1 8878 9452 8878 9452 0 _265_
rlabel metal1 8050 9554 8050 9554 0 _266_
rlabel metal1 8142 8364 8142 8364 0 _267_
rlabel metal2 8326 7004 8326 7004 0 _268_
rlabel metal1 6440 9010 6440 9010 0 _269_
rlabel metal1 7268 17714 7268 17714 0 _270_
rlabel metal1 5566 18836 5566 18836 0 _271_
rlabel metal1 8050 11526 8050 11526 0 _272_
rlabel metal1 8096 9010 8096 9010 0 _273_
rlabel metal1 7222 10132 7222 10132 0 _274_
rlabel metal1 8050 8534 8050 8534 0 _275_
rlabel metal1 7130 7514 7130 7514 0 _276_
rlabel metal1 7130 8908 7130 8908 0 _277_
rlabel metal1 6854 17170 6854 17170 0 _278_
rlabel metal1 7406 18326 7406 18326 0 _279_
rlabel metal1 8878 4794 8878 4794 0 _280_
rlabel metal1 13892 5202 13892 5202 0 _281_
rlabel via2 13478 6307 13478 6307 0 _282_
rlabel metal1 11914 5338 11914 5338 0 _283_
rlabel metal1 11040 5746 11040 5746 0 _284_
rlabel metal1 13064 6834 13064 6834 0 _285_
rlabel metal2 14122 10676 14122 10676 0 _286_
rlabel metal2 10902 18020 10902 18020 0 _287_
rlabel metal1 8280 4794 8280 4794 0 _288_
rlabel metal1 13616 2618 13616 2618 0 _289_
rlabel metal1 13892 4794 13892 4794 0 _290_
rlabel metal1 12420 6766 12420 6766 0 _291_
rlabel metal2 11730 6052 11730 6052 0 _292_
rlabel metal1 12834 7514 12834 7514 0 _293_
rlabel metal1 11822 11186 11822 11186 0 _294_
rlabel metal1 10442 17850 10442 17850 0 _295_
rlabel metal1 13386 19720 13386 19720 0 _296_
rlabel metal1 13018 19890 13018 19890 0 _297_
rlabel metal1 13570 19210 13570 19210 0 _298_
rlabel metal2 10902 20570 10902 20570 0 _299_
rlabel metal1 12627 17714 12627 17714 0 _300_
rlabel metal1 12926 11730 12926 11730 0 _301_
rlabel metal1 7452 20910 7452 20910 0 _302_
rlabel metal1 5658 20434 5658 20434 0 _303_
rlabel metal2 12834 19295 12834 19295 0 _304_
rlabel metal1 12558 19244 12558 19244 0 _305_
rlabel metal1 12650 19448 12650 19448 0 _306_
rlabel metal1 12052 19482 12052 19482 0 _307_
rlabel metal2 12098 17884 12098 17884 0 _308_
rlabel metal1 12834 11866 12834 11866 0 _309_
rlabel metal1 7452 20978 7452 20978 0 _310_
rlabel metal2 6118 19652 6118 19652 0 _311_
rlabel metal2 7958 823 7958 823 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 7222 1299 7222 1299 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 10672 22134 10672 22134 0 ccff_head
rlabel metal3 14636 23188 14636 23188 0 ccff_tail
rlabel metal3 751 2516 751 2516 0 chanx_left_in[0]
rlabel metal3 820 3604 820 3604 0 chanx_left_in[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_in[2]
rlabel metal3 1004 5780 1004 5780 0 chanx_left_in[3]
rlabel metal3 820 6868 820 6868 0 chanx_left_in[4]
rlabel metal3 1050 7956 1050 7956 0 chanx_left_in[5]
rlabel metal3 820 9044 820 9044 0 chanx_left_in[6]
rlabel metal3 1004 10132 1004 10132 0 chanx_left_in[7]
rlabel metal3 1050 11220 1050 11220 0 chanx_left_in[8]
rlabel metal3 820 14484 820 14484 0 chanx_left_out[0]
rlabel metal3 820 15572 820 15572 0 chanx_left_out[1]
rlabel metal3 820 16660 820 16660 0 chanx_left_out[2]
rlabel metal3 820 17748 820 17748 0 chanx_left_out[3]
rlabel metal3 820 18836 820 18836 0 chanx_left_out[4]
rlabel metal3 820 19924 820 19924 0 chanx_left_out[5]
rlabel metal3 820 21012 820 21012 0 chanx_left_out[6]
rlabel metal3 1096 22100 1096 22100 0 chanx_left_out[7]
rlabel metal3 1740 23188 1740 23188 0 chanx_left_out[8]
rlabel metal2 12052 340 12052 340 0 chanx_right_in[0]
rlabel metal3 13808 1428 13808 1428 0 chanx_right_in[1]
rlabel metal2 11868 2652 11868 2652 0 chanx_right_in[2]
rlabel metal1 13202 3536 13202 3536 0 chanx_right_in[3]
rlabel metal1 14628 5202 14628 5202 0 chanx_right_in[4]
rlabel metal2 14490 4403 14490 4403 0 chanx_right_in[5]
rlabel viali 13018 7377 13018 7377 0 chanx_right_in[6]
rlabel metal1 13110 6766 13110 6766 0 chanx_right_in[7]
rlabel metal1 12466 9588 12466 9588 0 chanx_right_in[8]
rlabel metal2 14398 10285 14398 10285 0 chanx_right_out[0]
rlabel metal1 14398 11254 14398 11254 0 chanx_right_out[1]
rlabel metal1 14674 12614 14674 12614 0 chanx_right_out[2]
rlabel metal1 14444 13702 14444 13702 0 chanx_right_out[3]
rlabel metal2 14398 14637 14398 14637 0 chanx_right_out[4]
rlabel metal2 14398 15725 14398 15725 0 chanx_right_out[5]
rlabel metal2 14398 16813 14398 16813 0 chanx_right_out[6]
rlabel metal1 14444 18054 14444 18054 0 chanx_right_out[7]
rlabel metal2 13938 18581 13938 18581 0 chanx_right_out[8]
rlabel metal2 598 1588 598 1588 0 chany_bottom_in[0]
rlabel metal2 1334 1554 1334 1554 0 chany_bottom_in[1]
rlabel metal2 2070 959 2070 959 0 chany_bottom_in[2]
rlabel metal2 2806 1384 2806 1384 0 chany_bottom_in[3]
rlabel metal2 3542 1761 3542 1761 0 chany_bottom_in[4]
rlabel metal1 4554 2822 4554 2822 0 chany_bottom_in[5]
rlabel metal2 5014 1554 5014 1554 0 chany_bottom_in[6]
rlabel metal1 6440 3910 6440 3910 0 chany_bottom_in[7]
rlabel metal2 6486 1299 6486 1299 0 chany_bottom_in[8]
rlabel metal2 8694 959 8694 959 0 chany_bottom_out[0]
rlabel metal1 9476 2822 9476 2822 0 chany_bottom_out[1]
rlabel metal2 10166 959 10166 959 0 chany_bottom_out[2]
rlabel metal2 10902 1792 10902 1792 0 chany_bottom_out[3]
rlabel metal2 11638 823 11638 823 0 chany_bottom_out[4]
rlabel metal2 12374 1520 12374 1520 0 chany_bottom_out[5]
rlabel metal2 13110 1520 13110 1520 0 chany_bottom_out[6]
rlabel metal1 14030 6086 14030 6086 0 chany_bottom_out[7]
rlabel metal1 14030 2822 14030 2822 0 chany_bottom_out[8]
rlabel metal2 1065 23324 1065 23324 0 chany_top_in[0]
rlabel metal2 1978 21505 1978 21505 0 chany_top_in[1]
rlabel metal2 2438 21940 2438 21940 0 chany_top_in[2]
rlabel metal2 3266 17612 3266 17612 0 chany_top_in[3]
rlabel metal1 4370 20026 4370 20026 0 chany_top_in[4]
rlabel metal2 4416 23324 4416 23324 0 chany_top_in[5]
rlabel metal2 5382 22695 5382 22695 0 chany_top_in[6]
rlabel metal1 5244 21454 5244 21454 0 chany_top_in[7]
rlabel metal1 6302 21590 6302 21590 0 chany_top_in[8]
rlabel metal2 7643 23324 7643 23324 0 chany_top_out[0]
rlabel metal2 8326 22695 8326 22695 0 chany_top_out[1]
rlabel metal1 9200 21658 9200 21658 0 chany_top_out[2]
rlabel metal1 9936 21658 9936 21658 0 chany_top_out[3]
rlabel metal2 10679 23324 10679 23324 0 chany_top_out[4]
rlabel metal2 11270 22695 11270 22695 0 chany_top_out[5]
rlabel metal1 11684 20026 11684 20026 0 chany_top_out[6]
rlabel metal1 12880 18938 12880 18938 0 chany_top_out[7]
rlabel metal1 12834 20264 12834 20264 0 chany_top_out[8]
rlabel metal1 8050 7446 8050 7446 0 clknet_0_prog_clk
rlabel metal2 2254 8942 2254 8942 0 clknet_2_0__leaf_prog_clk
rlabel metal1 13478 4114 13478 4114 0 clknet_2_1__leaf_prog_clk
rlabel metal1 2622 20468 2622 20468 0 clknet_2_2__leaf_prog_clk
rlabel metal2 13846 15572 13846 15572 0 clknet_2_3__leaf_prog_clk
rlabel metal3 820 12308 820 12308 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1326 1428 1326 1428 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 8786 11526 8786 11526 0 mem_bottom_track_1.DFF_0_.D
rlabel metal1 8602 10982 8602 10982 0 mem_bottom_track_1.DFF_0_.Q
rlabel metal1 6118 8466 6118 8466 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal1 4784 9894 4784 9894 0 mem_bottom_track_1.DFF_2_.Q
rlabel metal1 5060 2414 5060 2414 0 mem_bottom_track_1.DFF_3_.Q
rlabel metal1 10488 3638 10488 3638 0 mem_bottom_track_17.DFF_0_.D
rlabel metal1 10258 3162 10258 3162 0 mem_bottom_track_17.DFF_0_.Q
rlabel metal1 12834 5644 12834 5644 0 mem_bottom_track_17.DFF_1_.Q
rlabel metal1 13938 2448 13938 2448 0 mem_bottom_track_17.DFF_2_.Q
rlabel metal1 11040 4590 11040 4590 0 mem_bottom_track_17.DFF_3_.Q
rlabel metal1 5888 17170 5888 17170 0 mem_bottom_track_9.DFF_0_.Q
rlabel metal1 8602 5746 8602 5746 0 mem_bottom_track_9.DFF_1_.Q
rlabel metal1 8510 2414 8510 2414 0 mem_bottom_track_9.DFF_2_.Q
rlabel metal1 13616 4726 13616 4726 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 4738 8398 4738 8398 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 2392 6834 2392 6834 0 mem_left_track_1.DFF_2_.Q
rlabel metal2 3128 13294 3128 13294 0 mem_left_track_1.DFF_3_.Q
rlabel metal1 3864 20910 3864 20910 0 mem_left_track_17.DFF_0_.D
rlabel metal1 5612 20230 5612 20230 0 mem_left_track_17.DFF_0_.Q
rlabel metal2 12742 16864 12742 16864 0 mem_left_track_17.DFF_1_.Q
rlabel metal1 9706 17170 9706 17170 0 mem_left_track_17.DFF_2_.Q
rlabel metal1 6394 19244 6394 19244 0 mem_left_track_9.DFF_0_.Q
rlabel metal1 1702 19788 1702 19788 0 mem_left_track_9.DFF_1_.Q
rlabel metal1 2622 19380 2622 19380 0 mem_left_track_9.DFF_2_.Q
rlabel metal1 6946 11254 6946 11254 0 mem_right_track_0.DFF_0_.D
rlabel metal2 8602 14042 8602 14042 0 mem_right_track_0.DFF_0_.Q
rlabel metal2 12558 14144 12558 14144 0 mem_right_track_0.DFF_1_.Q
rlabel metal1 13110 15878 13110 15878 0 mem_right_track_0.DFF_2_.Q
rlabel metal2 14306 14926 14306 14926 0 mem_right_track_0.DFF_3_.Q
rlabel metal2 4830 17306 4830 17306 0 mem_right_track_16.DFF_0_.D
rlabel metal1 5428 18258 5428 18258 0 mem_right_track_16.DFF_0_.Q
rlabel metal1 7084 14926 7084 14926 0 mem_right_track_16.DFF_1_.Q
rlabel metal1 6762 9520 6762 9520 0 mem_right_track_16.DFF_2_.Q
rlabel metal1 5658 14246 5658 14246 0 mem_right_track_8.DFF_0_.Q
rlabel metal1 1702 13294 1702 13294 0 mem_right_track_8.DFF_1_.Q
rlabel metal1 2438 17238 2438 17238 0 mem_right_track_8.DFF_2_.Q
rlabel metal1 8970 20434 8970 20434 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 10948 12818 10948 12818 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 10350 14382 10350 14382 0 mem_top_track_0.DFF_2_.Q
rlabel metal1 10994 14382 10994 14382 0 mem_top_track_0.DFF_3_.Q
rlabel metal1 12098 7446 12098 7446 0 mem_top_track_16.DFF_0_.D
rlabel metal1 8694 6324 8694 6324 0 mem_top_track_16.DFF_0_.Q
rlabel metal2 1886 9792 1886 9792 0 mem_top_track_16.DFF_1_.Q
rlabel metal1 5796 10642 5796 10642 0 mem_top_track_16.DFF_2_.Q
rlabel metal1 12834 8500 12834 8500 0 mem_top_track_8.DFF_0_.Q
rlabel metal2 9982 10387 9982 10387 0 mem_top_track_8.DFF_1_.Q
rlabel metal2 12742 8160 12742 8160 0 mem_top_track_8.DFF_2_.Q
rlabel metal1 3910 12818 3910 12818 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 6164 13838 6164 13838 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 8280 17102 8280 17102 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 7636 14994 7636 14994 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 7038 2380 7038 2380 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 6348 2414 6348 2414 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 2024 13294 2024 13294 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal1 1932 12954 1932 12954 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 1932 8806 1932 8806 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal1 5198 12104 5198 12104 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7038 12920 7038 12920 0 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 5934 12138 5934 12138 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6118 2550 6118 2550 0 mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2254 10727 2254 10727 0 mux_bottom_track_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 3036 4726 3036 4726 0 mux_bottom_track_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 4922 2550 4922 2550 0 mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3404 3978 3404 3978 0 mux_bottom_track_1.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 5474 3536 5474 3536 0 mux_bottom_track_1.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 9982 18292 9982 18292 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 9982 18122 9982 18122 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 13156 12614 13156 12614 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal2 12558 10727 12558 10727 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 14122 6834 14122 6834 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 11868 14382 11868 14382 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal1 10902 5678 10902 5678 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal1 11960 12614 11960 12614 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal1 11546 18054 11546 18054 0 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14214 11050 14214 11050 0 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 13478 7344 13478 7344 0 mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 12650 5678 12650 5678 0 mux_bottom_track_17.mux_l2_in_2_.TGATE_0_.out
rlabel metal2 12558 6222 12558 6222 0 mux_bottom_track_17.mux_l2_in_3_.TGATE_0_.out
rlabel via1 13386 6222 13386 6222 0 mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 12880 5270 12880 5270 0 mux_bottom_track_17.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 12374 6290 12374 6290 0 mux_bottom_track_17.mux_l4_in_0_.TGATE_0_.out
rlabel metal2 5934 20468 5934 20468 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 5612 20366 5612 20366 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 5474 5066 5474 5066 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 6900 5202 6900 5202 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 6118 5134 6118 5134 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 7176 2414 7176 2414 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal1 8464 6766 8464 6766 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal1 9246 7820 9246 7820 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal1 2415 9894 2415 9894 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 7176 18122 7176 18122 0 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6946 4998 6946 4998 0 mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 7912 5338 7912 5338 0 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8004 2618 8004 2618 0 mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 8464 6086 8464 6086 0 mux_bottom_track_9.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 9936 5814 9936 5814 0 mux_bottom_track_9.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 10074 3978 10074 3978 0 mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 10442 4998 10442 4998 0 mux_bottom_track_9.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 9844 2550 9844 2550 0 mux_bottom_track_9.mux_l4_in_0_.TGATE_0_.out
rlabel metal2 1794 17476 1794 17476 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 5244 8942 5244 8942 0 mux_left_track_1.INVTX1_5_.out
rlabel metal1 5244 8874 5244 8874 0 mux_left_track_1.INVTX1_6_.out
rlabel metal1 6210 7310 6210 7310 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 3174 5202 3174 5202 0 mux_left_track_1.INVTX1_8_.out
rlabel metal2 3726 10030 3726 10030 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 4830 7140 4830 7140 0 mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4278 8602 4278 8602 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5014 6698 5014 6698 0 mux_left_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 4738 7242 4738 7242 0 mux_left_track_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 2392 5542 2392 5542 0 mux_left_track_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 4278 7378 4278 7378 0 mux_left_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 3266 6834 3266 6834 0 mux_left_track_1.mux_l3_in_1_.TGATE_0_.out
rlabel via2 2438 14365 2438 14365 0 mux_left_track_1.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 7222 20910 7222 20910 0 mux_left_track_17.INVTX1_2_.out
rlabel metal2 11914 16405 11914 16405 0 mux_left_track_17.INVTX1_5_.out
rlabel metal1 12466 17034 12466 17034 0 mux_left_track_17.INVTX1_6_.out
rlabel metal1 11638 14994 11638 14994 0 mux_left_track_17.INVTX1_7_.out
rlabel metal2 6210 20740 6210 20740 0 mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 12466 21420 12466 21420 0 mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 12696 13396 12696 13396 0 mux_left_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 12604 17850 12604 17850 0 mux_left_track_17.mux_l2_in_2_.TGATE_0_.out
rlabel metal2 12558 20298 12558 20298 0 mux_left_track_17.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 13662 20978 13662 20978 0 mux_left_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 13202 19754 13202 19754 0 mux_left_track_17.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 14030 19754 14030 19754 0 mux_left_track_17.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 7590 20434 7590 20434 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 6522 15470 6522 15470 0 mux_left_track_9.INVTX1_5_.out
rlabel metal1 2944 16558 2944 16558 0 mux_left_track_9.INVTX1_6_.out
rlabel metal1 2599 18190 2599 18190 0 mux_left_track_9.INVTX1_7_.out
rlabel metal2 2300 17068 2300 17068 0 mux_left_track_9.INVTX1_8_.out
rlabel metal1 9798 18938 9798 18938 0 mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 8694 17850 8694 17850 0 mux_left_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 7820 19414 7820 19414 0 mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6900 16558 6900 16558 0 mux_left_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2438 17952 2438 17952 0 mux_left_track_9.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 2438 18598 2438 18598 0 mux_left_track_9.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 5014 19754 5014 19754 0 mux_left_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3634 19278 3634 19278 0 mux_left_track_9.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 2162 15096 2162 15096 0 mux_left_track_9.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 13340 16558 13340 16558 0 mux_right_track_0.INVTX1_3_.out
rlabel metal2 11638 19176 11638 19176 0 mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 10764 20570 10764 20570 0 mux_right_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 12190 19040 12190 19040 0 mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 12788 17034 12788 17034 0 mux_right_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 12466 15300 12466 15300 0 mux_right_track_0.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 12558 14042 12558 14042 0 mux_right_track_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 13386 17680 13386 17680 0 mux_right_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 12834 15096 12834 15096 0 mux_right_track_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 13892 14518 13892 14518 0 mux_right_track_0.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 6808 18054 6808 18054 0 mux_right_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 7222 15402 7222 15402 0 mux_right_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7084 9078 7084 9078 0 mux_right_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 7728 7854 7728 7854 0 mux_right_track_16.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 8786 8806 8786 8806 0 mux_right_track_16.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 8326 9486 8326 9486 0 mux_right_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 8602 9690 8602 9690 0 mux_right_track_16.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 11776 15606 11776 15606 0 mux_right_track_16.mux_l4_in_0_.TGATE_0_.out
rlabel metal2 7038 14637 7038 14637 0 mux_right_track_8.INVTX1_3_.out
rlabel metal2 4278 13906 4278 13906 0 mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5704 13770 5704 13770 0 mux_right_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4416 14586 4416 14586 0 mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 4094 16558 4094 16558 0 mux_right_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2438 15470 2438 15470 0 mux_right_track_8.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 2484 14790 2484 14790 0 mux_right_track_8.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 4646 16218 4646 16218 0 mux_right_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3496 15606 3496 15606 0 mux_right_track_8.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 12650 15980 12650 15980 0 mux_right_track_8.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 9936 20026 9936 20026 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 9016 17306 9016 17306 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 8234 15674 8234 15674 0 mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9200 16218 9200 16218 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 7038 15776 7038 15776 0 mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 10396 13294 10396 13294 0 mux_top_track_0.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 10764 13838 10764 13838 0 mux_top_track_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 9522 15402 9522 15402 0 mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 11178 14042 11178 14042 0 mux_top_track_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 9706 15606 9706 15606 0 mux_top_track_0.mux_l4_in_0_.TGATE_0_.out
rlabel metal2 6670 6018 6670 6018 0 mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6762 6834 6762 6834 0 mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5750 9486 5750 9486 0 mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2530 11628 2530 11628 0 mux_top_track_16.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 3404 9690 3404 9690 0 mux_top_track_16.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 6992 10234 6992 10234 0 mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 4094 10234 4094 10234 0 mux_top_track_16.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 14352 19346 14352 19346 0 mux_top_track_16.mux_l4_in_0_.TGATE_0_.out
rlabel metal2 13754 12988 13754 12988 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 14076 10778 14076 10778 0 mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13478 8262 13478 8262 0 mux_top_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 13524 9350 13524 9350 0 mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 12834 9724 12834 9724 0 mux_top_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 9936 7718 9936 7718 0 mux_top_track_8.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 10212 9554 10212 9554 0 mux_top_track_8.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 12282 8840 12282 8840 0 mux_top_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 10902 8840 10902 8840 0 mux_top_track_8.mux_l3_in_1_.TGATE_0_.out
rlabel metal3 10695 19380 10695 19380 0 mux_top_track_8.mux_l4_in_0_.TGATE_0_.out
rlabel metal1 7406 3094 7406 3094 0 net1
rlabel metal1 10304 17102 10304 17102 0 net10
rlabel metal1 5515 17578 5515 17578 0 net100
rlabel metal1 4354 17238 4354 17238 0 net101
rlabel via1 10998 3026 10998 3026 0 net102
rlabel metal1 8525 14314 8525 14314 0 net103
rlabel viali 11090 6290 11090 6290 0 net104
rlabel metal1 12542 4522 12542 4522 0 net105
rlabel metal1 11495 12206 11495 12206 0 net106
rlabel metal1 6562 20502 6562 20502 0 net107
rlabel metal1 3588 13498 3588 13498 0 net108
rlabel metal1 8372 5134 8372 5134 0 net109
rlabel metal2 1794 9690 1794 9690 0 net11
rlabel metal1 13482 9962 13482 9962 0 net110
rlabel metal1 7360 9962 7360 9962 0 net111
rlabel metal1 11362 3162 11362 3162 0 net112
rlabel metal1 4058 13974 4058 13974 0 net113
rlabel metal1 8321 11118 8321 11118 0 net114
rlabel via1 9425 3434 9425 3434 0 net115
rlabel via1 2985 17170 2985 17170 0 net116
rlabel via1 13666 15062 13666 15062 0 net117
rlabel metal1 9420 13906 9420 13906 0 net118
rlabel metal1 4328 3094 4328 3094 0 net119
rlabel metal1 1978 9996 1978 9996 0 net12
rlabel metal2 7038 19618 7038 19618 0 net120
rlabel metal2 3082 7378 3082 7378 0 net121
rlabel via1 2893 20434 2893 20434 0 net122
rlabel metal1 8698 3026 8698 3026 0 net123
rlabel metal1 13473 20502 13473 20502 0 net124
rlabel metal1 5566 10778 5566 10778 0 net125
rlabel via1 10354 16082 10354 16082 0 net126
rlabel metal1 10529 7378 10529 7378 0 net127
rlabel metal1 9706 15062 9706 15062 0 net128
rlabel metal1 14030 3706 14030 3706 0 net129
rlabel metal2 10810 6069 10810 6069 0 net13
rlabel metal2 6394 3298 6394 3298 0 net130
rlabel via1 11817 16082 11817 16082 0 net131
rlabel metal1 2576 15674 2576 15674 0 net132
rlabel metal1 2714 7344 2714 7344 0 net133
rlabel metal1 12788 3706 12788 3706 0 net134
rlabel metal2 12466 8296 12466 8296 0 net135
rlabel metal1 11720 20434 11720 20434 0 net136
rlabel metal2 2438 6749 2438 6749 0 net137
rlabel metal2 2530 9282 2530 9282 0 net138
rlabel metal1 8597 13906 8597 13906 0 net139
rlabel metal1 8970 13226 8970 13226 0 net14
rlabel metal1 4692 19414 4692 19414 0 net140
rlabel metal2 6624 14790 6624 14790 0 net141
rlabel metal2 13570 13022 13570 13022 0 net15
rlabel metal1 12719 3638 12719 3638 0 net16
rlabel metal3 2415 19380 2415 19380 0 net17
rlabel metal2 14214 3196 14214 3196 0 net18
rlabel metal1 12834 10166 12834 10166 0 net19
rlabel metal2 2162 3808 2162 3808 0 net2
rlabel metal1 14076 2414 14076 2414 0 net20
rlabel metal1 14444 3502 14444 3502 0 net21
rlabel via2 2070 2533 2070 2533 0 net22
rlabel metal2 1702 2091 1702 2091 0 net23
rlabel metal1 8740 20910 8740 20910 0 net24
rlabel metal2 5750 9112 5750 9112 0 net25
rlabel metal1 3772 17646 3772 17646 0 net26
rlabel metal1 8832 17646 8832 17646 0 net27
rlabel metal2 4830 2244 4830 2244 0 net28
rlabel metal1 2898 2992 2898 2992 0 net29
rlabel metal2 7682 19618 7682 19618 0 net3
rlabel metal1 1840 3638 1840 3638 0 net30
rlabel metal1 3174 12852 3174 12852 0 net31
rlabel metal1 4922 20842 4922 20842 0 net32
rlabel metal3 8004 18904 8004 18904 0 net33
rlabel metal2 1472 20434 1472 20434 0 net34
rlabel metal1 7682 13294 7682 13294 0 net35
rlabel metal1 4922 21590 4922 21590 0 net36
rlabel metal2 9246 20638 9246 20638 0 net37
rlabel metal1 6118 21522 6118 21522 0 net38
rlabel metal1 7130 21590 7130 21590 0 net39
rlabel via2 1702 3043 1702 3043 0 net4
rlabel metal1 1886 12410 1886 12410 0 net40
rlabel metal1 6026 8330 6026 8330 0 net41
rlabel metal1 13340 16762 13340 16762 0 net42
rlabel metal1 13110 16626 13110 16626 0 net43
rlabel via1 10902 17051 10902 17051 0 net44
rlabel metal1 11178 17136 11178 17136 0 net45
rlabel metal1 13662 18734 13662 18734 0 net46
rlabel metal1 2024 14314 2024 14314 0 net47
rlabel metal2 1748 10540 1748 10540 0 net48
rlabel metal2 1748 16932 1748 16932 0 net49
rlabel metal1 13064 12750 13064 12750 0 net5
rlabel via2 1794 17595 1794 17595 0 net50
rlabel metal2 2024 16762 2024 16762 0 net51
rlabel metal1 2070 20502 2070 20502 0 net52
rlabel via3 2139 20740 2139 20740 0 net53
rlabel metal3 1863 20740 1863 20740 0 net54
rlabel metal1 2070 18904 2070 18904 0 net55
rlabel metal2 14306 9622 14306 9622 0 net56
rlabel metal1 14260 9146 14260 9146 0 net57
rlabel metal1 14122 12920 14122 12920 0 net58
rlabel metal2 14122 13158 14122 13158 0 net59
rlabel metal2 15042 9469 15042 9469 0 net6
rlabel metal1 14214 15062 14214 15062 0 net60
rlabel metal2 14214 17340 14214 17340 0 net61
rlabel metal1 14306 17170 14306 17170 0 net62
rlabel metal1 14122 18360 14122 18360 0 net63
rlabel metal2 12558 17238 12558 17238 0 net64
rlabel metal1 8924 2414 8924 2414 0 net65
rlabel metal3 7544 12716 7544 12716 0 net66
rlabel via2 11638 2363 11638 2363 0 net67
rlabel metal3 9867 19380 9867 19380 0 net68
rlabel metal1 12190 2448 12190 2448 0 net69
rlabel metal1 3404 5202 3404 5202 0 net7
rlabel metal2 12742 2159 12742 2159 0 net70
rlabel metal1 12880 2414 12880 2414 0 net71
rlabel metal2 14122 6239 14122 6239 0 net72
rlabel metal1 13248 3094 13248 3094 0 net73
rlabel metal1 7774 21488 7774 21488 0 net74
rlabel metal1 8004 21590 8004 21590 0 net75
rlabel metal2 8510 21318 8510 21318 0 net76
rlabel metal1 9384 21114 9384 21114 0 net77
rlabel metal1 10626 20026 10626 20026 0 net78
rlabel metal1 10120 21590 10120 21590 0 net79
rlabel metal1 13754 12886 13754 12886 0 net8
rlabel metal1 9154 17544 9154 17544 0 net80
rlabel via2 12926 18683 12926 18683 0 net81
rlabel metal2 14214 20026 14214 20026 0 net82
rlabel metal1 10166 12852 10166 12852 0 net83
rlabel metal1 10166 9690 10166 9690 0 net84
rlabel metal2 13386 13600 13386 13600 0 net85
rlabel metal1 2162 14994 2162 14994 0 net86
rlabel metal1 2231 4522 2231 4522 0 net87
rlabel via1 9798 4675 9798 4675 0 net88
rlabel metal1 1656 5746 1656 5746 0 net89
rlabel metal2 15318 16252 15318 16252 0 net9
rlabel metal2 1886 19754 1886 19754 0 net90
rlabel metal1 2530 9044 2530 9044 0 net91
rlabel metal1 8188 8466 8188 8466 0 net92
rlabel metal1 11776 4522 11776 4522 0 net93
rlabel metal1 11914 20910 11914 20910 0 net94
rlabel metal1 10176 11118 10176 11118 0 net95
rlabel via1 7677 13226 7677 13226 0 net96
rlabel metal1 6036 6290 6036 6290 0 net97
rlabel via1 4733 3434 4733 3434 0 net98
rlabel metal1 4595 20502 4595 20502 0 net99
rlabel via2 4094 13413 4094 13413 0 prog_clk
rlabel metal2 13570 18241 13570 18241 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 12098 20468 12098 20468 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 14214 22695 14214 22695 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 15003 23324 15003 23324 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
<< properties >>
string FIXED_BBOX 0 0 16000 24000
<< end >>
