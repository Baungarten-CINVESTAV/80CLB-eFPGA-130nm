magic
tech sky130A
magscale 1 2
timestamp 1708041177
<< viali >>
rect 1685 15657 1719 15691
rect 16221 15657 16255 15691
rect 1961 15453 1995 15487
rect 2789 15453 2823 15487
rect 3249 15453 3283 15487
rect 4353 15453 4387 15487
rect 5917 15453 5951 15487
rect 7481 15453 7515 15487
rect 9045 15453 9079 15487
rect 10793 15453 10827 15487
rect 12357 15453 12391 15487
rect 13921 15453 13955 15487
rect 14933 15453 14967 15487
rect 15209 15453 15243 15487
rect 2513 15385 2547 15419
rect 15669 15385 15703 15419
rect 15945 15385 15979 15419
rect 2237 15317 2271 15351
rect 2973 15317 3007 15351
rect 3065 15317 3099 15351
rect 4537 15317 4571 15351
rect 6101 15317 6135 15351
rect 7665 15317 7699 15351
rect 9229 15317 9263 15351
rect 10609 15317 10643 15351
rect 12173 15317 12207 15351
rect 13737 15317 13771 15351
rect 14749 15317 14783 15351
rect 15025 15317 15059 15351
rect 15577 15317 15611 15351
rect 1501 15113 1535 15147
rect 4997 15113 5031 15147
rect 11621 15113 11655 15147
rect 15761 15113 15795 15147
rect 16405 15113 16439 15147
rect 1777 14977 1811 15011
rect 2237 14977 2271 15011
rect 2329 14977 2363 15011
rect 2605 14977 2639 15011
rect 5181 14977 5215 15011
rect 7481 14977 7515 15011
rect 9965 14977 9999 15011
rect 11805 14977 11839 15011
rect 14381 14977 14415 15011
rect 14841 14977 14875 15011
rect 15301 14977 15335 15011
rect 15577 14977 15611 15011
rect 15669 14977 15703 15011
rect 16129 14977 16163 15011
rect 14473 14909 14507 14943
rect 10057 14841 10091 14875
rect 2513 14773 2547 14807
rect 7573 14773 7607 14807
rect 14933 14773 14967 14807
rect 15485 14773 15519 14807
rect 8769 14365 8803 14399
rect 9321 14365 9355 14399
rect 10333 14365 10367 14399
rect 10609 14365 10643 14399
rect 11989 14365 12023 14399
rect 13369 14365 13403 14399
rect 14841 14365 14875 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 16129 14365 16163 14399
rect 1409 14297 1443 14331
rect 1777 14297 1811 14331
rect 13277 14297 13311 14331
rect 16497 14297 16531 14331
rect 8585 14229 8619 14263
rect 9413 14229 9447 14263
rect 10517 14229 10551 14263
rect 10793 14229 10827 14263
rect 12081 14229 12115 14263
rect 14749 14229 14783 14263
rect 15209 14229 15243 14263
rect 15577 14229 15611 14263
rect 15761 14229 15795 14263
rect 10241 14025 10275 14059
rect 13553 14025 13587 14059
rect 13829 14025 13863 14059
rect 16129 13957 16163 13991
rect 1777 13889 1811 13923
rect 9045 13889 9079 13923
rect 9505 13889 9539 13923
rect 10057 13889 10091 13923
rect 10333 13889 10367 13923
rect 11069 13889 11103 13923
rect 12449 13889 12483 13923
rect 12541 13889 12575 13923
rect 13001 13889 13035 13923
rect 13369 13889 13403 13923
rect 13645 13889 13679 13923
rect 14473 13889 14507 13923
rect 14657 13889 14691 13923
rect 14749 13889 14783 13923
rect 14841 13889 14875 13923
rect 15393 13889 15427 13923
rect 16497 13889 16531 13923
rect 1501 13821 1535 13855
rect 8953 13821 8987 13855
rect 9321 13821 9355 13855
rect 11253 13821 11287 13855
rect 11529 13821 11563 13855
rect 13093 13821 13127 13855
rect 15117 13821 15151 13855
rect 15761 13821 15795 13855
rect 9229 13753 9263 13787
rect 9689 13685 9723 13719
rect 10425 13685 10459 13719
rect 10701 13685 10735 13719
rect 12173 13685 12207 13719
rect 12265 13685 12299 13719
rect 12633 13685 12667 13719
rect 12817 13685 12851 13719
rect 14289 13685 14323 13719
rect 8769 13481 8803 13515
rect 10701 13481 10735 13515
rect 13461 13481 13495 13515
rect 15117 13481 15151 13515
rect 15669 13481 15703 13515
rect 11529 13413 11563 13447
rect 12357 13413 12391 13447
rect 10333 13345 10367 13379
rect 11805 13345 11839 13379
rect 12725 13345 12759 13379
rect 12909 13345 12943 13379
rect 15209 13345 15243 13379
rect 15393 13345 15427 13379
rect 8585 13277 8619 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 10149 13277 10183 13311
rect 13645 13277 13679 13311
rect 13737 13277 13771 13311
rect 14197 13277 14231 13311
rect 14473 13277 14507 13311
rect 14657 13277 14691 13311
rect 16037 13277 16071 13311
rect 16405 13277 16439 13311
rect 10977 13209 11011 13243
rect 11069 13209 11103 13243
rect 11897 13209 11931 13243
rect 9229 13141 9263 13175
rect 10057 13141 10091 13175
rect 13369 13141 13403 13175
rect 13829 13141 13863 13175
rect 14381 13141 14415 13175
rect 2053 12937 2087 12971
rect 9505 12937 9539 12971
rect 11161 12937 11195 12971
rect 15301 12937 15335 12971
rect 4629 12869 4663 12903
rect 11796 12869 11830 12903
rect 15761 12869 15795 12903
rect 1777 12801 1811 12835
rect 2145 12801 2179 12835
rect 4537 12801 4571 12835
rect 5457 12801 5491 12835
rect 9045 12801 9079 12835
rect 9597 12801 9631 12835
rect 9864 12801 9898 12835
rect 11069 12801 11103 12835
rect 11529 12801 11563 12835
rect 13737 12801 13771 12835
rect 13921 12801 13955 12835
rect 15485 12801 15519 12835
rect 8861 12733 8895 12767
rect 13553 12733 13587 12767
rect 15025 12733 15059 12767
rect 15669 12733 15703 12767
rect 15945 12733 15979 12767
rect 5273 12665 5307 12699
rect 10977 12665 11011 12699
rect 14289 12665 14323 12699
rect 1501 12597 1535 12631
rect 12909 12597 12943 12631
rect 13001 12597 13035 12631
rect 14473 12597 14507 12631
rect 8953 12393 8987 12427
rect 12449 12393 12483 12427
rect 13921 12393 13955 12427
rect 7665 12257 7699 12291
rect 10333 12257 10367 12291
rect 12541 12257 12575 12291
rect 2145 12189 2179 12223
rect 7849 12189 7883 12223
rect 10609 12189 10643 12223
rect 11161 12189 11195 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 15485 12189 15519 12223
rect 16129 12189 16163 12223
rect 16497 12189 16531 12223
rect 1409 12121 1443 12155
rect 1777 12121 1811 12155
rect 10088 12121 10122 12155
rect 12808 12121 12842 12155
rect 15240 12121 15274 12155
rect 15577 12121 15611 12155
rect 1961 12053 1995 12087
rect 8309 12053 8343 12087
rect 10517 12053 10551 12087
rect 11345 12053 11379 12087
rect 14105 12053 14139 12087
rect 16313 12053 16347 12087
rect 6929 11849 6963 11883
rect 7021 11849 7055 11883
rect 8677 11849 8711 11883
rect 10333 11849 10367 11883
rect 12633 11849 12667 11883
rect 15393 11849 15427 11883
rect 8953 11781 8987 11815
rect 9045 11781 9079 11815
rect 14280 11781 14314 11815
rect 5733 11713 5767 11747
rect 6745 11713 6779 11747
rect 7205 11713 7239 11747
rect 7564 11713 7598 11747
rect 9781 11713 9815 11747
rect 10609 11713 10643 11747
rect 10885 11713 10919 11747
rect 12725 11713 12759 11747
rect 14013 11713 14047 11747
rect 16221 11713 16255 11747
rect 7297 11645 7331 11679
rect 9597 11645 9631 11679
rect 10701 11645 10735 11679
rect 11529 11645 11563 11679
rect 11713 11645 11747 11679
rect 13737 11645 13771 11679
rect 5641 11509 5675 11543
rect 10425 11509 10459 11543
rect 11345 11509 11379 11543
rect 11897 11509 11931 11543
rect 15669 11509 15703 11543
rect 7481 11305 7515 11339
rect 7573 11305 7607 11339
rect 9045 11305 9079 11339
rect 16221 11305 16255 11339
rect 2237 11237 2271 11271
rect 5641 11169 5675 11203
rect 6101 11169 6135 11203
rect 6285 11169 6319 11203
rect 7021 11169 7055 11203
rect 8585 11169 8619 11203
rect 11989 11169 12023 11203
rect 12633 11169 12667 11203
rect 13553 11169 13587 11203
rect 16037 11169 16071 11203
rect 1777 11101 1811 11135
rect 2421 11101 2455 11135
rect 2973 11101 3007 11135
rect 5457 11101 5491 11135
rect 6837 11101 6871 11135
rect 8217 11101 8251 11135
rect 8677 11101 8711 11135
rect 9137 11101 9171 11135
rect 9597 11101 9631 11135
rect 11161 11101 11195 11135
rect 12909 11101 12943 11135
rect 16129 11101 16163 11135
rect 1409 11033 1443 11067
rect 3065 11033 3099 11067
rect 6745 11033 6779 11067
rect 9505 11033 9539 11067
rect 9965 11033 9999 11067
rect 10057 11033 10091 11067
rect 10609 11033 10643 11067
rect 12081 11033 12115 11067
rect 13737 11033 13771 11067
rect 13829 11033 13863 11067
rect 14197 11033 14231 11067
rect 14565 11033 14599 11067
rect 15770 11033 15804 11067
rect 4997 10965 5031 10999
rect 9781 10965 9815 10999
rect 11345 10965 11379 10999
rect 13093 10965 13127 10999
rect 14657 10965 14691 10999
rect 4721 10761 4755 10795
rect 4813 10761 4847 10795
rect 7205 10761 7239 10795
rect 7481 10761 7515 10795
rect 12081 10761 12115 10795
rect 12541 10761 12575 10795
rect 12817 10761 12851 10795
rect 7021 10693 7055 10727
rect 15761 10693 15795 10727
rect 15853 10693 15887 10727
rect 1777 10625 1811 10659
rect 4261 10625 4295 10659
rect 4537 10625 4571 10659
rect 5273 10625 5307 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 6009 10625 6043 10659
rect 7297 10625 7331 10659
rect 8605 10625 8639 10659
rect 9045 10625 9079 10659
rect 9321 10625 9355 10659
rect 10333 10625 10367 10659
rect 10517 10625 10551 10659
rect 12173 10625 12207 10659
rect 12357 10625 12391 10659
rect 12633 10625 12667 10659
rect 12909 10625 12943 10659
rect 13277 10625 13311 10659
rect 13461 10625 13495 10659
rect 14749 10625 14783 10659
rect 5457 10557 5491 10591
rect 6377 10557 6411 10591
rect 6561 10557 6595 10591
rect 8861 10557 8895 10591
rect 10057 10557 10091 10591
rect 10241 10557 10275 10591
rect 14841 10557 14875 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 4445 10489 4479 10523
rect 6193 10489 6227 10523
rect 9137 10489 9171 10523
rect 13093 10489 13127 10523
rect 14105 10489 14139 10523
rect 1501 10421 1535 10455
rect 9505 10421 9539 10455
rect 9873 10421 9907 10455
rect 10701 10421 10735 10455
rect 13921 10421 13955 10455
rect 15209 10421 15243 10455
rect 6561 10217 6595 10251
rect 8953 10217 8987 10251
rect 9965 10217 9999 10251
rect 13829 10217 13863 10251
rect 6469 10149 6503 10183
rect 11713 10149 11747 10183
rect 4905 10081 4939 10115
rect 8033 10081 8067 10115
rect 13645 10081 13679 10115
rect 14105 10081 14139 10115
rect 14841 10081 14875 10115
rect 16313 10081 16347 10115
rect 3801 10013 3835 10047
rect 5089 10013 5123 10047
rect 5825 10015 5859 10049
rect 6101 10013 6135 10047
rect 6285 10013 6319 10047
rect 6737 10009 6771 10043
rect 6837 10013 6871 10047
rect 8217 10013 8251 10047
rect 8309 10013 8343 10047
rect 8769 10013 8803 10047
rect 9505 10013 9539 10047
rect 9689 10013 9723 10047
rect 10149 10013 10183 10047
rect 13389 10013 13423 10047
rect 13737 10013 13771 10047
rect 14657 10013 14691 10047
rect 15025 10013 15059 10047
rect 7481 9945 7515 9979
rect 10425 9945 10459 9979
rect 15669 9945 15703 9979
rect 16221 9945 16255 9979
rect 4445 9877 4479 9911
rect 5549 9877 5583 9911
rect 5733 9877 5767 9911
rect 5917 9877 5951 9911
rect 7573 9877 7607 9911
rect 8585 9877 8619 9911
rect 9873 9877 9907 9911
rect 12265 9877 12299 9911
rect 15485 9877 15519 9911
rect 14473 9673 14507 9707
rect 4160 9605 4194 9639
rect 5549 9605 5583 9639
rect 6101 9605 6135 9639
rect 10210 9605 10244 9639
rect 13216 9605 13250 9639
rect 16405 9605 16439 9639
rect 3545 9537 3579 9571
rect 6377 9537 6411 9571
rect 6644 9537 6678 9571
rect 7849 9537 7883 9571
rect 9137 9537 9171 9571
rect 9965 9537 9999 9571
rect 11621 9537 11655 9571
rect 11713 9537 11747 9571
rect 14381 9537 14415 9571
rect 14924 9537 14958 9571
rect 16313 9537 16347 9571
rect 3801 9469 3835 9503
rect 3893 9469 3927 9503
rect 5457 9469 5491 9503
rect 8125 9469 8159 9503
rect 8309 9469 8343 9503
rect 9229 9469 9263 9503
rect 9413 9469 9447 9503
rect 13461 9469 13495 9503
rect 14105 9469 14139 9503
rect 14657 9469 14691 9503
rect 2421 9401 2455 9435
rect 8033 9401 8067 9435
rect 9045 9401 9079 9435
rect 11345 9401 11379 9435
rect 5273 9333 5307 9367
rect 7757 9333 7791 9367
rect 8493 9333 8527 9367
rect 9873 9333 9907 9367
rect 12081 9333 12115 9367
rect 13553 9333 13587 9367
rect 16037 9333 16071 9367
rect 4721 9129 4755 9163
rect 6377 9129 6411 9163
rect 7205 9129 7239 9163
rect 7941 9129 7975 9163
rect 10609 9129 10643 9163
rect 16405 9129 16439 9163
rect 5917 9061 5951 9095
rect 11713 9061 11747 9095
rect 12081 9061 12115 9095
rect 13921 9061 13955 9095
rect 15301 9061 15335 9095
rect 7021 8993 7055 9027
rect 15853 8993 15887 9027
rect 1777 8925 1811 8959
rect 4629 8925 4663 8959
rect 6009 8925 6043 8959
rect 6285 8925 6319 8959
rect 7757 8925 7791 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 11529 8925 11563 8959
rect 12265 8925 12299 8959
rect 12449 8925 12483 8959
rect 12541 8925 12575 8959
rect 12808 8925 12842 8959
rect 14657 8925 14691 8959
rect 14933 8925 14967 8959
rect 1409 8857 1443 8891
rect 4905 8857 4939 8891
rect 5457 8857 5491 8891
rect 5549 8857 5583 8891
rect 6193 8857 6227 8891
rect 15761 8857 15795 8891
rect 16129 8857 16163 8891
rect 4169 8789 4203 8823
rect 9045 8789 9079 8823
rect 14105 8789 14139 8823
rect 15117 8789 15151 8823
rect 1777 8585 1811 8619
rect 5917 8585 5951 8619
rect 6193 8585 6227 8619
rect 8493 8585 8527 8619
rect 8677 8585 8711 8619
rect 9781 8585 9815 8619
rect 10517 8585 10551 8619
rect 12173 8585 12207 8619
rect 12817 8585 12851 8619
rect 14473 8585 14507 8619
rect 15209 8585 15243 8619
rect 15945 8585 15979 8619
rect 16221 8585 16255 8619
rect 16405 8585 16439 8619
rect 13093 8517 13127 8551
rect 13185 8517 13219 8551
rect 13737 8517 13771 8551
rect 1869 8449 1903 8483
rect 3709 8449 3743 8483
rect 3801 8449 3835 8483
rect 4077 8449 4111 8483
rect 5733 8449 5767 8483
rect 6009 8449 6043 8483
rect 6377 8449 6411 8483
rect 7297 8449 7331 8483
rect 8033 8449 8067 8483
rect 8769 8449 8803 8483
rect 9045 8449 9079 8483
rect 9321 8449 9355 8483
rect 9597 8449 9631 8483
rect 10057 8449 10091 8483
rect 10609 8449 10643 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12357 8449 12391 8483
rect 12633 8449 12667 8483
rect 12909 8449 12943 8483
rect 14013 8449 14047 8483
rect 14657 8449 14691 8483
rect 16037 8449 16071 8483
rect 16313 8449 16347 8483
rect 4261 8381 4295 8415
rect 4813 8381 4847 8415
rect 4997 8381 5031 8415
rect 6561 8381 6595 8415
rect 7113 8381 7147 8415
rect 7849 8381 7883 8415
rect 9873 8381 9907 8415
rect 10793 8381 10827 8415
rect 11621 8381 11655 8415
rect 13829 8381 13863 8415
rect 15301 8381 15335 8415
rect 15485 8381 15519 8415
rect 3985 8313 4019 8347
rect 4721 8313 4755 8347
rect 5181 8313 5215 8347
rect 7021 8313 7055 8347
rect 8861 8313 8895 8347
rect 9505 8313 9539 8347
rect 3525 8245 3559 8279
rect 7665 8245 7699 8279
rect 11161 8245 11195 8279
rect 11897 8245 11931 8279
rect 12449 8245 12483 8279
rect 3617 8041 3651 8075
rect 5181 8041 5215 8075
rect 5733 8041 5767 8075
rect 7113 8041 7147 8075
rect 7665 8041 7699 8075
rect 14473 8041 14507 8075
rect 4077 7973 4111 8007
rect 9045 7973 9079 8007
rect 13829 7973 13863 8007
rect 7941 7905 7975 7939
rect 8309 7905 8343 7939
rect 10425 7905 10459 7939
rect 12817 7905 12851 7939
rect 14841 7905 14875 7939
rect 2145 7837 2179 7871
rect 3157 7837 3191 7871
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 7297 7837 7331 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 8677 7837 8711 7871
rect 12909 7837 12943 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 15108 7837 15142 7871
rect 1409 7769 1443 7803
rect 1777 7769 1811 7803
rect 7021 7769 7055 7803
rect 10180 7769 10214 7803
rect 10517 7769 10551 7803
rect 11069 7769 11103 7803
rect 11161 7769 11195 7803
rect 12572 7769 12606 7803
rect 13277 7769 13311 7803
rect 13369 7769 13403 7803
rect 1961 7701 1995 7735
rect 3341 7701 3375 7735
rect 4445 7701 4479 7735
rect 8585 7701 8619 7735
rect 11437 7701 11471 7735
rect 13093 7701 13127 7735
rect 16221 7701 16255 7735
rect 3065 7497 3099 7531
rect 3801 7497 3835 7531
rect 3893 7497 3927 7531
rect 5549 7497 5583 7531
rect 5917 7497 5951 7531
rect 7757 7497 7791 7531
rect 7849 7497 7883 7531
rect 11529 7497 11563 7531
rect 13001 7497 13035 7531
rect 14197 7497 14231 7531
rect 9312 7429 9346 7463
rect 10517 7429 10551 7463
rect 11069 7429 11103 7463
rect 12909 7429 12943 7463
rect 14657 7429 14691 7463
rect 15393 7429 15427 7463
rect 1777 7361 1811 7395
rect 2881 7361 2915 7395
rect 3341 7361 3375 7395
rect 4353 7361 4387 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 5733 7361 5767 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6644 7361 6678 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 12449 7361 12483 7395
rect 13461 7361 13495 7395
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 14289 7361 14323 7395
rect 16313 7361 16347 7395
rect 3157 7293 3191 7327
rect 4537 7293 4571 7327
rect 8309 7293 8343 7327
rect 8493 7293 8527 7327
rect 11161 7293 11195 7327
rect 12081 7293 12115 7327
rect 12265 7293 12299 7327
rect 13645 7293 13679 7327
rect 15117 7293 15151 7327
rect 15301 7293 15335 7327
rect 15853 7293 15887 7327
rect 16037 7293 16071 7327
rect 14473 7225 14507 7259
rect 1501 7157 1535 7191
rect 5273 7157 5307 7191
rect 6193 7157 6227 7191
rect 8585 7157 8619 7191
rect 10425 7157 10459 7191
rect 13829 7157 13863 7191
rect 16129 7157 16163 7191
rect 6469 6953 6503 6987
rect 7573 6953 7607 6987
rect 10333 6953 10367 6987
rect 11069 6953 11103 6987
rect 13093 6953 13127 6987
rect 2973 6817 3007 6851
rect 4997 6817 5031 6851
rect 5641 6817 5675 6851
rect 9505 6817 9539 6851
rect 10885 6817 10919 6851
rect 13277 6817 13311 6851
rect 13829 6817 13863 6851
rect 14105 6817 14139 6851
rect 14841 6817 14875 6851
rect 15761 6817 15795 6851
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 4721 6749 4755 6783
rect 5457 6749 5491 6783
rect 6377 6749 6411 6783
rect 7113 6749 7147 6783
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 9413 6749 9447 6783
rect 11253 6749 11287 6783
rect 11621 6749 11655 6783
rect 11897 6749 11931 6783
rect 12265 6749 12299 6783
rect 12541 6749 12575 6783
rect 13461 6749 13495 6783
rect 13921 6749 13955 6783
rect 14565 6749 14599 6783
rect 15945 6749 15979 6783
rect 3065 6681 3099 6715
rect 3617 6681 3651 6715
rect 8677 6681 8711 6715
rect 11989 6681 12023 6715
rect 15393 6681 15427 6715
rect 15485 6681 15519 6715
rect 4353 6613 4387 6647
rect 4629 6613 4663 6647
rect 4905 6613 4939 6647
rect 5733 6613 5767 6647
rect 11345 6613 11379 6647
rect 11805 6613 11839 6647
rect 12449 6613 12483 6647
rect 12725 6613 12759 6647
rect 14381 6613 14415 6647
rect 16405 6613 16439 6647
rect 3249 6409 3283 6443
rect 4721 6409 4755 6443
rect 7021 6409 7055 6443
rect 7481 6409 7515 6443
rect 7849 6409 7883 6443
rect 10609 6409 10643 6443
rect 15393 6409 15427 6443
rect 15669 6409 15703 6443
rect 1777 6341 1811 6375
rect 12449 6341 12483 6375
rect 13001 6341 13035 6375
rect 14381 6341 14415 6375
rect 14933 6341 14967 6375
rect 3341 6273 3375 6307
rect 5926 6273 5960 6307
rect 6193 6273 6227 6307
rect 6561 6273 6595 6307
rect 7297 6273 7331 6307
rect 7573 6273 7607 6307
rect 8309 6273 8343 6307
rect 8493 6273 8527 6307
rect 8769 6273 8803 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9404 6273 9438 6307
rect 11253 6273 11287 6307
rect 13277 6273 13311 6307
rect 14105 6273 14139 6307
rect 15209 6273 15243 6307
rect 15509 6277 15543 6311
rect 15945 6273 15979 6307
rect 16313 6273 16347 6307
rect 4077 6205 4111 6239
rect 4261 6205 4295 6239
rect 6377 6205 6411 6239
rect 11069 6205 11103 6239
rect 11989 6205 12023 6239
rect 12173 6205 12207 6239
rect 13093 6205 13127 6239
rect 15025 6205 15059 6239
rect 7757 6137 7791 6171
rect 11529 6137 11563 6171
rect 13461 6137 13495 6171
rect 15761 6137 15795 6171
rect 1501 6069 1535 6103
rect 4813 6069 4847 6103
rect 8585 6069 8619 6103
rect 8861 6069 8895 6103
rect 10517 6069 10551 6103
rect 13553 6069 13587 6103
rect 16129 6069 16163 6103
rect 5181 5865 5215 5899
rect 7205 5865 7239 5899
rect 11897 5865 11931 5899
rect 12265 5865 12299 5899
rect 12725 5865 12759 5899
rect 13461 5865 13495 5899
rect 14749 5865 14783 5899
rect 15301 5865 15335 5899
rect 7481 5797 7515 5831
rect 8953 5797 8987 5831
rect 9413 5797 9447 5831
rect 8309 5729 8343 5763
rect 13093 5729 13127 5763
rect 14289 5729 14323 5763
rect 15025 5729 15059 5763
rect 2145 5661 2179 5695
rect 3801 5661 3835 5695
rect 7021 5661 7055 5695
rect 7113 5661 7147 5695
rect 7665 5661 7699 5695
rect 8493 5661 8527 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 10149 5661 10183 5695
rect 10425 5661 10459 5695
rect 12449 5657 12483 5691
rect 12541 5661 12575 5695
rect 13001 5661 13035 5695
rect 13277 5661 13311 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 14841 5661 14875 5695
rect 15577 5661 15611 5695
rect 16037 5661 16071 5695
rect 16221 5661 16255 5695
rect 16497 5661 16531 5695
rect 1777 5593 1811 5627
rect 2053 5593 2087 5627
rect 4068 5593 4102 5627
rect 9505 5593 9539 5627
rect 1501 5525 1535 5559
rect 5733 5525 5767 5559
rect 7757 5525 7791 5559
rect 8677 5525 8711 5559
rect 13921 5525 13955 5559
rect 16313 5525 16347 5559
rect 4261 5321 4295 5355
rect 8309 5321 8343 5355
rect 9873 5321 9907 5355
rect 10701 5321 10735 5355
rect 12357 5321 12391 5355
rect 15853 5321 15887 5355
rect 16405 5321 16439 5355
rect 5457 5253 5491 5287
rect 8953 5253 8987 5287
rect 3913 5185 3947 5219
rect 4169 5185 4203 5219
rect 4997 5185 5031 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 7573 5185 7607 5219
rect 7941 5185 7975 5219
rect 8033 5185 8067 5219
rect 8125 5185 8159 5219
rect 8861 5185 8895 5219
rect 9597 5185 9631 5219
rect 11161 5185 11195 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 13481 5185 13515 5219
rect 13737 5185 13771 5219
rect 14381 5185 14415 5219
rect 15669 5185 15703 5219
rect 15945 5185 15979 5219
rect 16221 5185 16255 5219
rect 16313 5185 16347 5219
rect 4813 5117 4847 5151
rect 5365 5117 5399 5151
rect 6837 5117 6871 5151
rect 7757 5117 7791 5151
rect 8585 5117 8619 5151
rect 9413 5117 9447 5151
rect 10425 5117 10459 5151
rect 11345 5117 11379 5151
rect 13829 5117 13863 5151
rect 15209 5117 15243 5151
rect 15393 5117 15427 5151
rect 5917 5049 5951 5083
rect 11805 5049 11839 5083
rect 2789 4981 2823 5015
rect 5181 4981 5215 5015
rect 6377 4981 6411 5015
rect 8769 4981 8803 5015
rect 11529 4981 11563 5015
rect 14749 4981 14783 5015
rect 15485 4981 15519 5015
rect 16129 4981 16163 5015
rect 4445 4777 4479 4811
rect 8677 4777 8711 4811
rect 10333 4777 10367 4811
rect 13369 4777 13403 4811
rect 14657 4777 14691 4811
rect 6009 4709 6043 4743
rect 15117 4709 15151 4743
rect 15853 4709 15887 4743
rect 4261 4641 4295 4675
rect 4629 4641 4663 4675
rect 5273 4641 5307 4675
rect 5457 4641 5491 4675
rect 8953 4641 8987 4675
rect 15485 4641 15519 4675
rect 16221 4641 16255 4675
rect 3801 4573 3835 4607
rect 4537 4573 4571 4607
rect 4813 4573 4847 4607
rect 6377 4573 6411 4607
rect 7021 4573 7055 4607
rect 8585 4573 8619 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 13461 4573 13495 4607
rect 13737 4573 13771 4607
rect 14197 4573 14231 4607
rect 14473 4573 14507 4607
rect 14749 4573 14783 4607
rect 14933 4573 14967 4607
rect 15669 4573 15703 4607
rect 1409 4505 1443 4539
rect 1777 4505 1811 4539
rect 5549 4505 5583 4539
rect 6929 4505 6963 4539
rect 7266 4505 7300 4539
rect 9220 4505 9254 4539
rect 11652 4505 11686 4539
rect 12234 4505 12268 4539
rect 3985 4437 4019 4471
rect 8401 4437 8435 4471
rect 10517 4437 10551 4471
rect 13553 4437 13587 4471
rect 13921 4437 13955 4471
rect 14381 4437 14415 4471
rect 4537 4233 4571 4267
rect 5273 4233 5307 4267
rect 6377 4233 6411 4267
rect 12081 4233 12115 4267
rect 14381 4233 14415 4267
rect 1777 4165 1811 4199
rect 8401 4165 8435 4199
rect 9229 4165 9263 4199
rect 15209 4165 15243 4199
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 4997 4097 5031 4131
rect 5457 4097 5491 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 7490 4097 7524 4131
rect 7941 4097 7975 4131
rect 9873 4097 9907 4131
rect 10241 4097 10275 4131
rect 10977 4097 11011 4131
rect 11805 4097 11839 4131
rect 12725 4097 12759 4131
rect 13277 4097 13311 4131
rect 13461 4097 13495 4131
rect 14013 4097 14047 4131
rect 14197 4097 14231 4131
rect 14289 4097 14323 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 16405 4097 16439 4131
rect 5089 4029 5123 4063
rect 7757 4029 7791 4063
rect 8309 4029 8343 4063
rect 9137 4029 9171 4063
rect 9781 4029 9815 4063
rect 11161 4029 11195 4063
rect 14565 4029 14599 4063
rect 14749 4029 14783 4063
rect 15761 4029 15795 4063
rect 15945 4029 15979 4063
rect 4721 3961 4755 3995
rect 8125 3961 8159 3995
rect 8861 3961 8895 3995
rect 10057 3961 10091 3995
rect 11989 3961 12023 3995
rect 1501 3893 1535 3927
rect 10333 3893 10367 3927
rect 10701 3893 10735 3927
rect 13093 3893 13127 3927
rect 13553 3893 13587 3927
rect 3801 3689 3835 3723
rect 9597 3689 9631 3723
rect 10701 3689 10735 3723
rect 14565 3689 14599 3723
rect 15117 3689 15151 3723
rect 15669 3689 15703 3723
rect 16129 3689 16163 3723
rect 16313 3689 16347 3723
rect 8033 3621 8067 3655
rect 8493 3621 8527 3655
rect 14289 3621 14323 3655
rect 7205 3553 7239 3587
rect 7573 3553 7607 3587
rect 10241 3553 10275 3587
rect 10425 3553 10459 3587
rect 11253 3553 11287 3587
rect 13277 3553 13311 3587
rect 15393 3553 15427 3587
rect 3985 3485 4019 3519
rect 6837 3485 6871 3519
rect 7113 3485 7147 3519
rect 7389 3485 7423 3519
rect 8125 3485 8159 3519
rect 8309 3485 8343 3519
rect 8953 3485 8987 3519
rect 11437 3485 11471 3519
rect 12081 3485 12115 3519
rect 12173 3485 12207 3519
rect 13093 3485 13127 3519
rect 13553 3485 13587 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 14381 3501 14415 3535
rect 14657 3485 14691 3519
rect 15025 3485 15059 3519
rect 15301 3485 15335 3519
rect 15577 3485 15611 3519
rect 16037 3485 16071 3519
rect 16497 3485 16531 3519
rect 7021 3349 7055 3383
rect 11897 3349 11931 3383
rect 12265 3349 12299 3383
rect 12633 3349 12667 3383
rect 13369 3349 13403 3383
rect 13921 3349 13955 3383
rect 14841 3349 14875 3383
rect 1961 3145 1995 3179
rect 2973 3145 3007 3179
rect 6929 3145 6963 3179
rect 7481 3145 7515 3179
rect 7665 3145 7699 3179
rect 8309 3145 8343 3179
rect 10977 3145 11011 3179
rect 11621 3145 11655 3179
rect 13001 3145 13035 3179
rect 13185 3145 13219 3179
rect 13461 3145 13495 3179
rect 13921 3145 13955 3179
rect 15669 3145 15703 3179
rect 15945 3145 15979 3179
rect 16313 3145 16347 3179
rect 1777 3077 1811 3111
rect 8033 3077 8067 3111
rect 2145 3009 2179 3043
rect 2881 3009 2915 3043
rect 6837 3009 6871 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 11069 3009 11103 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 13277 3009 13311 3043
rect 13369 3009 13403 3043
rect 14013 3009 14047 3043
rect 14289 3009 14323 3043
rect 14381 3009 14415 3043
rect 14657 3009 14691 3043
rect 16037 3009 16071 3043
rect 16497 3009 16531 3043
rect 12081 2941 12115 2975
rect 12357 2941 12391 2975
rect 12541 2941 12575 2975
rect 14473 2941 14507 2975
rect 15025 2941 15059 2975
rect 15209 2941 15243 2975
rect 14105 2873 14139 2907
rect 14841 2873 14875 2907
rect 1501 2805 1535 2839
rect 11345 2805 11379 2839
rect 2145 2601 2179 2635
rect 4077 2601 4111 2635
rect 5549 2601 5583 2635
rect 7021 2601 7055 2635
rect 8493 2601 8527 2635
rect 9781 2601 9815 2635
rect 11805 2601 11839 2635
rect 12449 2601 12483 2635
rect 13185 2601 13219 2635
rect 14197 2601 14231 2635
rect 14657 2601 14691 2635
rect 16037 2601 16071 2635
rect 2605 2533 2639 2567
rect 11069 2533 11103 2567
rect 12173 2533 12207 2567
rect 13645 2533 13679 2567
rect 14841 2533 14875 2567
rect 15117 2533 15151 2567
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 3893 2397 3927 2431
rect 5365 2397 5399 2431
rect 6837 2397 6871 2431
rect 8309 2397 8343 2431
rect 9965 2397 9999 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 10885 2397 10919 2431
rect 11345 2397 11379 2431
rect 11621 2397 11655 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13001 2397 13035 2431
rect 13461 2397 13495 2431
rect 13921 2397 13955 2431
rect 14381 2397 14415 2431
rect 14749 2397 14783 2431
rect 15025 2397 15059 2431
rect 15301 2397 15335 2431
rect 15669 2397 15703 2431
rect 15853 2397 15887 2431
rect 16129 2397 16163 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 10517 2261 10551 2295
rect 10793 2261 10827 2295
rect 11253 2261 11287 2295
rect 11897 2261 11931 2295
rect 12817 2261 12851 2295
rect 13737 2261 13771 2295
rect 15485 2261 15519 2295
rect 16221 2261 16255 2295
<< metal1 >>
rect 1104 15802 16836 15824
rect 1104 15750 2916 15802
rect 2968 15750 2980 15802
rect 3032 15750 3044 15802
rect 3096 15750 3108 15802
rect 3160 15750 3172 15802
rect 3224 15750 6849 15802
rect 6901 15750 6913 15802
rect 6965 15750 6977 15802
rect 7029 15750 7041 15802
rect 7093 15750 7105 15802
rect 7157 15750 10782 15802
rect 10834 15750 10846 15802
rect 10898 15750 10910 15802
rect 10962 15750 10974 15802
rect 11026 15750 11038 15802
rect 11090 15750 14715 15802
rect 14767 15750 14779 15802
rect 14831 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 16836 15802
rect 1104 15728 16836 15750
rect 934 15648 940 15700
rect 992 15688 998 15700
rect 1673 15691 1731 15697
rect 1673 15688 1685 15691
rect 992 15660 1685 15688
rect 992 15648 998 15660
rect 1673 15657 1685 15660
rect 1719 15657 1731 15691
rect 1673 15651 1731 15657
rect 16209 15691 16267 15697
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 16666 15688 16672 15700
rect 16255 15660 16672 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 11606 15552 11612 15564
rect 1964 15524 11612 15552
rect 1964 15493 1992 15524
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 13630 15512 13636 15564
rect 13688 15552 13694 15564
rect 16776 15552 16804 15648
rect 13688 15524 13952 15552
rect 13688 15512 13694 15524
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 2924 15456 3249 15484
rect 2924 15444 2930 15456
rect 3237 15453 3249 15456
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 4338 15444 4344 15496
rect 4396 15444 4402 15496
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 7466 15444 7472 15496
rect 7524 15444 7530 15496
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 10560 15456 10793 15484
rect 10560 15444 10566 15456
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 13924 15493 13952 15524
rect 14936 15524 16804 15552
rect 14936 15493 14964 15524
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12124 15456 12357 15484
rect 12124 15444 12130 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 15194 15444 15200 15496
rect 15252 15444 15258 15496
rect 2501 15419 2559 15425
rect 2501 15385 2513 15419
rect 2547 15416 2559 15419
rect 3786 15416 3792 15428
rect 2547 15388 3792 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 15657 15419 15715 15425
rect 15657 15385 15669 15419
rect 15703 15416 15715 15419
rect 15746 15416 15752 15428
rect 15703 15388 15752 15416
rect 15703 15385 15715 15388
rect 15657 15379 15715 15385
rect 15746 15376 15752 15388
rect 15804 15376 15810 15428
rect 15930 15376 15936 15428
rect 15988 15376 15994 15428
rect 2222 15308 2228 15360
rect 2280 15308 2286 15360
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2832 15320 2973 15348
rect 2832 15308 2838 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 2961 15311 3019 15317
rect 3050 15308 3056 15360
rect 3108 15308 3114 15360
rect 4522 15308 4528 15360
rect 4580 15308 4586 15360
rect 6089 15351 6147 15357
rect 6089 15317 6101 15351
rect 6135 15348 6147 15351
rect 6178 15348 6184 15360
rect 6135 15320 6184 15348
rect 6135 15317 6147 15320
rect 6089 15311 6147 15317
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 7650 15308 7656 15360
rect 7708 15308 7714 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 10594 15308 10600 15360
rect 10652 15308 10658 15360
rect 12158 15308 12164 15360
rect 12216 15308 12222 15360
rect 13722 15308 13728 15360
rect 13780 15308 13786 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 15102 15348 15108 15360
rect 15059 15320 15108 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 1104 15258 16995 15280
rect 1104 15206 4882 15258
rect 4934 15206 4946 15258
rect 4998 15206 5010 15258
rect 5062 15206 5074 15258
rect 5126 15206 5138 15258
rect 5190 15206 8815 15258
rect 8867 15206 8879 15258
rect 8931 15206 8943 15258
rect 8995 15206 9007 15258
rect 9059 15206 9071 15258
rect 9123 15206 12748 15258
rect 12800 15206 12812 15258
rect 12864 15206 12876 15258
rect 12928 15206 12940 15258
rect 12992 15206 13004 15258
rect 13056 15206 16681 15258
rect 16733 15206 16745 15258
rect 16797 15206 16809 15258
rect 16861 15206 16873 15258
rect 16925 15206 16937 15258
rect 16989 15206 16995 15258
rect 1104 15184 16995 15206
rect 1486 15104 1492 15156
rect 1544 15104 1550 15156
rect 3050 15104 3056 15156
rect 3108 15104 3114 15156
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 4985 15147 5043 15153
rect 4985 15144 4997 15147
rect 3844 15116 4997 15144
rect 3844 15104 3850 15116
rect 4985 15113 4997 15116
rect 5031 15113 5043 15147
rect 4985 15107 5043 15113
rect 7650 15104 7656 15156
rect 7708 15104 7714 15156
rect 11606 15104 11612 15156
rect 11664 15104 11670 15156
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 15654 15144 15660 15156
rect 13964 15116 15660 15144
rect 13964 15104 13970 15116
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 15746 15104 15752 15156
rect 15804 15104 15810 15156
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16482 15144 16488 15156
rect 16439 15116 16488 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 1118 15036 1124 15088
rect 1176 15076 1182 15088
rect 2866 15076 2872 15088
rect 1176 15048 2872 15076
rect 1176 15036 1182 15048
rect 2866 15036 2872 15048
rect 2924 15036 2930 15088
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 1811 14980 2237 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 15008 2651 15011
rect 3068 15008 3096 15104
rect 2639 14980 3096 15008
rect 5169 15011 5227 15017
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 5718 15008 5724 15020
rect 5215 14980 5724 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 2332 14940 2360 14971
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7668 15008 7696 15104
rect 12158 15036 12164 15088
rect 12216 15036 12222 15088
rect 7515 14980 7696 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 9950 14968 9956 15020
rect 10008 14968 10014 15020
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 12176 15008 12204 15036
rect 11839 14980 12204 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14056 14980 14381 15008
rect 14056 14968 14062 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 14792 14980 14841 15008
rect 14792 14968 14798 14980
rect 14829 14977 14841 14980
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15010 14968 15016 15020
rect 15068 15008 15074 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 15068 14980 15301 15008
rect 15068 14968 15074 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15528 14980 15577 15008
rect 15528 14968 15534 14980
rect 15565 14977 15577 14980
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 8110 14940 8116 14952
rect 2332 14912 8116 14940
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 14461 14943 14519 14949
rect 14461 14909 14473 14943
rect 14507 14940 14519 14943
rect 15930 14940 15936 14952
rect 14507 14912 15936 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 10045 14875 10103 14881
rect 10045 14841 10057 14875
rect 10091 14872 10103 14875
rect 16132 14872 16160 14971
rect 10091 14844 16160 14872
rect 10091 14841 10103 14844
rect 10045 14835 10103 14841
rect 2501 14807 2559 14813
rect 2501 14773 2513 14807
rect 2547 14804 2559 14807
rect 3694 14804 3700 14816
rect 2547 14776 3700 14804
rect 2547 14773 2559 14776
rect 2501 14767 2559 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 7558 14764 7564 14816
rect 7616 14764 7622 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14608 14776 14933 14804
rect 14608 14764 14614 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 15470 14764 15476 14816
rect 15528 14764 15534 14816
rect 1104 14714 16836 14736
rect 1104 14662 2916 14714
rect 2968 14662 2980 14714
rect 3032 14662 3044 14714
rect 3096 14662 3108 14714
rect 3160 14662 3172 14714
rect 3224 14662 6849 14714
rect 6901 14662 6913 14714
rect 6965 14662 6977 14714
rect 7029 14662 7041 14714
rect 7093 14662 7105 14714
rect 7157 14662 10782 14714
rect 10834 14662 10846 14714
rect 10898 14662 10910 14714
rect 10962 14662 10974 14714
rect 11026 14662 11038 14714
rect 11090 14662 14715 14714
rect 14767 14662 14779 14714
rect 14831 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 16836 14714
rect 1104 14640 16836 14662
rect 10594 14600 10600 14612
rect 6886 14572 10600 14600
rect 5718 14424 5724 14476
rect 5776 14464 5782 14476
rect 6886 14464 6914 14572
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 15102 14560 15108 14612
rect 15160 14560 15166 14612
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 15528 14572 16160 14600
rect 15528 14560 15534 14572
rect 15120 14464 15148 14560
rect 5776 14436 6914 14464
rect 14844 14436 15148 14464
rect 5776 14424 5782 14436
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 9214 14396 9220 14408
rect 8803 14368 9220 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 9214 14356 9220 14368
rect 9272 14396 9278 14408
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 9272 14368 9321 14396
rect 9272 14356 9278 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 11514 14396 11520 14408
rect 10643 14368 11520 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12158 14396 12164 14408
rect 12023 14368 12164 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 13722 14396 13728 14408
rect 13403 14368 13728 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 14844 14405 14872 14436
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1397 14331 1455 14337
rect 1397 14328 1409 14331
rect 992 14300 1409 14328
rect 992 14288 998 14300
rect 1397 14297 1409 14300
rect 1443 14297 1455 14331
rect 1397 14291 1455 14297
rect 1765 14331 1823 14337
rect 1765 14297 1777 14331
rect 1811 14328 1823 14331
rect 1811 14300 6914 14328
rect 1811 14297 1823 14300
rect 1765 14291 1823 14297
rect 6886 14260 6914 14300
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 11480 14300 13277 14328
rect 11480 14288 11486 14300
rect 13265 14297 13277 14300
rect 13311 14297 13323 14331
rect 13265 14291 13323 14297
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 15120 14328 15148 14359
rect 15378 14356 15384 14408
rect 15436 14356 15442 14408
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 16132 14405 16160 14572
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 13688 14300 15148 14328
rect 13688 14288 13694 14300
rect 16482 14288 16488 14340
rect 16540 14288 16546 14340
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 6886 14232 8585 14260
rect 8573 14229 8585 14232
rect 8619 14229 8631 14263
rect 8573 14223 8631 14229
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 10042 14260 10048 14272
rect 9447 14232 10048 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 10778 14220 10784 14272
rect 10836 14220 10842 14272
rect 12069 14263 12127 14269
rect 12069 14229 12081 14263
rect 12115 14260 12127 14263
rect 12434 14260 12440 14272
rect 12115 14232 12440 14260
rect 12115 14229 12127 14232
rect 12069 14223 12127 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 14734 14220 14740 14272
rect 14792 14220 14798 14272
rect 15197 14263 15255 14269
rect 15197 14229 15209 14263
rect 15243 14260 15255 14263
rect 15470 14260 15476 14272
rect 15243 14232 15476 14260
rect 15243 14229 15255 14232
rect 15197 14223 15255 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 15562 14220 15568 14272
rect 15620 14220 15626 14272
rect 15746 14220 15752 14272
rect 15804 14220 15810 14272
rect 1104 14170 16995 14192
rect 1104 14118 4882 14170
rect 4934 14118 4946 14170
rect 4998 14118 5010 14170
rect 5062 14118 5074 14170
rect 5126 14118 5138 14170
rect 5190 14118 8815 14170
rect 8867 14118 8879 14170
rect 8931 14118 8943 14170
rect 8995 14118 9007 14170
rect 9059 14118 9071 14170
rect 9123 14118 12748 14170
rect 12800 14118 12812 14170
rect 12864 14118 12876 14170
rect 12928 14118 12940 14170
rect 12992 14118 13004 14170
rect 13056 14118 16681 14170
rect 16733 14118 16745 14170
rect 16797 14118 16809 14170
rect 16861 14118 16873 14170
rect 16925 14118 16937 14170
rect 16989 14118 16995 14170
rect 1104 14096 16995 14118
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 10229 14059 10287 14065
rect 9364 14028 10088 14056
rect 9364 14016 9370 14028
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 6236 13960 9720 13988
rect 6236 13948 6242 13960
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 9030 13880 9036 13932
rect 9088 13880 9094 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9416 13892 9505 13920
rect 1486 13812 1492 13864
rect 1544 13812 1550 13864
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8987 13824 9321 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 9217 13787 9275 13793
rect 9217 13753 9229 13787
rect 9263 13784 9275 13787
rect 9416 13784 9444 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9692 13852 9720 13960
rect 10060 13929 10088 14028
rect 10229 14025 10241 14059
rect 10275 14056 10287 14059
rect 10318 14056 10324 14068
rect 10275 14028 10324 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 10502 14016 10508 14068
rect 10560 14016 10566 14068
rect 10778 14016 10784 14068
rect 10836 14016 10842 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 13817 14059 13875 14065
rect 13817 14025 13829 14059
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 10091 13892 10333 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10520 13920 10548 14016
rect 10796 13988 10824 14016
rect 10796 13960 12480 13988
rect 12452 13929 12480 13960
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 10520 13892 11069 13920
rect 10321 13883 10379 13889
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 12437 13923 12495 13929
rect 11057 13883 11115 13889
rect 11164 13892 11652 13920
rect 11164 13852 11192 13892
rect 9692 13824 11192 13852
rect 11241 13855 11299 13861
rect 11241 13821 11253 13855
rect 11287 13852 11299 13855
rect 11422 13852 11428 13864
rect 11287 13824 11428 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 11624 13852 11652 13892
rect 12437 13889 12449 13923
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13889 12587 13923
rect 12529 13883 12587 13889
rect 12544 13852 12572 13883
rect 12986 13880 12992 13932
rect 13044 13880 13050 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13556 13920 13584 14019
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13556 13892 13645 13920
rect 13357 13883 13415 13889
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13832 13920 13860 14019
rect 14734 14016 14740 14068
rect 14792 14016 14798 14068
rect 15746 14016 15752 14068
rect 15804 14016 15810 14068
rect 14752 13988 14780 14016
rect 14660 13960 14780 13988
rect 15764 13988 15792 14016
rect 16117 13991 16175 13997
rect 16117 13988 16129 13991
rect 15764 13960 16129 13988
rect 14660 13929 14688 13960
rect 16117 13957 16129 13960
rect 16163 13957 16175 13991
rect 16117 13951 16175 13957
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 13832 13892 14473 13920
rect 13633 13883 13691 13889
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15286 13920 15292 13932
rect 14875 13892 15292 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 11624 13824 12572 13852
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12768 13824 13093 13852
rect 12768 13812 12774 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13372 13852 13400 13883
rect 14752 13852 14780 13883
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16390 13920 16396 13932
rect 15427 13892 16396 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 16482 13880 16488 13932
rect 16540 13880 16546 13932
rect 13372 13824 13584 13852
rect 13081 13815 13139 13821
rect 9263 13756 9444 13784
rect 9263 13753 9275 13756
rect 9217 13747 9275 13753
rect 13556 13728 13584 13824
rect 14476 13824 14780 13852
rect 14476 13728 14504 13824
rect 15102 13812 15108 13864
rect 15160 13812 15166 13864
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 9674 13676 9680 13728
rect 9732 13676 9738 13728
rect 10410 13676 10416 13728
rect 10468 13676 10474 13728
rect 10686 13676 10692 13728
rect 10744 13676 10750 13728
rect 12158 13676 12164 13728
rect 12216 13676 12222 13728
rect 12250 13676 12256 13728
rect 12308 13676 12314 13728
rect 12618 13676 12624 13728
rect 12676 13676 12682 13728
rect 12802 13676 12808 13728
rect 12860 13676 12866 13728
rect 13538 13676 13544 13728
rect 13596 13676 13602 13728
rect 14274 13676 14280 13728
rect 14332 13676 14338 13728
rect 14458 13676 14464 13728
rect 14516 13676 14522 13728
rect 1104 13626 16836 13648
rect 1104 13574 2916 13626
rect 2968 13574 2980 13626
rect 3032 13574 3044 13626
rect 3096 13574 3108 13626
rect 3160 13574 3172 13626
rect 3224 13574 6849 13626
rect 6901 13574 6913 13626
rect 6965 13574 6977 13626
rect 7029 13574 7041 13626
rect 7093 13574 7105 13626
rect 7157 13574 10782 13626
rect 10834 13574 10846 13626
rect 10898 13574 10910 13626
rect 10962 13574 10974 13626
rect 11026 13574 11038 13626
rect 11090 13574 14715 13626
rect 14767 13574 14779 13626
rect 14831 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 16836 13626
rect 1104 13552 16836 13574
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9030 13512 9036 13524
rect 8803 13484 9036 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10686 13472 10692 13524
rect 10744 13472 10750 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13044 13484 13461 13512
rect 13044 13472 13050 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 15654 13512 15660 13524
rect 15151 13484 15660 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 10321 13379 10379 13385
rect 9692 13348 10272 13376
rect 9692 13320 9720 13348
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 9306 13308 9312 13320
rect 8619 13280 9312 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 9306 13268 9312 13280
rect 9364 13308 9370 13320
rect 9401 13311 9459 13317
rect 9401 13308 9413 13311
rect 9364 13280 9413 13308
rect 9364 13268 9370 13280
rect 9401 13277 9413 13280
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 10152 13240 10180 13271
rect 8536 13212 10180 13240
rect 10244 13240 10272 13348
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10410 13376 10416 13388
rect 10367 13348 10416 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 10704 13376 10732 13472
rect 11517 13447 11575 13453
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 12345 13447 12403 13453
rect 12345 13444 12357 13447
rect 11563 13416 12357 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 12345 13413 12357 13416
rect 12391 13444 12403 13447
rect 13630 13444 13636 13456
rect 12391 13416 13636 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 14332 13416 15240 13444
rect 14332 13404 14338 13416
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 10704 13348 11805 13376
rect 11793 13345 11805 13348
rect 11839 13345 11851 13379
rect 11793 13339 11851 13345
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 15212 13385 15240 13416
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12860 13348 12909 13376
rect 12860 13336 12866 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 15197 13379 15255 13385
rect 12897 13339 12955 13345
rect 13372 13348 14320 13376
rect 10965 13243 11023 13249
rect 10965 13240 10977 13243
rect 10244 13212 10977 13240
rect 8536 13200 8542 13212
rect 10965 13209 10977 13212
rect 11011 13209 11023 13243
rect 10965 13203 11023 13209
rect 11057 13243 11115 13249
rect 11057 13209 11069 13243
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 9214 13132 9220 13184
rect 9272 13132 9278 13184
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10045 13175 10103 13181
rect 10045 13172 10057 13175
rect 9916 13144 10057 13172
rect 9916 13132 9922 13144
rect 10045 13141 10057 13144
rect 10091 13141 10103 13175
rect 11072 13172 11100 13203
rect 11882 13200 11888 13252
rect 11940 13200 11946 13252
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 12268 13172 12296 13200
rect 11072 13144 12296 13172
rect 10045 13135 10103 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 13372 13181 13400 13348
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13556 13280 13645 13308
rect 13556 13184 13584 13280
rect 13633 13277 13645 13280
rect 13679 13308 13691 13311
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13679 13280 13737 13308
rect 13679 13277 13691 13280
rect 13633 13271 13691 13277
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 14185 13311 14243 13317
rect 14185 13277 14197 13311
rect 14231 13277 14243 13311
rect 14292 13308 14320 13348
rect 15197 13345 15209 13379
rect 15243 13345 15255 13379
rect 15197 13339 15255 13345
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 15344 13348 15393 13376
rect 15344 13336 15350 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 14292 13280 14473 13308
rect 14185 13271 14243 13277
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14200 13240 14228 13271
rect 14642 13268 14648 13320
rect 14700 13268 14706 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15528 13280 16037 13308
rect 15528 13268 15534 13280
rect 16025 13277 16037 13280
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16574 13308 16580 13320
rect 16439 13280 16580 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 14200 13212 14504 13240
rect 14476 13184 14504 13212
rect 13357 13175 13415 13181
rect 13357 13172 13369 13175
rect 12584 13144 13369 13172
rect 12584 13132 12590 13144
rect 13357 13141 13369 13144
rect 13403 13141 13415 13175
rect 13357 13135 13415 13141
rect 13538 13132 13544 13184
rect 13596 13132 13602 13184
rect 13814 13132 13820 13184
rect 13872 13132 13878 13184
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 14458 13132 14464 13184
rect 14516 13132 14522 13184
rect 1104 13082 16995 13104
rect 1104 13030 4882 13082
rect 4934 13030 4946 13082
rect 4998 13030 5010 13082
rect 5062 13030 5074 13082
rect 5126 13030 5138 13082
rect 5190 13030 8815 13082
rect 8867 13030 8879 13082
rect 8931 13030 8943 13082
rect 8995 13030 9007 13082
rect 9059 13030 9071 13082
rect 9123 13030 12748 13082
rect 12800 13030 12812 13082
rect 12864 13030 12876 13082
rect 12928 13030 12940 13082
rect 12992 13030 13004 13082
rect 13056 13030 16681 13082
rect 16733 13030 16745 13082
rect 16797 13030 16809 13082
rect 16861 13030 16873 13082
rect 16925 13030 16937 13082
rect 16989 13030 16995 13082
rect 1104 13008 16995 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 2041 12971 2099 12977
rect 2041 12968 2053 12971
rect 1820 12940 2053 12968
rect 1820 12928 1826 12940
rect 2041 12937 2053 12940
rect 2087 12937 2099 12971
rect 2041 12931 2099 12937
rect 4522 12928 4528 12980
rect 4580 12928 4586 12980
rect 8478 12968 8484 12980
rect 6886 12940 8484 12968
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 3326 12832 3332 12844
rect 2179 12804 3332 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 1780 12764 1808 12795
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 4540 12841 4568 12928
rect 4617 12903 4675 12909
rect 4617 12869 4629 12903
rect 4663 12900 4675 12903
rect 5350 12900 5356 12912
rect 4663 12872 5356 12900
rect 4663 12869 4675 12872
rect 4617 12863 4675 12869
rect 5350 12860 5356 12872
rect 5408 12900 5414 12912
rect 6886 12900 6914 12940
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 9214 12928 9220 12980
rect 9272 12928 9278 12980
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 9674 12968 9680 12980
rect 9539 12940 9680 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11882 12968 11888 12980
rect 11195 12940 11888 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 14366 12928 14372 12980
rect 14424 12928 14430 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 15289 12971 15347 12977
rect 15289 12968 15301 12971
rect 14700 12940 15301 12968
rect 14700 12928 14706 12940
rect 15289 12937 15301 12940
rect 15335 12937 15347 12971
rect 15289 12931 15347 12937
rect 5408 12872 6914 12900
rect 5408 12860 5414 12872
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 6178 12832 6184 12844
rect 5491 12804 6184 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9232 12832 9260 12928
rect 11784 12903 11842 12909
rect 9692 12872 11560 12900
rect 9692 12844 9720 12872
rect 9079 12804 9260 12832
rect 9585 12835 9643 12841
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9858 12841 9864 12844
rect 9852 12832 9864 12841
rect 9819 12804 9864 12832
rect 9852 12795 9864 12804
rect 9858 12792 9864 12795
rect 9916 12792 9922 12844
rect 11532 12841 11560 12872
rect 11784 12869 11796 12903
rect 11830 12900 11842 12903
rect 12158 12900 12164 12912
rect 11830 12872 12164 12900
rect 11830 12869 11842 12872
rect 11784 12863 11842 12869
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 1780 12736 5304 12764
rect 5276 12705 5304 12736
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 8536 12736 8861 12764
rect 8536 12724 8542 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8849 12727 8907 12733
rect 5261 12699 5319 12705
rect 5261 12665 5273 12699
rect 5307 12665 5319 12699
rect 5261 12659 5319 12665
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12696 11023 12699
rect 11072 12696 11100 12795
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 13630 12832 13636 12844
rect 12676 12804 13636 12832
rect 12676 12792 12682 12804
rect 13630 12792 13636 12804
rect 13688 12832 13694 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13688 12804 13737 12832
rect 13688 12792 13694 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13832 12832 13860 12928
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13832 12804 13921 12832
rect 13725 12795 13783 12801
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 14384 12832 14412 12928
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 16114 12900 16120 12912
rect 15795 12872 16120 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 14384 12804 15485 12832
rect 13909 12795 13967 12801
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 13538 12764 13544 12776
rect 12912 12736 13544 12764
rect 11514 12696 11520 12708
rect 11011 12668 11520 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 934 12588 940 12640
rect 992 12628 998 12640
rect 1489 12631 1547 12637
rect 1489 12628 1501 12631
rect 992 12600 1501 12628
rect 992 12588 998 12600
rect 1489 12597 1501 12600
rect 1535 12597 1547 12631
rect 1489 12591 1547 12597
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 12912 12637 12940 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14240 12736 15025 12764
rect 14240 12724 14246 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15252 12736 15669 12764
rect 15252 12724 15258 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15896 12736 15945 12764
rect 15896 12724 15902 12736
rect 15933 12733 15945 12736
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 14274 12656 14280 12708
rect 14332 12656 14338 12708
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12676 12600 12909 12628
rect 12676 12588 12682 12600
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 12897 12591 12955 12597
rect 12986 12588 12992 12640
rect 13044 12588 13050 12640
rect 14458 12588 14464 12640
rect 14516 12588 14522 12640
rect 1104 12538 16836 12560
rect 1104 12486 2916 12538
rect 2968 12486 2980 12538
rect 3032 12486 3044 12538
rect 3096 12486 3108 12538
rect 3160 12486 3172 12538
rect 3224 12486 6849 12538
rect 6901 12486 6913 12538
rect 6965 12486 6977 12538
rect 7029 12486 7041 12538
rect 7093 12486 7105 12538
rect 7157 12486 10782 12538
rect 10834 12486 10846 12538
rect 10898 12486 10910 12538
rect 10962 12486 10974 12538
rect 11026 12486 11038 12538
rect 11090 12486 14715 12538
rect 14767 12486 14779 12538
rect 14831 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 16836 12538
rect 1104 12464 16836 12486
rect 8941 12427 8999 12433
rect 8941 12393 8953 12427
rect 8987 12424 8999 12427
rect 9306 12424 9312 12436
rect 8987 12396 9312 12424
rect 8987 12393 8999 12396
rect 8941 12387 8999 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 12526 12424 12532 12436
rect 12483 12396 12532 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 14366 12424 14372 12436
rect 13955 12396 14372 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 7650 12248 7656 12300
rect 7708 12248 7714 12300
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 12526 12288 12532 12300
rect 10367 12260 12532 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 4522 12220 4528 12232
rect 2179 12192 4528 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 6972 12192 7849 12220
rect 6972 12180 6978 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10336 12220 10364 12251
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 15620 12260 16528 12288
rect 15620 12248 15626 12260
rect 9732 12192 10364 12220
rect 10597 12223 10655 12229
rect 9732 12180 9738 12192
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 10643 12192 11161 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 934 12112 940 12164
rect 992 12152 998 12164
rect 1397 12155 1455 12161
rect 1397 12152 1409 12155
rect 992 12124 1409 12152
rect 992 12112 998 12124
rect 1397 12121 1409 12124
rect 1443 12121 1455 12155
rect 1397 12115 1455 12121
rect 1765 12155 1823 12161
rect 1765 12121 1777 12155
rect 1811 12152 1823 12155
rect 10076 12155 10134 12161
rect 1811 12124 1992 12152
rect 1811 12121 1823 12124
rect 1765 12115 1823 12121
rect 1964 12093 1992 12124
rect 10076 12121 10088 12155
rect 10122 12152 10134 12155
rect 10318 12152 10324 12164
rect 10122 12124 10324 12152
rect 10122 12121 10134 12124
rect 10076 12115 10134 12121
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 11164 12152 11192 12183
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11664 12192 11805 12220
rect 11664 12180 11670 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 12544 12220 12572 12248
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 12544 12192 15485 12220
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 15654 12220 15660 12232
rect 15519 12192 15660 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 16500 12229 16528 12260
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12189 16543 12223
rect 16485 12183 16543 12189
rect 12796 12155 12854 12161
rect 11164 12124 12434 12152
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7524 12056 8309 12084
rect 7524 12044 7530 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8297 12047 8355 12053
rect 10502 12044 10508 12096
rect 10560 12044 10566 12096
rect 11330 12044 11336 12096
rect 11388 12044 11394 12096
rect 12406 12084 12434 12124
rect 12796 12121 12808 12155
rect 12842 12152 12854 12155
rect 12986 12152 12992 12164
rect 12842 12124 12992 12152
rect 12842 12121 12854 12124
rect 12796 12115 12854 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 15228 12155 15286 12161
rect 15228 12121 15240 12155
rect 15274 12152 15286 12155
rect 15565 12155 15623 12161
rect 15565 12152 15577 12155
rect 15274 12124 15577 12152
rect 15274 12121 15286 12124
rect 15228 12115 15286 12121
rect 15565 12121 15577 12124
rect 15611 12121 15623 12155
rect 15565 12115 15623 12121
rect 14090 12084 14096 12096
rect 12406 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 16132 12084 16160 12183
rect 14424 12056 16160 12084
rect 14424 12044 14430 12056
rect 16298 12044 16304 12096
rect 16356 12044 16362 12096
rect 1104 11994 16995 12016
rect 1104 11942 4882 11994
rect 4934 11942 4946 11994
rect 4998 11942 5010 11994
rect 5062 11942 5074 11994
rect 5126 11942 5138 11994
rect 5190 11942 8815 11994
rect 8867 11942 8879 11994
rect 8931 11942 8943 11994
rect 8995 11942 9007 11994
rect 9059 11942 9071 11994
rect 9123 11942 12748 11994
rect 12800 11942 12812 11994
rect 12864 11942 12876 11994
rect 12928 11942 12940 11994
rect 12992 11942 13004 11994
rect 13056 11942 16681 11994
rect 16733 11942 16745 11994
rect 16797 11942 16809 11994
rect 16861 11942 16873 11994
rect 16925 11942 16937 11994
rect 16989 11942 16995 11994
rect 1104 11920 16995 11942
rect 6914 11840 6920 11892
rect 6972 11840 6978 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11849 7067 11883
rect 7009 11843 7067 11849
rect 8665 11883 8723 11889
rect 8665 11849 8677 11883
rect 8711 11880 8723 11883
rect 9122 11880 9128 11892
rect 8711 11852 9128 11880
rect 8711 11849 8723 11852
rect 8665 11843 8723 11849
rect 5718 11704 5724 11756
rect 5776 11704 5782 11756
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 7024 11744 7052 11843
rect 9122 11840 9128 11852
rect 9180 11880 9186 11892
rect 9180 11852 9812 11880
rect 9180 11840 9186 11852
rect 7466 11772 7472 11824
rect 7524 11812 7530 11824
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 7524 11784 8953 11812
rect 7524 11772 7530 11784
rect 8941 11781 8953 11784
rect 8987 11781 8999 11815
rect 8941 11775 8999 11781
rect 9030 11772 9036 11824
rect 9088 11772 9094 11824
rect 6779 11716 7052 11744
rect 7193 11747 7251 11753
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 7374 11744 7380 11756
rect 7239 11716 7380 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7558 11753 7564 11756
rect 7552 11707 7564 11753
rect 7558 11704 7564 11707
rect 7616 11704 7622 11756
rect 9784 11753 9812 11852
rect 10318 11840 10324 11892
rect 10376 11840 10382 11892
rect 10502 11840 10508 11892
rect 10560 11840 10566 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12621 11883 12679 11889
rect 12621 11880 12633 11883
rect 12032 11852 12633 11880
rect 12032 11840 12038 11852
rect 12621 11849 12633 11852
rect 12667 11849 12679 11883
rect 12621 11843 12679 11849
rect 15378 11840 15384 11892
rect 15436 11840 15442 11892
rect 10520 11812 10548 11840
rect 14268 11815 14326 11821
rect 10520 11784 10916 11812
rect 10888 11753 10916 11784
rect 12544 11784 14044 11812
rect 12544 11756 12572 11784
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11744 9827 11747
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 9815 11716 10609 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 14016 11753 14044 11784
rect 14268 11781 14280 11815
rect 14314 11812 14326 11815
rect 14458 11812 14464 11824
rect 14314 11784 14464 11812
rect 14314 11781 14326 11784
rect 14268 11775 14326 11781
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 15396 11744 15424 11840
rect 16206 11744 16212 11756
rect 15396 11716 16212 11744
rect 14001 11707 14059 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6512 11648 7297 11676
rect 6512 11636 6518 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 10134 11676 10140 11688
rect 9631 11648 10140 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10284 11648 10701 11676
rect 10284 11636 10290 11648
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 11514 11636 11520 11688
rect 11572 11636 11578 11688
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13320 11648 13737 11676
rect 13320 11636 13326 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 11974 11608 11980 11620
rect 9600 11580 11980 11608
rect 5626 11500 5632 11552
rect 5684 11500 5690 11552
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 9600 11540 9628 11580
rect 11974 11568 11980 11580
rect 12032 11568 12038 11620
rect 8260 11512 9628 11540
rect 8260 11500 8266 11512
rect 10410 11500 10416 11552
rect 10468 11500 10474 11552
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11379 11512 11897 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11885 11509 11897 11512
rect 11931 11540 11943 11543
rect 15194 11540 15200 11552
rect 11931 11512 15200 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15620 11512 15669 11540
rect 15620 11500 15626 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 15657 11503 15715 11509
rect 1104 11450 16836 11472
rect 1104 11398 2916 11450
rect 2968 11398 2980 11450
rect 3032 11398 3044 11450
rect 3096 11398 3108 11450
rect 3160 11398 3172 11450
rect 3224 11398 6849 11450
rect 6901 11398 6913 11450
rect 6965 11398 6977 11450
rect 7029 11398 7041 11450
rect 7093 11398 7105 11450
rect 7157 11398 10782 11450
rect 10834 11398 10846 11450
rect 10898 11398 10910 11450
rect 10962 11398 10974 11450
rect 11026 11398 11038 11450
rect 11090 11398 14715 11450
rect 14767 11398 14779 11450
rect 14831 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 16836 11450
rect 1104 11376 16836 11398
rect 5626 11296 5632 11348
rect 5684 11296 5690 11348
rect 7466 11296 7472 11348
rect 7524 11296 7530 11348
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 9030 11296 9036 11348
rect 9088 11296 9094 11348
rect 9122 11296 9128 11348
rect 9180 11296 9186 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 11330 11296 11336 11348
rect 11388 11296 11394 11348
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 15712 11308 16068 11336
rect 15712 11296 15718 11308
rect 2225 11271 2283 11277
rect 2225 11237 2237 11271
rect 2271 11237 2283 11271
rect 2225 11231 2283 11237
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2240 11132 2268 11231
rect 5644 11209 5672 11296
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 5675 11172 6101 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6914 11200 6920 11212
rect 6319 11172 6920 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 7055 11172 8585 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 8573 11169 8585 11172
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 1811 11104 2268 11132
rect 2409 11135 2467 11141
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2774 11132 2780 11144
rect 2455 11104 2780 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2832 11104 2973 11132
rect 2832 11092 2838 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 4764 11104 5457 11132
rect 4764 11092 4770 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 5445 11095 5503 11101
rect 6380 11104 6837 11132
rect 1394 11024 1400 11076
rect 1452 11024 1458 11076
rect 3053 11067 3111 11073
rect 3053 11033 3065 11067
rect 3099 11064 3111 11067
rect 6380 11064 6408 11104
rect 6825 11101 6837 11104
rect 6871 11132 6883 11135
rect 6871 11104 7420 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 3099 11036 6408 11064
rect 6733 11067 6791 11073
rect 3099 11033 3111 11036
rect 3053 11027 3111 11033
rect 6733 11033 6745 11067
rect 6779 11064 6791 11067
rect 7392 11064 7420 11104
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 9140 11141 9168 11296
rect 10428 11200 10456 11296
rect 9600 11172 10456 11200
rect 9600 11141 9628 11172
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 7524 11104 8217 11132
rect 7524 11092 7530 11104
rect 8205 11101 8217 11104
rect 8251 11132 8263 11135
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 8251 11104 8677 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8665 11101 8677 11104
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11348 11132 11376 11296
rect 11195 11104 11376 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 8294 11064 8300 11076
rect 6779 11036 7052 11064
rect 7392 11036 8300 11064
rect 6779 11033 6791 11036
rect 6733 11027 6791 11033
rect 7024 11008 7052 11036
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 8680 11064 8708 11095
rect 9493 11067 9551 11073
rect 8680 11036 9260 11064
rect 9232 11008 9260 11036
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9674 11064 9680 11076
rect 9539 11036 9680 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 9950 11024 9956 11076
rect 10008 11024 10014 11076
rect 10045 11067 10103 11073
rect 10045 11033 10057 11067
rect 10091 11033 10103 11067
rect 10045 11027 10103 11033
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 4985 10999 5043 11005
rect 4985 10996 4997 10999
rect 4856 10968 4997 10996
rect 4856 10956 4862 10968
rect 4985 10965 4997 10968
rect 5031 10965 5043 10999
rect 4985 10959 5043 10965
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 9214 10956 9220 11008
rect 9272 10956 9278 11008
rect 9769 10999 9827 11005
rect 9769 10965 9781 10999
rect 9815 10996 9827 10999
rect 10060 10996 10088 11027
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 10597 11067 10655 11073
rect 10597 11064 10609 11067
rect 10192 11036 10609 11064
rect 10192 11024 10198 11036
rect 10597 11033 10609 11036
rect 10643 11064 10655 11067
rect 10686 11064 10692 11076
rect 10643 11036 10692 11064
rect 10643 11033 10655 11036
rect 10597 11027 10655 11033
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 11716 11064 11744 11296
rect 13906 11228 13912 11280
rect 13964 11228 13970 11280
rect 11974 11160 11980 11212
rect 12032 11160 12038 11212
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 12667 11172 13553 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13541 11169 13553 11172
rect 13587 11200 13599 11203
rect 13924 11200 13952 11228
rect 16040 11209 16068 11308
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16172 11308 16221 11336
rect 16172 11296 16178 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 13587 11172 13952 11200
rect 16025 11203 16083 11209
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 16025 11169 16037 11203
rect 16071 11169 16083 11203
rect 16206 11200 16212 11212
rect 16025 11163 16083 11169
rect 16132 11172 16212 11200
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 13078 11132 13084 11144
rect 12943 11104 13084 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 16132 11141 16160 11172
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 11348 11036 11744 11064
rect 11348 11005 11376 11036
rect 12066 11024 12072 11076
rect 12124 11024 12130 11076
rect 13722 11024 13728 11076
rect 13780 11024 13786 11076
rect 13817 11067 13875 11073
rect 13817 11033 13829 11067
rect 13863 11033 13875 11067
rect 13817 11027 13875 11033
rect 9815 10968 10088 10996
rect 11333 10999 11391 11005
rect 9815 10965 9827 10968
rect 9769 10959 9827 10965
rect 11333 10965 11345 10999
rect 11379 10965 11391 10999
rect 11333 10959 11391 10965
rect 13081 10999 13139 11005
rect 13081 10965 13093 10999
rect 13127 10996 13139 10999
rect 13354 10996 13360 11008
rect 13127 10968 13360 10996
rect 13127 10965 13139 10968
rect 13081 10959 13139 10965
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 13832 10996 13860 11027
rect 14182 11024 14188 11076
rect 14240 11024 14246 11076
rect 14550 11024 14556 11076
rect 14608 11024 14614 11076
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 15758 11067 15816 11073
rect 15758 11064 15770 11067
rect 15620 11036 15770 11064
rect 15620 11024 15626 11036
rect 15758 11033 15770 11036
rect 15804 11033 15816 11067
rect 15758 11027 15816 11033
rect 13906 10996 13912 11008
rect 13832 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14366 10956 14372 11008
rect 14424 10996 14430 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 14424 10968 14657 10996
rect 14424 10956 14430 10968
rect 14645 10965 14657 10968
rect 14691 10965 14703 10999
rect 14645 10959 14703 10965
rect 1104 10906 16995 10928
rect 1104 10854 4882 10906
rect 4934 10854 4946 10906
rect 4998 10854 5010 10906
rect 5062 10854 5074 10906
rect 5126 10854 5138 10906
rect 5190 10854 8815 10906
rect 8867 10854 8879 10906
rect 8931 10854 8943 10906
rect 8995 10854 9007 10906
rect 9059 10854 9071 10906
rect 9123 10854 12748 10906
rect 12800 10854 12812 10906
rect 12864 10854 12876 10906
rect 12928 10854 12940 10906
rect 12992 10854 13004 10906
rect 13056 10854 16681 10906
rect 16733 10854 16745 10906
rect 16797 10854 16809 10906
rect 16861 10854 16873 10906
rect 16925 10854 16937 10906
rect 16989 10854 16995 10906
rect 1104 10832 16995 10854
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 4798 10752 4804 10804
rect 4856 10752 4862 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7193 10795 7251 10801
rect 7193 10792 7205 10795
rect 6972 10764 7205 10792
rect 6972 10752 6978 10764
rect 7193 10761 7205 10764
rect 7239 10761 7251 10795
rect 7193 10755 7251 10761
rect 7466 10752 7472 10804
rect 7524 10752 7530 10804
rect 8202 10752 8208 10804
rect 8260 10752 8266 10804
rect 8312 10764 11284 10792
rect 7006 10684 7012 10736
rect 7064 10724 7070 10736
rect 8220 10724 8248 10752
rect 7064 10696 8248 10724
rect 7064 10684 7070 10696
rect 1762 10616 1768 10668
rect 1820 10616 1826 10668
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10625 4307 10659
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4249 10619 4307 10625
rect 4448 10628 4537 10656
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 992 10424 1501 10452
rect 992 10412 998 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 4264 10452 4292 10619
rect 4448 10529 4476 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5307 10628 5641 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5442 10548 5448 10600
rect 5500 10548 5506 10600
rect 4433 10523 4491 10529
rect 4433 10489 4445 10523
rect 4479 10489 4491 10523
rect 5736 10520 5764 10619
rect 5994 10616 6000 10668
rect 6052 10616 6058 10668
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6696 10628 7297 10656
rect 6696 10616 6702 10628
rect 7285 10625 7297 10628
rect 7331 10656 7343 10659
rect 8312 10656 8340 10764
rect 9508 10696 10548 10724
rect 9508 10668 9536 10696
rect 7331 10628 8340 10656
rect 8593 10659 8651 10665
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 8593 10625 8605 10659
rect 8639 10656 8651 10659
rect 8938 10656 8944 10668
rect 8639 10628 8944 10656
rect 8639 10625 8651 10628
rect 8593 10619 8651 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9122 10656 9128 10668
rect 9079 10628 9128 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10520 10665 10548 10696
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 9732 10628 10333 10656
rect 9732 10616 9738 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 11256 10656 11284 10764
rect 12066 10752 12072 10804
rect 12124 10752 12130 10804
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10761 12587 10795
rect 12529 10755 12587 10761
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 13078 10792 13084 10804
rect 12851 10764 13084 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 12544 10724 12572 10755
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 16298 10752 16304 10804
rect 16356 10752 16362 10804
rect 13814 10724 13820 10736
rect 12544 10696 12940 10724
rect 12161 10659 12219 10665
rect 11256 10628 12112 10656
rect 10505 10619 10563 10625
rect 6362 10548 6368 10600
rect 6420 10548 6426 10600
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10588 8907 10591
rect 9858 10588 9864 10600
rect 8895 10560 9864 10588
rect 8895 10557 8907 10560
rect 8849 10551 8907 10557
rect 4433 10483 4491 10489
rect 4540 10492 5764 10520
rect 4540 10464 4568 10492
rect 4522 10452 4528 10464
rect 4264 10424 4528 10452
rect 1489 10415 1547 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 5736 10452 5764 10492
rect 6181 10523 6239 10529
rect 6181 10489 6193 10523
rect 6227 10520 6239 10523
rect 6564 10520 6592 10551
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 11974 10588 11980 10600
rect 10275 10560 11980 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 6227 10492 6592 10520
rect 9125 10523 9183 10529
rect 6227 10489 6239 10492
rect 6181 10483 6239 10489
rect 9125 10489 9137 10523
rect 9171 10520 9183 10523
rect 10060 10520 10088 10551
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 12084 10588 12112 10628
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12250 10656 12256 10668
rect 12207 10628 12256 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 12912 10665 12940 10696
rect 13004 10696 13820 10724
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12308 10628 12357 10656
rect 12308 10616 12314 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12621 10659 12679 10665
rect 12621 10625 12633 10659
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12636 10588 12664 10619
rect 13004 10588 13032 10696
rect 13814 10684 13820 10696
rect 13872 10724 13878 10736
rect 14366 10724 14372 10736
rect 13872 10696 14372 10724
rect 13872 10684 13878 10696
rect 14366 10684 14372 10696
rect 14424 10724 14430 10736
rect 14424 10696 14780 10724
rect 14424 10684 14430 10696
rect 13262 10616 13268 10668
rect 13320 10616 13326 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 14752 10665 14780 10696
rect 15746 10684 15752 10736
rect 15804 10684 15810 10736
rect 15841 10727 15899 10733
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 16316 10724 16344 10752
rect 15887 10696 16344 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13412 10628 13461 10656
rect 13412 10616 13418 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 13722 10588 13728 10600
rect 12084 10560 13032 10588
rect 13096 10560 13728 10588
rect 13096 10529 13124 10560
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 14826 10548 14832 10600
rect 14884 10548 14890 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 9171 10492 10088 10520
rect 13081 10523 13139 10529
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 13081 10489 13093 10523
rect 13127 10489 13139 10523
rect 13081 10483 13139 10489
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 13596 10492 14105 10520
rect 13596 10480 13602 10492
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 14093 10483 14151 10489
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 15028 10520 15056 10551
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15988 10560 16037 10588
rect 15988 10548 15994 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 14424 10492 15056 10520
rect 14424 10480 14430 10492
rect 7374 10452 7380 10464
rect 5736 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9490 10412 9496 10464
rect 9548 10412 9554 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 9950 10452 9956 10464
rect 9907 10424 9956 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 9950 10412 9956 10424
rect 10008 10452 10014 10464
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10008 10424 10701 10452
rect 10008 10412 10014 10424
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 13964 10424 15209 10452
rect 13964 10412 13970 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 1104 10362 16836 10384
rect 1104 10310 2916 10362
rect 2968 10310 2980 10362
rect 3032 10310 3044 10362
rect 3096 10310 3108 10362
rect 3160 10310 3172 10362
rect 3224 10310 6849 10362
rect 6901 10310 6913 10362
rect 6965 10310 6977 10362
rect 7029 10310 7041 10362
rect 7093 10310 7105 10362
rect 7157 10310 10782 10362
rect 10834 10310 10846 10362
rect 10898 10310 10910 10362
rect 10962 10310 10974 10362
rect 11026 10310 11038 10362
rect 11090 10310 14715 10362
rect 14767 10310 14779 10362
rect 14831 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 16836 10362
rect 1104 10288 16836 10310
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6052 10220 6561 10248
rect 6052 10208 6058 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 8938 10208 8944 10260
rect 8996 10208 9002 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9364 10220 9965 10248
rect 9364 10208 9370 10220
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 12526 10248 12532 10260
rect 9953 10211 10011 10217
rect 11716 10220 12532 10248
rect 6457 10183 6515 10189
rect 6457 10149 6469 10183
rect 6503 10180 6515 10183
rect 6638 10180 6644 10192
rect 6503 10152 6644 10180
rect 6503 10149 6515 10152
rect 6457 10143 6515 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 6880 10152 8064 10180
rect 6880 10140 6886 10152
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4856 10084 4905 10112
rect 4856 10072 4862 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 6546 10072 6552 10124
rect 6604 10112 6610 10124
rect 8036 10121 8064 10152
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 11716 10189 11744 10220
rect 12526 10208 12532 10220
rect 12584 10248 12590 10260
rect 13817 10251 13875 10257
rect 12584 10220 13676 10248
rect 12584 10208 12590 10220
rect 11701 10183 11759 10189
rect 11701 10180 11713 10183
rect 9916 10152 11713 10180
rect 9916 10140 9922 10152
rect 11701 10149 11713 10152
rect 11747 10149 11759 10183
rect 11701 10143 11759 10149
rect 13648 10124 13676 10220
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 14366 10248 14372 10260
rect 13863 10220 14372 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 8021 10115 8079 10121
rect 6604 10084 6684 10112
rect 6604 10072 6610 10084
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 2832 10016 3801 10044
rect 2832 10004 2838 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 4764 10016 5089 10044
rect 4764 10004 4770 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5810 10004 5816 10056
rect 5868 10046 5874 10056
rect 5868 10018 5911 10046
rect 5868 10004 5874 10018
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6270 10004 6276 10056
rect 6328 10004 6334 10056
rect 6656 10040 6684 10084
rect 8021 10081 8033 10115
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8168 10084 12664 10112
rect 8168 10072 8174 10084
rect 6725 10043 6783 10049
rect 6725 10040 6737 10043
rect 6656 10012 6737 10040
rect 6725 10009 6737 10012
rect 6771 10009 6783 10043
rect 6725 10003 6783 10009
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10020 6883 10047
rect 8205 10047 8263 10053
rect 6871 10013 6914 10020
rect 6825 10007 6914 10013
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8251 10016 8309 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 6840 9992 6914 10007
rect 8386 10004 8392 10056
rect 8444 10044 8450 10056
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 8444 10016 8769 10044
rect 8444 10004 8450 10016
rect 8757 10013 8769 10016
rect 8803 10044 8815 10047
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 8803 10016 9505 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 5258 9868 5264 9920
rect 5316 9908 5322 9920
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 5316 9880 5549 9908
rect 5316 9868 5322 9880
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 5537 9871 5595 9877
rect 5718 9868 5724 9920
rect 5776 9868 5782 9920
rect 5902 9868 5908 9920
rect 5960 9868 5966 9920
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6886 9908 6914 9992
rect 7469 9979 7527 9985
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 8662 9976 8668 9988
rect 7515 9948 8668 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 8662 9936 8668 9948
rect 8720 9936 8726 9988
rect 9122 9936 9128 9988
rect 9180 9976 9186 9988
rect 10152 9976 10180 10007
rect 9180 9948 10180 9976
rect 9180 9936 9186 9948
rect 10410 9936 10416 9988
rect 10468 9936 10474 9988
rect 12636 9976 12664 10084
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 13814 10112 13820 10124
rect 13740 10084 13820 10112
rect 13377 10047 13435 10053
rect 13377 10013 13389 10047
rect 13423 10040 13435 10047
rect 13538 10044 13544 10056
rect 13464 10040 13544 10044
rect 13423 10016 13544 10040
rect 13423 10013 13492 10016
rect 13377 10012 13492 10013
rect 13377 10007 13435 10012
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13740 10053 13768 10084
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 14090 10072 14096 10124
rect 14148 10072 14154 10124
rect 14458 10072 14464 10124
rect 14516 10112 14522 10124
rect 14829 10115 14887 10121
rect 14829 10112 14841 10115
rect 14516 10084 14841 10112
rect 14516 10072 14522 10084
rect 14829 10081 14841 10084
rect 14875 10081 14887 10115
rect 14829 10075 14887 10081
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15712 10084 16313 10112
rect 15712 10072 15718 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 13262 9976 13268 9988
rect 12636 9948 13268 9976
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 15286 9976 15292 9988
rect 13556 9948 15292 9976
rect 13556 9920 13584 9948
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 15657 9979 15715 9985
rect 15657 9976 15669 9979
rect 15344 9948 15669 9976
rect 15344 9936 15350 9948
rect 15657 9945 15669 9948
rect 15703 9945 15715 9979
rect 15657 9939 15715 9945
rect 16206 9936 16212 9988
rect 16264 9936 16270 9988
rect 6052 9880 6914 9908
rect 6052 9868 6058 9880
rect 7558 9868 7564 9920
rect 7616 9868 7622 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9824 9880 9873 9908
rect 9824 9868 9830 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 12250 9868 12256 9920
rect 12308 9868 12314 9920
rect 13538 9868 13544 9920
rect 13596 9868 13602 9920
rect 15470 9868 15476 9920
rect 15528 9868 15534 9920
rect 1104 9818 16995 9840
rect 1104 9766 4882 9818
rect 4934 9766 4946 9818
rect 4998 9766 5010 9818
rect 5062 9766 5074 9818
rect 5126 9766 5138 9818
rect 5190 9766 8815 9818
rect 8867 9766 8879 9818
rect 8931 9766 8943 9818
rect 8995 9766 9007 9818
rect 9059 9766 9071 9818
rect 9123 9766 12748 9818
rect 12800 9766 12812 9818
rect 12864 9766 12876 9818
rect 12928 9766 12940 9818
rect 12992 9766 13004 9818
rect 13056 9766 16681 9818
rect 16733 9766 16745 9818
rect 16797 9766 16809 9818
rect 16861 9766 16873 9818
rect 16925 9766 16937 9818
rect 16989 9766 16995 9818
rect 1104 9744 16995 9766
rect 5460 9676 5856 9704
rect 5460 9648 5488 9676
rect 4148 9639 4206 9645
rect 4148 9605 4160 9639
rect 4194 9636 4206 9639
rect 4430 9636 4436 9648
rect 4194 9608 4436 9636
rect 4194 9605 4206 9608
rect 4148 9599 4206 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 5442 9596 5448 9648
rect 5500 9596 5506 9648
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 5718 9636 5724 9648
rect 5583 9608 5724 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 5828 9636 5856 9676
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 7282 9704 7288 9716
rect 6328 9676 7288 9704
rect 6328 9664 6334 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 8570 9704 8576 9716
rect 8220 9676 8576 9704
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 5828 9608 6101 9636
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 6089 9599 6147 9605
rect 3533 9571 3591 9577
rect 3533 9537 3545 9571
rect 3579 9568 3591 9571
rect 4982 9568 4988 9580
rect 3579 9540 4988 9568
rect 3579 9537 3591 9540
rect 3533 9531 3591 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 6454 9568 6460 9580
rect 6411 9540 6460 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3835 9472 3893 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 2774 9432 2780 9444
rect 2455 9404 2780 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 2774 9392 2780 9404
rect 2832 9392 2838 9444
rect 3896 9364 3924 9463
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5316 9472 5457 9500
rect 5316 9460 5322 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 6380 9500 6408 9531
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6632 9571 6690 9577
rect 6632 9537 6644 9571
rect 6678 9568 6690 9571
rect 7190 9568 7196 9580
rect 6678 9540 7196 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8220 9568 8248 9676
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 14461 9707 14519 9713
rect 13096 9676 13492 9704
rect 13096 9648 13124 9676
rect 13464 9674 13492 9676
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8352 9608 8432 9636
rect 8352 9596 8358 9608
rect 7883 9540 8248 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 5445 9463 5503 9469
rect 5552 9472 6408 9500
rect 7576 9500 7604 9528
rect 7926 9500 7932 9512
rect 7576 9472 7932 9500
rect 5552 9432 5580 9472
rect 7926 9460 7932 9472
rect 7984 9500 7990 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7984 9472 8125 9500
rect 7984 9460 7990 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9469 8355 9503
rect 8404 9500 8432 9608
rect 8662 9596 8668 9648
rect 8720 9636 8726 9648
rect 10198 9639 10256 9645
rect 10198 9636 10210 9639
rect 8720 9608 10210 9636
rect 8720 9596 8726 9608
rect 10198 9605 10210 9608
rect 10244 9605 10256 9639
rect 13078 9636 13084 9648
rect 10198 9599 10256 9605
rect 11624 9608 13084 9636
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9171 9540 9628 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 8404 9472 9229 9500
rect 8297 9463 8355 9469
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 4816 9404 5580 9432
rect 4816 9364 4844 9404
rect 5718 9392 5724 9444
rect 5776 9392 5782 9444
rect 8021 9435 8079 9441
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8312 9432 8340 9463
rect 8067 9404 8340 9432
rect 9033 9435 9091 9441
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 9033 9401 9045 9435
rect 9079 9432 9091 9435
rect 9416 9432 9444 9463
rect 9079 9404 9444 9432
rect 9079 9401 9091 9404
rect 9033 9395 9091 9401
rect 3896 9336 4844 9364
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 5736 9364 5764 9392
rect 9600 9376 9628 9540
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 11624 9577 11652 9608
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 13170 9596 13176 9648
rect 13228 9645 13234 9648
rect 13464 9646 13584 9674
rect 14461 9673 14473 9707
rect 14507 9704 14519 9707
rect 15010 9704 15016 9716
rect 14507 9676 15016 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 16356 9676 16436 9704
rect 16356 9664 16362 9676
rect 13228 9639 13262 9645
rect 13250 9605 13262 9639
rect 13228 9599 13262 9605
rect 13228 9596 13234 9599
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9916 9540 9965 9568
rect 9916 9528 9922 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 11609 9571 11667 9577
rect 11609 9537 11621 9571
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 13354 9568 13360 9580
rect 11747 9540 13360 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 11624 9432 11652 9531
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9469 13507 9503
rect 13556 9500 13584 9646
rect 16408 9645 16436 9676
rect 16393 9639 16451 9645
rect 16393 9605 16405 9639
rect 16439 9605 16451 9639
rect 16393 9599 16451 9605
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 14369 9571 14427 9577
rect 13688 9540 14228 9568
rect 13688 9528 13694 9540
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 13556 9472 14105 9500
rect 13449 9463 13507 9469
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14200 9500 14228 9540
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14550 9568 14556 9580
rect 14415 9540 14556 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14912 9571 14970 9577
rect 14912 9537 14924 9571
rect 14958 9568 14970 9571
rect 15194 9568 15200 9580
rect 14958 9540 15200 9568
rect 14958 9537 14970 9540
rect 14912 9531 14970 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 14200 9472 14657 9500
rect 14093 9463 14151 9469
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 11379 9404 11652 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 5307 9336 5764 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 6052 9336 7757 9364
rect 6052 9324 6058 9336
rect 7745 9333 7757 9336
rect 7791 9364 7803 9367
rect 8386 9364 8392 9376
rect 7791 9336 8392 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8478 9324 8484 9376
rect 8536 9324 8542 9376
rect 9582 9324 9588 9376
rect 9640 9324 9646 9376
rect 9858 9324 9864 9376
rect 9916 9324 9922 9376
rect 12069 9367 12127 9373
rect 12069 9333 12081 9367
rect 12115 9364 12127 9367
rect 12342 9364 12348 9376
rect 12115 9336 12348 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13464 9364 13492 9463
rect 12768 9336 13492 9364
rect 12768 9324 12774 9336
rect 13538 9324 13544 9376
rect 13596 9324 13602 9376
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16114 9364 16120 9376
rect 16071 9336 16120 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 1104 9274 16836 9296
rect 1104 9222 2916 9274
rect 2968 9222 2980 9274
rect 3032 9222 3044 9274
rect 3096 9222 3108 9274
rect 3160 9222 3172 9274
rect 3224 9222 6849 9274
rect 6901 9222 6913 9274
rect 6965 9222 6977 9274
rect 7029 9222 7041 9274
rect 7093 9222 7105 9274
rect 7157 9222 10782 9274
rect 10834 9222 10846 9274
rect 10898 9222 10910 9274
rect 10962 9222 10974 9274
rect 11026 9222 11038 9274
rect 11090 9222 14715 9274
rect 14767 9222 14779 9274
rect 14831 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 16836 9274
rect 1104 9200 16836 9222
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4614 9160 4620 9172
rect 3844 9132 4620 9160
rect 3844 9120 3850 9132
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4706 9120 4712 9172
rect 4764 9120 4770 9172
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 5040 9132 6377 9160
rect 5040 9120 5046 9132
rect 6365 9129 6377 9132
rect 6411 9129 6423 9163
rect 6365 9123 6423 9129
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7926 9120 7932 9172
rect 7984 9120 7990 9172
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10468 9132 10609 9160
rect 10468 9120 10474 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13170 9160 13176 9172
rect 12584 9132 13176 9160
rect 12584 9120 12590 9132
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13538 9120 13544 9172
rect 13596 9120 13602 9172
rect 16114 9160 16120 9172
rect 14936 9132 16120 9160
rect 5810 9092 5816 9104
rect 1780 9064 5816 9092
rect 1780 8965 1808 9064
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5905 9095 5963 9101
rect 5905 9061 5917 9095
rect 5951 9092 5963 9095
rect 6822 9092 6828 9104
rect 5951 9064 6828 9092
rect 5951 9061 5963 9064
rect 5905 9055 5963 9061
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 7374 9092 7380 9104
rect 7024 9064 7380 9092
rect 7024 9033 7052 9064
rect 7374 9052 7380 9064
rect 7432 9092 7438 9104
rect 8662 9092 8668 9104
rect 7432 9064 8668 9092
rect 7432 9052 7438 9064
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 11701 9095 11759 9101
rect 11701 9061 11713 9095
rect 11747 9061 11759 9095
rect 11701 9055 11759 9061
rect 12069 9095 12127 9101
rect 12069 9061 12081 9095
rect 12115 9092 12127 9095
rect 12434 9092 12440 9104
rect 12115 9064 12440 9092
rect 12115 9061 12127 9064
rect 12069 9055 12127 9061
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 5902 8916 5908 8968
rect 5960 8916 5966 8968
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 7190 8956 7196 8968
rect 6328 8928 7196 8956
rect 6328 8916 6334 8928
rect 7190 8916 7196 8928
rect 7248 8956 7254 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7248 8928 7757 8956
rect 7248 8916 7254 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 5350 8888 5356 8900
rect 4939 8860 5356 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 5445 8891 5503 8897
rect 5445 8857 5457 8891
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 5460 8820 5488 8851
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 5920 8888 5948 8916
rect 5644 8860 5948 8888
rect 6181 8891 6239 8897
rect 5644 8820 5672 8860
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 8404 8888 8432 8919
rect 8478 8916 8484 8968
rect 8536 8916 8542 8968
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 6227 8860 8432 8888
rect 8496 8888 8524 8916
rect 8956 8888 8984 8919
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 11514 8916 11520 8968
rect 11572 8916 11578 8968
rect 8496 8860 8984 8888
rect 11716 8888 11744 9055
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12544 9024 12572 9120
rect 12452 8996 12572 9024
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 12452 8965 12480 8996
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 12618 8956 12624 8968
rect 12575 8928 12624 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12796 8959 12854 8965
rect 12796 8925 12808 8959
rect 12842 8956 12854 8959
rect 13556 8956 13584 9120
rect 13909 9095 13967 9101
rect 13909 9061 13921 9095
rect 13955 9061 13967 9095
rect 13909 9055 13967 9061
rect 13924 9024 13952 9055
rect 14550 9024 14556 9036
rect 13924 8996 14556 9024
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 12842 8928 13584 8956
rect 12842 8925 12854 8928
rect 12796 8919 12854 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14936 8965 14964 9132
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16393 9163 16451 9169
rect 16393 9129 16405 9163
rect 16439 9160 16451 9163
rect 16758 9160 16764 9172
rect 16439 9132 16764 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 15286 9052 15292 9104
rect 15344 9052 15350 9104
rect 15470 9052 15476 9104
rect 15528 9052 15534 9104
rect 15488 9024 15516 9052
rect 15841 9027 15899 9033
rect 15841 9024 15853 9027
rect 15488 8996 15853 9024
rect 15841 8993 15853 8996
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 14240 8928 14657 8956
rect 14240 8916 14246 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 15749 8891 15807 8897
rect 11716 8860 14044 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 14016 8832 14044 8860
rect 15749 8857 15761 8891
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 5460 8792 5672 8820
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 5868 8792 9045 8820
rect 5868 8780 5874 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 9033 8783 9091 8789
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 13814 8820 13820 8832
rect 10744 8792 13820 8820
rect 10744 8780 10750 8792
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 13998 8780 14004 8832
rect 14056 8780 14062 8832
rect 14090 8780 14096 8832
rect 14148 8780 14154 8832
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15562 8820 15568 8832
rect 15151 8792 15568 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 15764 8820 15792 8851
rect 16114 8848 16120 8900
rect 16172 8848 16178 8900
rect 16206 8820 16212 8832
rect 15764 8792 16212 8820
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 1104 8730 16995 8752
rect 1104 8678 4882 8730
rect 4934 8678 4946 8730
rect 4998 8678 5010 8730
rect 5062 8678 5074 8730
rect 5126 8678 5138 8730
rect 5190 8678 8815 8730
rect 8867 8678 8879 8730
rect 8931 8678 8943 8730
rect 8995 8678 9007 8730
rect 9059 8678 9071 8730
rect 9123 8678 12748 8730
rect 12800 8678 12812 8730
rect 12864 8678 12876 8730
rect 12928 8678 12940 8730
rect 12992 8678 13004 8730
rect 13056 8678 16681 8730
rect 16733 8678 16745 8730
rect 16797 8678 16809 8730
rect 16861 8678 16873 8730
rect 16925 8678 16937 8730
rect 16989 8678 16995 8730
rect 1104 8656 16995 8678
rect 1762 8576 1768 8628
rect 1820 8576 1826 8628
rect 2774 8576 2780 8628
rect 2832 8576 2838 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8616 5963 8619
rect 6086 8616 6092 8628
rect 5951 8588 6092 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6227 8588 8432 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2792 8480 2820 8576
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 2792 8452 3709 8480
rect 1857 8443 1915 8449
rect 3697 8449 3709 8452
rect 3743 8480 3755 8483
rect 3786 8480 3792 8492
rect 3743 8452 3792 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 1872 8344 1900 8443
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4172 8480 4200 8576
rect 5736 8489 5764 8576
rect 6270 8548 6276 8560
rect 6012 8520 6276 8548
rect 6012 8489 6040 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 8404 8548 8432 8588
rect 8478 8576 8484 8628
rect 8536 8576 8542 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8665 8619 8723 8625
rect 8665 8616 8677 8619
rect 8628 8588 8677 8616
rect 8628 8576 8634 8588
rect 8665 8585 8677 8588
rect 8711 8585 8723 8619
rect 8665 8579 8723 8585
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 9732 8588 9781 8616
rect 9732 8576 9738 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 9769 8579 9827 8585
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 9916 8588 10517 8616
rect 9916 8576 9922 8588
rect 10505 8585 10517 8588
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 6880 8520 8064 8548
rect 8404 8520 9076 8548
rect 6880 8508 6886 8520
rect 8036 8489 8064 8520
rect 9048 8489 9076 8520
rect 9692 8520 10456 8548
rect 4111 8452 4200 8480
rect 5721 8483 5779 8489
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 7285 8483 7343 8489
rect 6411 8452 6776 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6748 8424 6776 8452
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 9033 8483 9091 8489
rect 8803 8452 8984 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 4246 8372 4252 8424
rect 4304 8372 4310 8424
rect 4798 8372 4804 8424
rect 4856 8372 4862 8424
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 3973 8347 4031 8353
rect 1872 8316 3944 8344
rect 3510 8236 3516 8288
rect 3568 8236 3574 8288
rect 3916 8276 3944 8316
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4154 8344 4160 8356
rect 4019 8316 4160 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4709 8347 4767 8353
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 5169 8347 5227 8353
rect 5169 8344 5181 8347
rect 4755 8316 5181 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 5169 8313 5181 8316
rect 5215 8344 5227 8347
rect 5534 8344 5540 8356
rect 5215 8316 5540 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6564 8344 6592 8375
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7300 8412 7328 8443
rect 7147 8384 7181 8412
rect 7300 8384 7604 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 5868 8316 6592 8344
rect 7009 8347 7067 8353
rect 5868 8304 5874 8316
rect 7009 8313 7021 8347
rect 7055 8344 7067 8347
rect 7116 8344 7144 8375
rect 7374 8344 7380 8356
rect 7055 8316 7380 8344
rect 7055 8313 7067 8316
rect 7009 8307 7067 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7576 8344 7604 8384
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 7708 8384 7849 8412
rect 7708 8372 7714 8384
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 7837 8375 7895 8381
rect 8849 8347 8907 8353
rect 8849 8344 8861 8347
rect 7576 8316 8861 8344
rect 8849 8313 8861 8316
rect 8895 8313 8907 8347
rect 8956 8344 8984 8452
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9324 8412 9352 8443
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 9692 8424 9720 8520
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9824 8452 10057 8480
rect 9824 8440 9830 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 9674 8412 9680 8424
rect 9324 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10226 8412 10232 8424
rect 9907 8384 10232 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10428 8412 10456 8520
rect 10520 8480 10548 8579
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11572 8588 12173 8616
rect 11572 8576 11578 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12308 8588 12817 8616
rect 12308 8576 12314 8588
rect 12805 8585 12817 8588
rect 12851 8585 12863 8619
rect 13262 8616 13268 8628
rect 12805 8579 12863 8585
rect 13096 8588 13268 8616
rect 10704 8520 11836 8548
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10520 8452 10609 8480
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10704 8412 10732 8520
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11808 8489 11836 8520
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 13096 8557 13124 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13906 8616 13912 8628
rect 13740 8588 13912 8616
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 12492 8520 13093 8548
rect 12492 8508 12498 8520
rect 13081 8517 13093 8520
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 13173 8551 13231 8557
rect 13173 8517 13185 8551
rect 13219 8548 13231 8551
rect 13538 8548 13544 8560
rect 13219 8520 13544 8548
rect 13219 8517 13231 8520
rect 13173 8511 13231 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 13740 8557 13768 8588
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 15194 8576 15200 8628
rect 15252 8576 15258 8628
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 15528 8588 15945 8616
rect 15528 8576 15534 8588
rect 15933 8585 15945 8588
rect 15979 8585 15991 8619
rect 15933 8579 15991 8585
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 16298 8616 16304 8628
rect 16255 8588 16304 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 16390 8576 16396 8628
rect 16448 8576 16454 8628
rect 13725 8551 13783 8557
rect 13725 8517 13737 8551
rect 13771 8517 13783 8551
rect 13725 8511 13783 8517
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13872 8520 16344 8548
rect 13872 8508 13878 8520
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 10428 8384 10732 8412
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 10827 8384 11621 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 9493 8347 9551 8353
rect 8956 8316 9444 8344
rect 8849 8307 8907 8313
rect 9416 8288 9444 8316
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 11330 8344 11336 8356
rect 9539 8316 11336 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12360 8344 12388 8443
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12584 8452 12633 8480
rect 12584 8440 12590 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12894 8480 12900 8492
rect 12621 8443 12679 8449
rect 12728 8452 12900 8480
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 12728 8412 12756 8452
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13998 8440 14004 8492
rect 14056 8440 14062 8492
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14608 8452 14657 8480
rect 14608 8440 14614 8452
rect 14645 8449 14657 8452
rect 14691 8480 14703 8483
rect 15746 8480 15752 8492
rect 14691 8452 15752 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 16316 8489 16344 8520
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 12492 8384 12756 8412
rect 13817 8415 13875 8421
rect 12492 8372 12498 8384
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 12360 8316 13124 8344
rect 13096 8288 13124 8316
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 13832 8344 13860 8375
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15470 8372 15476 8424
rect 15528 8372 15534 8424
rect 16040 8412 16068 8443
rect 16482 8412 16488 8424
rect 16040 8384 16488 8412
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 13228 8316 13860 8344
rect 13228 8304 13234 8316
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16390 8344 16396 8356
rect 16172 8316 16396 8344
rect 16172 8304 16178 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 5718 8276 5724 8288
rect 3916 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 7650 8236 7656 8288
rect 7708 8236 7714 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 11146 8236 11152 8288
rect 11204 8236 11210 8288
rect 11882 8236 11888 8288
rect 11940 8236 11946 8288
rect 12434 8236 12440 8288
rect 12492 8236 12498 8288
rect 13078 8236 13084 8288
rect 13136 8236 13142 8288
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 14274 8276 14280 8288
rect 13412 8248 14280 8276
rect 13412 8236 13418 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 1104 8186 16836 8208
rect 1104 8134 2916 8186
rect 2968 8134 2980 8186
rect 3032 8134 3044 8186
rect 3096 8134 3108 8186
rect 3160 8134 3172 8186
rect 3224 8134 6849 8186
rect 6901 8134 6913 8186
rect 6965 8134 6977 8186
rect 7029 8134 7041 8186
rect 7093 8134 7105 8186
rect 7157 8134 10782 8186
rect 10834 8134 10846 8186
rect 10898 8134 10910 8186
rect 10962 8134 10974 8186
rect 11026 8134 11038 8186
rect 11090 8134 14715 8186
rect 14767 8134 14779 8186
rect 14831 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 16836 8186
rect 1104 8112 16836 8134
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 4246 8072 4252 8084
rect 3651 8044 4252 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4982 8072 4988 8084
rect 4356 8044 4988 8072
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 4356 8004 4384 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5169 8075 5227 8081
rect 5169 8041 5181 8075
rect 5215 8072 5227 8075
rect 5258 8072 5264 8084
rect 5215 8044 5264 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 6454 8072 6460 8084
rect 5767 8044 6460 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7282 8072 7288 8084
rect 7147 8044 7288 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 11790 8072 11796 8084
rect 7760 8044 9444 8072
rect 4111 7976 4384 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 7760 7936 7788 8044
rect 9416 8016 9444 8044
rect 10428 8044 11796 8072
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 8680 7976 9045 8004
rect 2148 7908 7788 7936
rect 7929 7939 7987 7945
rect 2148 7877 2176 7908
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 7975 7908 8309 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8297 7905 8309 7908
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 8680 7880 8708 7976
rect 9033 7973 9045 7976
rect 9079 7973 9091 8007
rect 9033 7967 9091 7973
rect 9398 7964 9404 8016
rect 9456 7964 9462 8016
rect 10428 7945 10456 8044
rect 11790 8032 11796 8044
rect 11848 8072 11854 8084
rect 12618 8072 12624 8084
rect 11848 8044 12624 8072
rect 11848 8032 11854 8044
rect 12618 8032 12624 8044
rect 12676 8072 12682 8084
rect 12676 8044 12848 8072
rect 12676 8032 12682 8044
rect 12820 8004 12848 8044
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 14090 8072 14096 8084
rect 13044 8044 14096 8072
rect 13044 8032 13050 8044
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14458 8032 14464 8084
rect 14516 8032 14522 8084
rect 13817 8007 13875 8013
rect 12820 7976 13308 8004
rect 12820 7945 12848 7976
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7905 10471 7939
rect 10413 7899 10471 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7905 12863 7939
rect 13280 7936 13308 7976
rect 13817 7973 13829 8007
rect 13863 8004 13875 8007
rect 13906 8004 13912 8016
rect 13863 7976 13912 8004
rect 13863 7973 13875 7976
rect 13817 7967 13875 7973
rect 13906 7964 13912 7976
rect 13964 7964 13970 8016
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13280 7908 14841 7936
rect 12805 7899 12863 7905
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3510 7868 3516 7880
rect 3467 7840 3516 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3844 7840 3985 7868
rect 3844 7828 3850 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4212 7840 4261 7868
rect 4212 7828 4218 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4614 7868 4620 7880
rect 4571 7840 4620 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1397 7803 1455 7809
rect 1397 7800 1409 7803
rect 992 7772 1409 7800
rect 992 7760 998 7772
rect 1397 7769 1409 7772
rect 1443 7769 1455 7803
rect 1397 7763 1455 7769
rect 1765 7803 1823 7809
rect 1765 7769 1777 7803
rect 1811 7800 1823 7803
rect 1811 7772 1992 7800
rect 1811 7769 1823 7772
rect 1765 7763 1823 7769
rect 1964 7741 1992 7772
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7701 2007 7735
rect 1949 7695 2007 7701
rect 3326 7692 3332 7744
rect 3384 7692 3390 7744
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4724 7732 4752 7831
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 5718 7760 5724 7812
rect 5776 7760 5782 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7190 7800 7196 7812
rect 7055 7772 7196 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7300 7800 7328 7828
rect 8220 7800 8248 7831
rect 8662 7828 8668 7880
rect 8720 7828 8726 7880
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 10168 7803 10226 7809
rect 7300 7772 8248 7800
rect 8312 7772 9674 7800
rect 4479 7704 4752 7732
rect 5736 7732 5764 7760
rect 8312 7732 8340 7772
rect 5736 7704 8340 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 8570 7692 8576 7744
rect 8628 7692 8634 7744
rect 9646 7732 9674 7772
rect 10168 7769 10180 7803
rect 10214 7800 10226 7803
rect 10318 7800 10324 7812
rect 10214 7772 10324 7800
rect 10214 7769 10226 7772
rect 10168 7763 10226 7769
rect 10318 7760 10324 7772
rect 10376 7760 10382 7812
rect 10502 7760 10508 7812
rect 10560 7760 10566 7812
rect 11057 7803 11115 7809
rect 11057 7769 11069 7803
rect 11103 7769 11115 7803
rect 11057 7763 11115 7769
rect 10520 7732 10548 7760
rect 9646 7704 10548 7732
rect 11072 7732 11100 7763
rect 11146 7760 11152 7812
rect 11204 7760 11210 7812
rect 11882 7800 11888 7812
rect 11256 7772 11888 7800
rect 11256 7732 11284 7772
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 12560 7803 12618 7809
rect 12560 7769 12572 7803
rect 12606 7800 12618 7803
rect 12986 7800 12992 7812
rect 12606 7772 12992 7800
rect 12606 7769 12618 7772
rect 12560 7763 12618 7769
rect 12986 7760 12992 7772
rect 13044 7760 13050 7812
rect 13262 7760 13268 7812
rect 13320 7760 13326 7812
rect 13354 7760 13360 7812
rect 13412 7760 13418 7812
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14108 7800 14136 7831
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 15096 7871 15154 7877
rect 15096 7837 15108 7871
rect 15142 7868 15154 7871
rect 17218 7868 17224 7880
rect 15142 7840 17224 7868
rect 15142 7837 15154 7840
rect 15096 7831 15154 7837
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 13780 7772 14136 7800
rect 13780 7760 13786 7772
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 17126 7800 17132 7812
rect 15620 7772 17132 7800
rect 15620 7760 15626 7772
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 11072 7704 11284 7732
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 13081 7735 13139 7741
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13998 7732 14004 7744
rect 13127 7704 14004 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 16209 7735 16267 7741
rect 16209 7732 16221 7735
rect 15436 7704 16221 7732
rect 15436 7692 15442 7704
rect 16209 7701 16221 7704
rect 16255 7701 16267 7735
rect 16209 7695 16267 7701
rect 1104 7642 16995 7664
rect 1104 7590 4882 7642
rect 4934 7590 4946 7642
rect 4998 7590 5010 7642
rect 5062 7590 5074 7642
rect 5126 7590 5138 7642
rect 5190 7590 8815 7642
rect 8867 7590 8879 7642
rect 8931 7590 8943 7642
rect 8995 7590 9007 7642
rect 9059 7590 9071 7642
rect 9123 7590 12748 7642
rect 12800 7590 12812 7642
rect 12864 7590 12876 7642
rect 12928 7590 12940 7642
rect 12992 7590 13004 7642
rect 13056 7590 16681 7642
rect 16733 7590 16745 7642
rect 16797 7590 16809 7642
rect 16861 7590 16873 7642
rect 16925 7590 16937 7642
rect 16989 7590 16995 7642
rect 1104 7568 16995 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3142 7528 3148 7540
rect 3099 7500 3148 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 3326 7488 3332 7540
rect 3384 7488 3390 7540
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3835 7500 3893 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 3881 7497 3893 7500
rect 3927 7528 3939 7531
rect 4798 7528 4804 7540
rect 3927 7500 4804 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5810 7528 5816 7540
rect 5583 7500 5816 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7497 5963 7531
rect 5905 7491 5963 7497
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 3344 7401 3372 7488
rect 4522 7460 4528 7472
rect 3896 7432 4528 7460
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3329 7395 3387 7401
rect 2915 7364 3096 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 3068 7256 3096 7364
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3234 7324 3240 7336
rect 3191 7296 3240 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 3896 7256 3924 7432
rect 4522 7420 4528 7432
rect 4580 7460 4586 7472
rect 4580 7432 4844 7460
rect 4580 7420 4586 7432
rect 4816 7401 4844 7432
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4387 7364 4721 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4709 7361 4721 7364
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5350 7392 5356 7404
rect 5215 7364 5356 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5500 7364 5733 7392
rect 5500 7352 5506 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5920 7392 5948 7491
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7340 7500 7757 7528
rect 7340 7488 7346 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 8110 7528 8116 7540
rect 7883 7500 8116 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8662 7488 8668 7540
rect 8720 7488 8726 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 10428 7500 11529 7528
rect 6730 7460 6736 7472
rect 6104 7432 6736 7460
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5920 7364 6009 7392
rect 5721 7355 5779 7361
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 6104 7324 6132 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6454 7392 6460 7404
rect 6411 7364 6460 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6638 7401 6644 7404
rect 6632 7355 6644 7401
rect 6638 7352 6644 7355
rect 6696 7352 6702 7404
rect 8680 7392 8708 7488
rect 9300 7463 9358 7469
rect 9300 7429 9312 7463
rect 9346 7460 9358 7463
rect 10428 7460 10456 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13262 7528 13268 7540
rect 13035 7500 13268 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 17034 7528 17040 7540
rect 14231 7500 17040 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 9346 7432 10456 7460
rect 9346 7429 9358 7432
rect 9300 7423 9358 7429
rect 10502 7420 10508 7472
rect 10560 7420 10566 7472
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11146 7460 11152 7472
rect 11103 7432 11152 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11146 7420 11152 7432
rect 11204 7420 11210 7472
rect 12897 7463 12955 7469
rect 12897 7429 12909 7463
rect 12943 7460 12955 7463
rect 13170 7460 13176 7472
rect 12943 7432 13176 7460
rect 12943 7429 12955 7432
rect 12897 7423 12955 7429
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 14108 7460 14136 7488
rect 13924 7432 14136 7460
rect 14645 7463 14703 7469
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8680 7364 8769 7392
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9122 7392 9128 7404
rect 9079 7364 9128 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 13722 7392 13728 7404
rect 13495 7364 13728 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 13924 7401 13952 7432
rect 14645 7429 14657 7463
rect 14691 7460 14703 7463
rect 15381 7463 15439 7469
rect 15381 7460 15393 7463
rect 14691 7432 15393 7460
rect 14691 7429 14703 7432
rect 14645 7423 14703 7429
rect 15381 7429 15393 7432
rect 15427 7460 15439 7463
rect 15654 7460 15660 7472
rect 15427 7432 15660 7460
rect 15427 7429 15439 7432
rect 15381 7423 15439 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14182 7392 14188 7404
rect 14047 7364 14188 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 15804 7364 16313 7392
rect 15804 7352 15810 7364
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 4571 7296 6132 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 8294 7284 8300 7336
rect 8352 7284 8358 7336
rect 8478 7284 8484 7336
rect 8536 7284 8542 7336
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10744 7296 11161 7324
rect 10744 7284 10750 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 11882 7324 11888 7336
rect 11756 7296 11888 7324
rect 11756 7284 11762 7296
rect 11882 7284 11888 7296
rect 11940 7324 11946 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11940 7296 12081 7324
rect 11940 7284 11946 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 14090 7324 14096 7336
rect 13679 7296 14096 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15194 7324 15200 7336
rect 15151 7296 15200 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 15562 7324 15568 7336
rect 15335 7296 15568 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7293 15899 7327
rect 15841 7287 15899 7293
rect 14461 7259 14519 7265
rect 3068 7228 3924 7256
rect 4632 7228 6408 7256
rect 4632 7200 4660 7228
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 4614 7148 4620 7200
rect 4672 7148 4678 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6270 7188 6276 7200
rect 6227 7160 6276 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6380 7188 6408 7228
rect 14461 7225 14473 7259
rect 14507 7256 14519 7259
rect 15856 7256 15884 7287
rect 16022 7284 16028 7336
rect 16080 7284 16086 7336
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 16316 7324 16344 7355
rect 16264 7296 16344 7324
rect 16264 7284 16270 7296
rect 14507 7228 15884 7256
rect 14507 7225 14519 7228
rect 14461 7219 14519 7225
rect 7834 7188 7840 7200
rect 6380 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8386 7148 8392 7200
rect 8444 7188 8450 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8444 7160 8585 7188
rect 8444 7148 8450 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 8573 7151 8631 7157
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 9732 7160 10425 7188
rect 9732 7148 9738 7160
rect 10413 7157 10425 7160
rect 10459 7188 10471 7191
rect 10502 7188 10508 7200
rect 10459 7160 10508 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13596 7160 13829 7188
rect 13596 7148 13602 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 16114 7148 16120 7200
rect 16172 7148 16178 7200
rect 1104 7098 16836 7120
rect 1104 7046 2916 7098
rect 2968 7046 2980 7098
rect 3032 7046 3044 7098
rect 3096 7046 3108 7098
rect 3160 7046 3172 7098
rect 3224 7046 6849 7098
rect 6901 7046 6913 7098
rect 6965 7046 6977 7098
rect 7029 7046 7041 7098
rect 7093 7046 7105 7098
rect 7157 7046 10782 7098
rect 10834 7046 10846 7098
rect 10898 7046 10910 7098
rect 10962 7046 10974 7098
rect 11026 7046 11038 7098
rect 11090 7046 14715 7098
rect 14767 7046 14779 7098
rect 14831 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 16836 7098
rect 1104 7024 16836 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 6457 6987 6515 6993
rect 1820 6956 6408 6984
rect 1820 6944 1826 6956
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 6380 6916 6408 6956
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6638 6984 6644 6996
rect 6503 6956 6644 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 7561 6987 7619 6993
rect 7561 6953 7573 6987
rect 7607 6984 7619 6987
rect 8110 6984 8116 6996
rect 7607 6956 8116 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 10318 6944 10324 6996
rect 10376 6944 10382 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11146 6984 11152 6996
rect 11103 6956 11152 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 11606 6984 11612 6996
rect 11348 6956 11612 6984
rect 8662 6916 8668 6928
rect 5500 6888 5764 6916
rect 6380 6888 8668 6916
rect 5500 6876 5506 6888
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3694 6848 3700 6860
rect 3007 6820 3700 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4672 6820 4997 6848
rect 4672 6808 4678 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 5460 6848 5488 6876
rect 4985 6811 5043 6817
rect 5184 6820 5488 6848
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4246 6780 4252 6792
rect 4203 6752 4252 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4356 6752 4445 6780
rect 3050 6672 3056 6724
rect 3108 6672 3114 6724
rect 3605 6715 3663 6721
rect 3605 6681 3617 6715
rect 3651 6681 3663 6715
rect 3605 6675 3663 6681
rect 3620 6644 3648 6675
rect 4062 6644 4068 6656
rect 3620 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4356 6653 4384 6752
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 5184 6780 5212 6820
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 5736 6848 5764 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 11348 6916 11376 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 13081 6987 13139 6993
rect 13081 6953 13093 6987
rect 13127 6984 13139 6987
rect 13262 6984 13268 6996
rect 13127 6956 13268 6984
rect 13127 6953 13139 6956
rect 13081 6947 13139 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 14918 6984 14924 6996
rect 13412 6956 14924 6984
rect 13412 6944 13418 6956
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 11256 6888 11376 6916
rect 9493 6851 9551 6857
rect 5736 6820 7144 6848
rect 4764 6752 5212 6780
rect 5445 6783 5503 6789
rect 4764 6740 4770 6752
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5460 6712 5488 6743
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5592 6752 6377 6780
rect 5592 6740 5598 6752
rect 6365 6749 6377 6752
rect 6411 6780 6423 6783
rect 6454 6780 6460 6792
rect 6411 6752 6460 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7116 6789 7144 6820
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9582 6848 9588 6860
rect 9539 6820 9588 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9582 6808 9588 6820
rect 9640 6848 9646 6860
rect 9640 6820 10364 6848
rect 9640 6808 9646 6820
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7282 6780 7288 6792
rect 7147 6752 7288 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7984 6752 8033 6780
rect 7984 6740 7990 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 10336 6780 10364 6820
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10873 6851 10931 6857
rect 10873 6848 10885 6851
rect 10560 6820 10885 6848
rect 10560 6808 10566 6820
rect 10873 6817 10885 6820
rect 10919 6817 10931 6851
rect 11256 6848 11284 6888
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 14182 6916 14188 6928
rect 11480 6888 14188 6916
rect 11480 6876 11486 6888
rect 10873 6811 10931 6817
rect 10980 6820 11284 6848
rect 10980 6780 11008 6820
rect 11330 6808 11336 6860
rect 11388 6808 11394 6860
rect 12342 6808 12348 6860
rect 12400 6808 12406 6860
rect 13265 6851 13323 6857
rect 13265 6817 13277 6851
rect 13311 6848 13323 6851
rect 13538 6848 13544 6860
rect 13311 6820 13544 6848
rect 13311 6817 13323 6820
rect 13265 6811 13323 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13688 6820 13829 6848
rect 13688 6808 13694 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 9447 6752 9812 6780
rect 10336 6752 11008 6780
rect 11241 6783 11299 6789
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 4632 6684 5488 6712
rect 4632 6653 4660 6684
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 7892 6684 8677 6712
rect 7892 6672 7898 6684
rect 8665 6681 8677 6684
rect 8711 6681 8723 6715
rect 8665 6675 8723 6681
rect 9784 6656 9812 6752
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11348 6780 11376 6808
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11287 6752 11376 6780
rect 11440 6752 11621 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11146 6672 11152 6724
rect 11204 6712 11210 6724
rect 11440 6712 11468 6752
rect 11609 6749 11621 6752
rect 11655 6780 11667 6783
rect 11882 6780 11888 6792
rect 11655 6752 11888 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12360 6780 12388 6808
rect 12299 6752 12388 6780
rect 12529 6783 12587 6789
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 11204 6684 11468 6712
rect 11204 6672 11210 6684
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 11977 6715 12035 6721
rect 11977 6712 11989 6715
rect 11572 6684 11989 6712
rect 11572 6672 11578 6684
rect 11977 6681 11989 6684
rect 12023 6681 12035 6715
rect 11977 6675 12035 6681
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12544 6712 12572 6743
rect 13446 6740 13452 6792
rect 13504 6740 13510 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 13924 6789 13952 6888
rect 14182 6876 14188 6888
rect 14240 6876 14246 6928
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14792 6888 14964 6916
rect 14792 6876 14798 6888
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 14826 6848 14832 6860
rect 14424 6820 14832 6848
rect 14424 6808 14430 6820
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 14936 6848 14964 6888
rect 15010 6876 15016 6928
rect 15068 6916 15074 6928
rect 15378 6916 15384 6928
rect 15068 6888 15384 6916
rect 15068 6876 15074 6888
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 14936 6820 15761 6848
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 15749 6811 15807 6817
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14056 6752 14565 6780
rect 14056 6740 14062 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 13630 6712 13636 6724
rect 12124 6684 13636 6712
rect 12124 6672 12130 6684
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6613 4399 6647
rect 4341 6607 4399 6613
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 4893 6647 4951 6653
rect 4893 6644 4905 6647
rect 4856 6616 4905 6644
rect 4856 6604 4862 6616
rect 4893 6613 4905 6616
rect 4939 6613 4951 6647
rect 4893 6607 4951 6613
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 5902 6644 5908 6656
rect 5767 6616 5908 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11112 6616 11345 6644
rect 11112 6604 11118 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 12158 6644 12164 6656
rect 11839 6616 12164 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12526 6644 12532 6656
rect 12483 6616 12532 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12676 6616 12725 6644
rect 12676 6604 12682 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 13740 6644 13768 6740
rect 14090 6672 14096 6724
rect 14148 6712 14154 6724
rect 15010 6712 15016 6724
rect 14148 6684 15016 6712
rect 14148 6672 14154 6684
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15378 6672 15384 6724
rect 15436 6672 15442 6724
rect 15473 6715 15531 6721
rect 15473 6681 15485 6715
rect 15519 6712 15531 6715
rect 15519 6684 15608 6712
rect 15519 6681 15531 6684
rect 15473 6675 15531 6681
rect 15580 6656 15608 6684
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 13740 6616 14381 6644
rect 12713 6607 12771 6613
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 15562 6604 15568 6656
rect 15620 6604 15626 6656
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 15712 6616 16405 6644
rect 15712 6604 15718 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 1104 6554 16995 6576
rect 1104 6502 4882 6554
rect 4934 6502 4946 6554
rect 4998 6502 5010 6554
rect 5062 6502 5074 6554
rect 5126 6502 5138 6554
rect 5190 6502 8815 6554
rect 8867 6502 8879 6554
rect 8931 6502 8943 6554
rect 8995 6502 9007 6554
rect 9059 6502 9071 6554
rect 9123 6502 12748 6554
rect 12800 6502 12812 6554
rect 12864 6502 12876 6554
rect 12928 6502 12940 6554
rect 12992 6502 13004 6554
rect 13056 6502 16681 6554
rect 16733 6502 16745 6554
rect 16797 6502 16809 6554
rect 16861 6502 16873 6554
rect 16925 6502 16937 6554
rect 16989 6502 16995 6554
rect 1104 6480 16995 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 3108 6412 3249 6440
rect 3108 6400 3114 6412
rect 3237 6409 3249 6412
rect 3283 6409 3295 6443
rect 3237 6403 3295 6409
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4672 6412 4721 6440
rect 4672 6400 4678 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 7009 6443 7067 6449
rect 4856 6412 6776 6440
rect 4856 6400 4862 6412
rect 1765 6375 1823 6381
rect 1765 6341 1777 6375
rect 1811 6372 1823 6375
rect 5074 6372 5080 6384
rect 1811 6344 5080 6372
rect 1811 6341 1823 6344
rect 1765 6335 1823 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 3326 6264 3332 6316
rect 3384 6264 3390 6316
rect 5902 6264 5908 6316
rect 5960 6313 5966 6316
rect 5960 6304 5972 6313
rect 5960 6276 6005 6304
rect 5960 6267 5972 6276
rect 5960 6264 5966 6267
rect 6178 6264 6184 6316
rect 6236 6264 6242 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6328 6276 6561 6304
rect 6328 6264 6334 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6748 6304 6776 6412
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7374 6440 7380 6452
rect 7055 6412 7380 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7742 6440 7748 6452
rect 7515 6412 7748 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 7834 6400 7840 6452
rect 7892 6400 7898 6452
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10980 6412 11468 6440
rect 8404 6372 8432 6400
rect 10980 6372 11008 6412
rect 7576 6344 8432 6372
rect 8680 6344 11008 6372
rect 7576 6313 7604 6344
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 6748 6276 7297 6304
rect 6549 6267 6607 6273
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8343 6276 8432 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4430 6236 4436 6248
rect 4295 6208 4436 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 6362 6196 6368 6248
rect 6420 6196 6426 6248
rect 8404 6236 8432 6276
rect 8478 6264 8484 6316
rect 8536 6264 8542 6316
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8588 6236 8616 6264
rect 6472 6208 8340 6236
rect 8404 6208 8616 6236
rect 4080 6168 4108 6196
rect 4080 6140 4936 6168
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 992 6072 1501 6100
rect 992 6060 998 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1489 6063 1547 6069
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4764 6072 4813 6100
rect 4764 6060 4770 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4908 6100 4936 6140
rect 6472 6100 6500 6208
rect 7745 6171 7803 6177
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 8202 6168 8208 6180
rect 7791 6140 8208 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 8312 6168 8340 6208
rect 8680 6168 8708 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11440 6372 11468 6412
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 14826 6440 14832 6452
rect 11664 6412 14832 6440
rect 11664 6400 11670 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15470 6440 15476 6452
rect 15427 6412 15476 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 15657 6443 15715 6449
rect 15657 6409 15669 6443
rect 15703 6440 15715 6443
rect 15838 6440 15844 6452
rect 15703 6412 15844 6440
rect 15703 6409 15715 6412
rect 15657 6403 15715 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16574 6400 16580 6452
rect 16632 6400 16638 6452
rect 12437 6375 12495 6381
rect 12437 6372 12449 6375
rect 11112 6344 11284 6372
rect 11440 6344 12449 6372
rect 11112 6332 11118 6344
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9214 6304 9220 6316
rect 9171 6276 9220 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 8312 6140 8708 6168
rect 4908 6072 6500 6100
rect 4801 6063 4859 6069
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8720 6072 8861 6100
rect 8720 6060 8726 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 9048 6100 9076 6267
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9392 6307 9450 6313
rect 9392 6273 9404 6307
rect 9438 6304 9450 6307
rect 9858 6304 9864 6316
rect 9438 6276 9864 6304
rect 9438 6273 9450 6276
rect 9392 6267 9450 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 11256 6313 11284 6344
rect 12437 6341 12449 6344
rect 12483 6341 12495 6375
rect 12437 6335 12495 6341
rect 12986 6332 12992 6384
rect 13044 6332 13050 6384
rect 14274 6332 14280 6384
rect 14332 6332 14338 6384
rect 14366 6332 14372 6384
rect 14424 6332 14430 6384
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 14921 6375 14979 6381
rect 14921 6372 14933 6375
rect 14700 6344 14933 6372
rect 14700 6332 14706 6344
rect 14921 6341 14933 6344
rect 14967 6341 14979 6375
rect 16592 6372 16620 6400
rect 14921 6335 14979 6341
rect 15672 6344 16620 6372
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11422 6236 11428 6248
rect 11103 6208 11428 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 11974 6196 11980 6248
rect 12032 6196 12038 6248
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 13081 6239 13139 6245
rect 12207 6208 12434 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11296 6140 11529 6168
rect 11296 6128 11302 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 12406 6168 12434 6208
rect 13081 6205 13093 6239
rect 13127 6236 13139 6239
rect 13998 6236 14004 6248
rect 13127 6208 14004 6236
rect 13127 6205 13139 6208
rect 13081 6199 13139 6205
rect 12894 6168 12900 6180
rect 12406 6140 12900 6168
rect 11517 6131 11575 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 9766 6100 9772 6112
rect 9048 6072 9772 6100
rect 8849 6063 8907 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 10100 6072 10517 6100
rect 10100 6060 10106 6072
rect 10505 6069 10517 6072
rect 10551 6100 10563 6103
rect 11146 6100 11152 6112
rect 10551 6072 11152 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 13096 6100 13124 6199
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14292 6236 14320 6332
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 15497 6311 15555 6317
rect 15497 6277 15509 6311
rect 15543 6308 15555 6311
rect 15672 6308 15700 6344
rect 17034 6332 17040 6384
rect 17092 6332 17098 6384
rect 15543 6280 15700 6308
rect 15543 6277 15555 6280
rect 15497 6271 15555 6277
rect 14366 6236 14372 6248
rect 14292 6208 14372 6236
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 14608 6208 15025 6236
rect 14608 6196 14614 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 15212 6236 15240 6267
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15804 6276 15945 6304
rect 15804 6264 15810 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17052 6304 17080 6332
rect 16347 6276 17080 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16132 6236 16160 6264
rect 15212 6208 16160 6236
rect 15013 6199 15071 6205
rect 16206 6196 16212 6248
rect 16264 6236 16270 6248
rect 16574 6236 16580 6248
rect 16264 6208 16580 6236
rect 16264 6196 16270 6208
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 13449 6171 13507 6177
rect 13449 6137 13461 6171
rect 13495 6168 13507 6171
rect 13814 6168 13820 6180
rect 13495 6140 13820 6168
rect 13495 6137 13507 6140
rect 13449 6131 13507 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 15749 6171 15807 6177
rect 15749 6168 15761 6171
rect 14292 6140 15761 6168
rect 11940 6072 13124 6100
rect 11940 6060 11946 6072
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14292 6100 14320 6140
rect 15749 6137 15761 6140
rect 15795 6137 15807 6171
rect 15749 6131 15807 6137
rect 13780 6072 14320 6100
rect 13780 6060 13786 6072
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 14976 6072 16129 6100
rect 14976 6060 14982 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16117 6063 16175 6069
rect 1104 6010 16836 6032
rect 1104 5958 2916 6010
rect 2968 5958 2980 6010
rect 3032 5958 3044 6010
rect 3096 5958 3108 6010
rect 3160 5958 3172 6010
rect 3224 5958 6849 6010
rect 6901 5958 6913 6010
rect 6965 5958 6977 6010
rect 7029 5958 7041 6010
rect 7093 5958 7105 6010
rect 7157 5958 10782 6010
rect 10834 5958 10846 6010
rect 10898 5958 10910 6010
rect 10962 5958 10974 6010
rect 11026 5958 11038 6010
rect 11090 5958 14715 6010
rect 14767 5958 14779 6010
rect 14831 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 16836 6010
rect 1104 5936 16836 5958
rect 2148 5868 5028 5896
rect 2148 5701 2176 5868
rect 5000 5760 5028 5868
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5534 5896 5540 5908
rect 5215 5868 5540 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 7193 5899 7251 5905
rect 7193 5865 7205 5899
rect 7239 5896 7251 5899
rect 8294 5896 8300 5908
rect 7239 5868 8300 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8404 5868 10548 5896
rect 5092 5828 5120 5856
rect 7469 5831 7527 5837
rect 7469 5828 7481 5831
rect 5092 5800 7481 5828
rect 7469 5797 7481 5800
rect 7515 5797 7527 5831
rect 8404 5828 8432 5868
rect 7469 5791 7527 5797
rect 8312 5800 8432 5828
rect 5718 5760 5724 5772
rect 5000 5732 5724 5760
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 7190 5760 7196 5772
rect 7024 5732 7196 5760
rect 7024 5701 7052 5732
rect 7190 5720 7196 5732
rect 7248 5760 7254 5772
rect 7834 5760 7840 5772
rect 7248 5732 7840 5760
rect 7248 5720 7254 5732
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 8312 5769 8340 5800
rect 8938 5788 8944 5840
rect 8996 5788 9002 5840
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 9306 5828 9312 5840
rect 9180 5800 9312 5828
rect 9180 5788 9186 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 9401 5831 9459 5837
rect 9401 5797 9413 5831
rect 9447 5828 9459 5831
rect 10318 5828 10324 5840
rect 9447 5800 10324 5828
rect 9447 5797 9459 5800
rect 9401 5791 9459 5797
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 8297 5763 8355 5769
rect 8297 5760 8309 5763
rect 8076 5732 8309 5760
rect 8076 5720 8082 5732
rect 8297 5729 8309 5732
rect 8343 5729 8355 5763
rect 8297 5723 8355 5729
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 10520 5760 10548 5868
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 11606 5896 11612 5908
rect 10652 5868 11612 5896
rect 10652 5856 10658 5868
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11848 5868 11897 5896
rect 11848 5856 11854 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 11900 5828 11928 5859
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 12032 5868 12265 5896
rect 12032 5856 12038 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 12986 5896 12992 5908
rect 12759 5868 12992 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 13320 5868 13461 5896
rect 13320 5856 13326 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14737 5899 14795 5905
rect 13872 5868 14688 5896
rect 13872 5856 13878 5868
rect 12526 5828 12532 5840
rect 11900 5800 12532 5828
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 14660 5828 14688 5868
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15286 5896 15292 5908
rect 14783 5868 15292 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 14660 5800 15056 5828
rect 12066 5760 12072 5772
rect 8720 5732 10456 5760
rect 10520 5732 12072 5760
rect 8720 5720 8726 5732
rect 10428 5704 10456 5732
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12216 5732 12480 5760
rect 12216 5720 12222 5732
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7282 5692 7288 5704
rect 7147 5664 7288 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5624 1823 5627
rect 2041 5627 2099 5633
rect 2041 5624 2053 5627
rect 1811 5596 2053 5624
rect 1811 5593 1823 5596
rect 1765 5587 1823 5593
rect 2041 5593 2053 5596
rect 2087 5593 2099 5627
rect 2041 5587 2099 5593
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 3804 5556 3832 5655
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 8202 5692 8208 5704
rect 7699 5664 8208 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8404 5664 8493 5692
rect 4056 5627 4114 5633
rect 4056 5593 4068 5627
rect 4102 5624 4114 5627
rect 4246 5624 4252 5636
rect 4102 5596 4252 5624
rect 4102 5593 4114 5596
rect 4056 5587 4114 5593
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 6914 5584 6920 5636
rect 6972 5624 6978 5636
rect 6972 5596 7328 5624
rect 6972 5584 6978 5596
rect 4154 5556 4160 5568
rect 3804 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5556 4218 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 4212 5528 5733 5556
rect 4212 5516 4218 5528
rect 5721 5525 5733 5528
rect 5767 5556 5779 5559
rect 6178 5556 6184 5568
rect 5767 5528 6184 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6178 5516 6184 5528
rect 6236 5556 6242 5568
rect 7190 5556 7196 5568
rect 6236 5528 7196 5556
rect 6236 5516 6242 5528
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 7300 5556 7328 5596
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7300 5528 7757 5556
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 8404 5556 8432 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 10042 5692 10048 5704
rect 9263 5664 10048 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10183 5664 10364 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 9490 5584 9496 5636
rect 9548 5584 9554 5636
rect 8478 5556 8484 5568
rect 8404 5528 8484 5556
rect 7745 5519 7803 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 10336 5556 10364 5664
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 12452 5697 12480 5732
rect 12618 5720 12624 5772
rect 12676 5720 12682 5772
rect 12894 5720 12900 5772
rect 12952 5720 12958 5772
rect 15028 5769 15056 5800
rect 15654 5788 15660 5840
rect 15712 5828 15718 5840
rect 16206 5828 16212 5840
rect 15712 5800 16212 5828
rect 15712 5788 15718 5800
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13127 5732 14289 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14277 5723 14335 5729
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 12437 5691 12495 5697
rect 12437 5657 12449 5691
rect 12483 5657 12495 5691
rect 12437 5651 12495 5657
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12636 5692 12664 5720
rect 12575 5664 12664 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12912 5624 12940 5720
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 13044 5664 13277 5692
rect 13044 5652 13050 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 13998 5652 14004 5704
rect 14056 5694 14062 5704
rect 14093 5695 14151 5701
rect 14093 5694 14105 5695
rect 14056 5666 14105 5694
rect 14056 5652 14062 5666
rect 14093 5661 14105 5666
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14829 5695 14887 5701
rect 14829 5692 14841 5695
rect 14516 5664 14841 5692
rect 14516 5652 14522 5664
rect 14829 5661 14841 5664
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 15488 5664 15577 5692
rect 13814 5624 13820 5636
rect 12912 5596 13820 5624
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 15396 5624 15424 5652
rect 15488 5636 15516 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15712 5664 16037 5692
rect 15712 5652 15718 5664
rect 16025 5661 16037 5664
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16209 5695 16267 5701
rect 16209 5692 16221 5695
rect 16172 5664 16221 5692
rect 16172 5652 16178 5664
rect 16209 5661 16221 5664
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 13924 5596 15424 5624
rect 11330 5556 11336 5568
rect 10336 5528 11336 5556
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 13924 5565 13952 5596
rect 15470 5584 15476 5636
rect 15528 5584 15534 5636
rect 16500 5624 16528 5655
rect 16574 5624 16580 5636
rect 16500 5596 16580 5624
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5525 13967 5559
rect 13909 5519 13967 5525
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 14424 5528 16313 5556
rect 14424 5516 14430 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 1104 5466 16995 5488
rect 1104 5414 4882 5466
rect 4934 5414 4946 5466
rect 4998 5414 5010 5466
rect 5062 5414 5074 5466
rect 5126 5414 5138 5466
rect 5190 5414 8815 5466
rect 8867 5414 8879 5466
rect 8931 5414 8943 5466
rect 8995 5414 9007 5466
rect 9059 5414 9071 5466
rect 9123 5414 12748 5466
rect 12800 5414 12812 5466
rect 12864 5414 12876 5466
rect 12928 5414 12940 5466
rect 12992 5414 13004 5466
rect 13056 5414 16681 5466
rect 16733 5414 16745 5466
rect 16797 5414 16809 5466
rect 16861 5414 16873 5466
rect 16925 5414 16937 5466
rect 16989 5414 16995 5466
rect 1104 5392 16995 5414
rect 4246 5312 4252 5364
rect 4304 5312 4310 5364
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 5074 5352 5080 5364
rect 4672 5324 5080 5352
rect 4672 5312 4678 5324
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 8297 5355 8355 5361
rect 5368 5324 6960 5352
rect 5368 5284 5396 5324
rect 6932 5296 6960 5324
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8478 5352 8484 5364
rect 8343 5324 8484 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8680 5324 9674 5352
rect 4080 5256 5396 5284
rect 3901 5219 3959 5225
rect 3901 5185 3913 5219
rect 3947 5216 3959 5219
rect 4080 5216 4108 5256
rect 5442 5244 5448 5296
rect 5500 5244 5506 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 3947 5188 4108 5216
rect 3947 5185 3959 5188
rect 3901 5179 3959 5185
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 4356 5148 4384 5176
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4356 5120 4813 5148
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5000 5080 5028 5179
rect 5074 5176 5080 5228
rect 5132 5176 5138 5228
rect 7009 5219 7067 5225
rect 6564 5188 6960 5216
rect 5092 5148 5120 5176
rect 6564 5160 6592 5188
rect 5353 5151 5411 5157
rect 5353 5148 5365 5151
rect 5092 5120 5365 5148
rect 5353 5117 5365 5120
rect 5399 5117 5411 5151
rect 5353 5111 5411 5117
rect 5460 5120 6040 5148
rect 5460 5080 5488 5120
rect 5000 5052 5488 5080
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 5905 5083 5963 5089
rect 5905 5080 5917 5083
rect 5776 5052 5917 5080
rect 5776 5040 5782 5052
rect 5905 5049 5917 5052
rect 5951 5049 5963 5083
rect 6012 5080 6040 5120
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6932 5148 6960 5188
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 7055 5188 7113 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 7101 5185 7113 5188
rect 7147 5216 7159 5219
rect 7374 5216 7380 5228
rect 7147 5188 7380 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7607 5188 7941 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7929 5185 7941 5188
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 8076 5188 8125 5216
rect 8076 5176 8082 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8680 5216 8708 5324
rect 8938 5244 8944 5296
rect 8996 5244 9002 5296
rect 9646 5284 9674 5324
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 10686 5312 10692 5364
rect 10744 5312 10750 5364
rect 12250 5352 12256 5364
rect 10796 5324 12256 5352
rect 10796 5284 10824 5324
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12345 5355 12403 5361
rect 12345 5321 12357 5355
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 9646 5256 10824 5284
rect 10888 5256 11836 5284
rect 8113 5179 8171 5185
rect 8496 5188 8708 5216
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 6932 5120 7757 5148
rect 6825 5111 6883 5117
rect 7745 5117 7757 5120
rect 7791 5148 7803 5151
rect 8496 5148 8524 5188
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8812 5188 8861 5216
rect 8812 5176 8818 5188
rect 8849 5185 8861 5188
rect 8895 5216 8907 5219
rect 9306 5216 9312 5228
rect 8895 5188 9312 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 10888 5216 10916 5256
rect 10376 5188 10916 5216
rect 11149 5219 11207 5225
rect 10376 5176 10382 5188
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11514 5216 11520 5228
rect 11195 5188 11520 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11808 5216 11836 5256
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12360 5284 12388 5315
rect 13814 5312 13820 5364
rect 13872 5312 13878 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 14608 5324 15853 5352
rect 14608 5312 14614 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 15841 5315 15899 5321
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16356 5324 16405 5352
rect 16356 5312 16362 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 16482 5312 16488 5364
rect 16540 5312 16546 5364
rect 13832 5284 13860 5312
rect 16500 5284 16528 5312
rect 12124 5256 12388 5284
rect 12544 5256 13768 5284
rect 13832 5256 14596 5284
rect 12124 5244 12130 5256
rect 12544 5228 12572 5256
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11808 5188 11989 5216
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12526 5176 12532 5228
rect 12584 5176 12590 5228
rect 13740 5225 13768 5256
rect 14568 5228 14596 5256
rect 15672 5256 16528 5284
rect 13469 5219 13527 5225
rect 13469 5185 13481 5219
rect 13515 5216 13527 5219
rect 13725 5219 13783 5225
rect 13515 5188 13676 5216
rect 13515 5185 13527 5188
rect 13469 5179 13527 5185
rect 7791 5120 8524 5148
rect 8573 5151 8631 5157
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8478 5080 8484 5092
rect 6012 5052 8484 5080
rect 5905 5043 5963 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 8588 5080 8616 5111
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 8720 5120 9413 5148
rect 8720 5108 8726 5120
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9692 5148 9720 5176
rect 10410 5148 10416 5160
rect 9692 5120 10416 5148
rect 9401 5111 9459 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 13648 5148 13676 5188
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13725 5179 13783 5185
rect 13924 5188 14381 5216
rect 13817 5151 13875 5157
rect 13817 5148 13829 5151
rect 11379 5120 12434 5148
rect 13648 5120 13829 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 9122 5080 9128 5092
rect 8588 5052 9128 5080
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 11793 5083 11851 5089
rect 11793 5080 11805 5083
rect 11480 5052 11805 5080
rect 11480 5040 11486 5052
rect 11793 5049 11805 5052
rect 11839 5049 11851 5083
rect 11793 5043 11851 5049
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 4338 5012 4344 5024
rect 2823 4984 4344 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 5012 5227 5015
rect 5534 5012 5540 5024
rect 5215 4984 5540 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8628 4984 8769 5012
rect 8628 4972 8634 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 8846 4972 8852 5024
rect 8904 5012 8910 5024
rect 11238 5012 11244 5024
rect 8904 4984 11244 5012
rect 8904 4972 8910 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 12406 5012 12434 5120
rect 13817 5117 13829 5120
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 13722 5040 13728 5092
rect 13780 5080 13786 5092
rect 13924 5080 13952 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 15470 5216 15476 5228
rect 15120 5188 15476 5216
rect 15120 5148 15148 5188
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 15672 5225 15700 5256
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15804 5188 15945 5216
rect 15804 5176 15810 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16390 5216 16396 5228
rect 16347 5188 16396 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 13780 5052 13952 5080
rect 14108 5120 15148 5148
rect 13780 5040 13786 5052
rect 14108 5012 14136 5120
rect 15194 5108 15200 5160
rect 15252 5108 15258 5160
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15381 5151 15439 5157
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 16114 5148 16120 5160
rect 15427 5120 16120 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 16224 5148 16252 5179
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 16574 5148 16580 5160
rect 16224 5120 16580 5148
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 15304 5080 15332 5108
rect 15304 5052 16160 5080
rect 12406 4984 14136 5012
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14737 5015 14795 5021
rect 14737 5012 14749 5015
rect 14240 4984 14749 5012
rect 14240 4972 14246 4984
rect 14737 4981 14749 4984
rect 14783 4981 14795 5015
rect 14737 4975 14795 4981
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 16132 5021 16160 5052
rect 16117 5015 16175 5021
rect 16117 4981 16129 5015
rect 16163 4981 16175 5015
rect 16117 4975 16175 4981
rect 1104 4922 16836 4944
rect 1104 4870 2916 4922
rect 2968 4870 2980 4922
rect 3032 4870 3044 4922
rect 3096 4870 3108 4922
rect 3160 4870 3172 4922
rect 3224 4870 6849 4922
rect 6901 4870 6913 4922
rect 6965 4870 6977 4922
rect 7029 4870 7041 4922
rect 7093 4870 7105 4922
rect 7157 4870 10782 4922
rect 10834 4870 10846 4922
rect 10898 4870 10910 4922
rect 10962 4870 10974 4922
rect 11026 4870 11038 4922
rect 11090 4870 14715 4922
rect 14767 4870 14779 4922
rect 14831 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 16836 4922
rect 1104 4848 16836 4870
rect 4430 4768 4436 4820
rect 4488 4768 4494 4820
rect 6362 4768 6368 4820
rect 6420 4768 6426 4820
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 8846 4808 8852 4820
rect 8711 4780 8852 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9214 4808 9220 4820
rect 8956 4780 9220 4808
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 5997 4743 6055 4749
rect 5997 4740 6009 4743
rect 5776 4712 6009 4740
rect 5776 4700 5782 4712
rect 5997 4709 6009 4712
rect 6043 4709 6055 4743
rect 5997 4703 6055 4709
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4295 4644 4629 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5307 4644 5457 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5445 4641 5457 4644
rect 5491 4672 5503 4675
rect 6380 4672 6408 4768
rect 5491 4644 6408 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8956 4681 8984 4780
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 10410 4808 10416 4820
rect 10367 4780 10416 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13722 4808 13728 4820
rect 13403 4780 13728 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 15194 4808 15200 4820
rect 14691 4780 15200 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 15105 4743 15163 4749
rect 15105 4740 15117 4743
rect 14240 4712 15117 4740
rect 14240 4700 14246 4712
rect 15105 4709 15117 4712
rect 15151 4709 15163 4743
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 15105 4703 15163 4709
rect 15212 4712 15853 4740
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8076 4644 8953 4672
rect 8076 4632 8082 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 14274 4632 14280 4684
rect 14332 4632 14338 4684
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15212 4672 15240 4712
rect 15841 4709 15853 4712
rect 15887 4709 15899 4743
rect 15841 4703 15899 4709
rect 14700 4644 15240 4672
rect 15473 4675 15531 4681
rect 14700 4632 14706 4644
rect 15473 4641 15485 4675
rect 15519 4672 15531 4675
rect 15519 4644 15792 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 4338 4604 4344 4616
rect 3835 4576 4344 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4338 4564 4344 4576
rect 4396 4604 4402 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4396 4576 4537 4604
rect 4396 4564 4402 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7098 4604 7104 4616
rect 7055 4576 7104 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7098 4564 7104 4576
rect 7156 4604 7162 4616
rect 8036 4604 8064 4632
rect 7156 4576 8064 4604
rect 7156 4564 7162 4576
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8352 4576 8585 4604
rect 8352 4564 8358 4576
rect 8573 4573 8585 4576
rect 8619 4604 8631 4607
rect 11885 4607 11943 4613
rect 8619 4576 8892 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1397 4539 1455 4545
rect 1397 4536 1409 4539
rect 992 4508 1409 4536
rect 992 4496 998 4508
rect 1397 4505 1409 4508
rect 1443 4505 1455 4539
rect 1397 4499 1455 4505
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 5258 4536 5264 4548
rect 1811 4508 5264 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5534 4496 5540 4548
rect 5592 4496 5598 4548
rect 6917 4539 6975 4545
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 7254 4539 7312 4545
rect 7254 4536 7266 4539
rect 6963 4508 7266 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 7254 4505 7266 4508
rect 7300 4505 7312 4539
rect 7254 4499 7312 4505
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4154 4468 4160 4480
rect 4019 4440 4160 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 8389 4471 8447 4477
rect 8389 4437 8401 4471
rect 8435 4468 8447 4471
rect 8662 4468 8668 4480
rect 8435 4440 8668 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 8864 4468 8892 4576
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11931 4576 11989 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 11977 4573 11989 4576
rect 12023 4604 12035 4607
rect 12526 4604 12532 4616
rect 12023 4576 12532 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 13136 4576 13461 4604
rect 13136 4564 13142 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 13538 4564 13544 4616
rect 13596 4564 13602 4616
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 14292 4604 14320 4632
rect 15764 4616 15792 4644
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 16080 4644 16221 4672
rect 16080 4632 16086 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 14231 4576 14320 4604
rect 14384 4576 14473 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 9208 4539 9266 4545
rect 9208 4505 9220 4539
rect 9254 4536 9266 4539
rect 9582 4536 9588 4548
rect 9254 4508 9588 4536
rect 9254 4505 9266 4508
rect 9208 4499 9266 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 11640 4539 11698 4545
rect 11640 4505 11652 4539
rect 11686 4536 11698 4539
rect 11686 4508 12020 4536
rect 11686 4505 11698 4508
rect 11640 4499 11698 4505
rect 9306 4468 9312 4480
rect 8864 4440 9312 4468
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 10505 4471 10563 4477
rect 10505 4437 10517 4471
rect 10551 4468 10563 4471
rect 11422 4468 11428 4480
rect 10551 4440 11428 4468
rect 10551 4437 10563 4440
rect 10505 4431 10563 4437
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 11992 4468 12020 4508
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 12222 4539 12280 4545
rect 12222 4536 12234 4539
rect 12124 4508 12234 4536
rect 12124 4496 12130 4508
rect 12222 4505 12234 4508
rect 12268 4505 12280 4539
rect 13556 4536 13584 4564
rect 12222 4499 12280 4505
rect 12406 4508 13584 4536
rect 12406 4468 12434 4508
rect 11992 4440 12434 4468
rect 13354 4428 13360 4480
rect 13412 4468 13418 4480
rect 13541 4471 13599 4477
rect 13541 4468 13553 4471
rect 13412 4440 13553 4468
rect 13412 4428 13418 4440
rect 13541 4437 13553 4440
rect 13587 4437 13599 4471
rect 13541 4431 13599 4437
rect 13906 4428 13912 4480
rect 13964 4428 13970 4480
rect 14384 4477 14412 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 14737 4607 14795 4613
rect 14737 4604 14749 4607
rect 14608 4576 14749 4604
rect 14608 4564 14614 4576
rect 14737 4573 14749 4576
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 14918 4564 14924 4616
rect 14976 4564 14982 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15657 4607 15715 4613
rect 15657 4604 15669 4607
rect 15436 4576 15669 4604
rect 15436 4564 15442 4576
rect 15657 4573 15669 4576
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 15746 4564 15752 4616
rect 15804 4564 15810 4616
rect 14369 4471 14427 4477
rect 14369 4437 14381 4471
rect 14415 4437 14427 4471
rect 14369 4431 14427 4437
rect 1104 4378 16995 4400
rect 1104 4326 4882 4378
rect 4934 4326 4946 4378
rect 4998 4326 5010 4378
rect 5062 4326 5074 4378
rect 5126 4326 5138 4378
rect 5190 4326 8815 4378
rect 8867 4326 8879 4378
rect 8931 4326 8943 4378
rect 8995 4326 9007 4378
rect 9059 4326 9071 4378
rect 9123 4326 12748 4378
rect 12800 4326 12812 4378
rect 12864 4326 12876 4378
rect 12928 4326 12940 4378
rect 12992 4326 13004 4378
rect 13056 4326 16681 4378
rect 16733 4326 16745 4378
rect 16797 4326 16809 4378
rect 16861 4326 16873 4378
rect 16925 4326 16937 4378
rect 16989 4326 16995 4378
rect 1104 4304 16995 4326
rect 4154 4224 4160 4276
rect 4212 4224 4218 4276
rect 4338 4224 4344 4276
rect 4396 4224 4402 4276
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 4798 4264 4804 4276
rect 4571 4236 4804 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5258 4224 5264 4276
rect 5316 4224 5322 4276
rect 6362 4224 6368 4276
rect 6420 4224 6426 4276
rect 7834 4224 7840 4276
rect 7892 4224 7898 4276
rect 8570 4264 8576 4276
rect 8404 4236 8576 4264
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4196 1823 4199
rect 3786 4196 3792 4208
rect 1811 4168 3792 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 4172 4128 4200 4224
rect 4356 4196 4384 4224
rect 4356 4168 5028 4196
rect 5000 4137 5028 4168
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4172 4100 4353 4128
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5534 4128 5540 4140
rect 5491 4100 5540 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4632 4060 4660 4091
rect 5534 4088 5540 4100
rect 5592 4128 5598 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5592 4100 6009 4128
rect 5592 4088 5598 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6270 4128 6276 4140
rect 6135 4100 6276 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6730 4088 6736 4140
rect 6788 4088 6794 4140
rect 7466 4088 7472 4140
rect 7524 4137 7530 4140
rect 7524 4128 7536 4137
rect 7852 4128 7880 4224
rect 8404 4205 8432 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 12066 4224 12072 4276
rect 12124 4224 12130 4276
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 14274 4264 14280 4276
rect 13188 4236 14280 4264
rect 8389 4199 8447 4205
rect 8389 4165 8401 4199
rect 8435 4165 8447 4199
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 8389 4159 8447 4165
rect 8956 4168 9229 4196
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7524 4100 7569 4128
rect 7852 4100 7941 4128
rect 7524 4091 7536 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 7524 4088 7530 4091
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 4120 4032 4660 4060
rect 5077 4063 5135 4069
rect 4120 4020 4126 4032
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 6748 4060 6776 4088
rect 5123 4032 6776 4060
rect 7745 4063 7803 4069
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 8036 4060 8064 4088
rect 7791 4032 8064 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 8294 4020 8300 4072
rect 8352 4020 8358 4072
rect 8956 4060 8984 4168
rect 9217 4165 9229 4168
rect 9263 4165 9275 4199
rect 9217 4159 9275 4165
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 13096 4196 13124 4224
rect 11480 4168 11836 4196
rect 11480 4156 11486 4168
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 9907 4100 10241 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10229 4097 10241 4100
rect 10275 4128 10287 4131
rect 10778 4128 10784 4140
rect 10275 4100 10784 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11514 4128 11520 4140
rect 11011 4100 11520 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11808 4137 11836 4168
rect 12728 4168 13124 4196
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12158 4128 12164 4140
rect 11839 4100 12164 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12158 4088 12164 4100
rect 12216 4128 12222 4140
rect 12728 4137 12756 4168
rect 12713 4131 12771 4137
rect 12713 4128 12725 4131
rect 12216 4100 12725 4128
rect 12216 4088 12222 4100
rect 12713 4097 12725 4100
rect 12759 4097 12771 4131
rect 13188 4128 13216 4236
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 14369 4267 14427 4273
rect 14369 4233 14381 4267
rect 14415 4264 14427 4267
rect 14918 4264 14924 4276
rect 14415 4236 14924 4264
rect 14415 4233 14427 4236
rect 14369 4227 14427 4233
rect 14918 4224 14924 4236
rect 14976 4224 14982 4276
rect 15470 4224 15476 4276
rect 15528 4224 15534 4276
rect 13464 4168 14412 4196
rect 12713 4091 12771 4097
rect 12912 4100 13216 4128
rect 13265 4131 13323 4137
rect 8772 4032 8984 4060
rect 9125 4063 9183 4069
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 6546 3992 6552 4004
rect 4755 3964 6552 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 8113 3995 8171 4001
rect 8113 3961 8125 3995
rect 8159 3992 8171 3995
rect 8772 3992 8800 4032
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9214 4060 9220 4072
rect 9171 4032 9220 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 9950 4060 9956 4072
rect 9815 4032 9956 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 8159 3964 8800 3992
rect 8849 3995 8907 4001
rect 8159 3961 8171 3964
rect 8113 3955 8171 3961
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 9784 3992 9812 4023
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4060 11207 4063
rect 11238 4060 11244 4072
rect 11195 4032 11244 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11698 4020 11704 4072
rect 11756 4020 11762 4072
rect 12912 4060 12940 4100
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13354 4128 13360 4140
rect 13311 4100 13360 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13464 4137 13492 4168
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13964 4100 14013 4128
rect 13964 4088 13970 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14274 4088 14280 4140
rect 14332 4088 14338 4140
rect 14384 4128 14412 4168
rect 14642 4156 14648 4208
rect 14700 4196 14706 4208
rect 15197 4199 15255 4205
rect 15197 4196 15209 4199
rect 14700 4168 15209 4196
rect 14700 4156 14706 4168
rect 15197 4165 15209 4168
rect 15243 4165 15255 4199
rect 15197 4159 15255 4165
rect 15488 4137 15516 4224
rect 15473 4131 15531 4137
rect 14384 4100 15424 4128
rect 11808 4032 12940 4060
rect 8895 3964 9812 3992
rect 10045 3995 10103 4001
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 11716 3992 11744 4020
rect 10091 3964 11744 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 992 3896 1501 3924
rect 992 3884 998 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 9490 3924 9496 3936
rect 7524 3896 9496 3924
rect 7524 3884 7530 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 10318 3884 10324 3936
rect 10376 3884 10382 3936
rect 10686 3884 10692 3936
rect 10744 3884 10750 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11808 3924 11836 4032
rect 12986 4020 12992 4072
rect 13044 4060 13050 4072
rect 14550 4060 14556 4072
rect 13044 4032 14556 4060
rect 13044 4020 13050 4032
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14700 4032 14749 4060
rect 14700 4020 14706 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 15396 4060 15424 4100
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 15562 4088 15568 4140
rect 15620 4088 15626 4140
rect 16206 4128 16212 4140
rect 15672 4100 16212 4128
rect 15672 4060 15700 4100
rect 16206 4088 16212 4100
rect 16264 4128 16270 4140
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 16264 4100 16405 4128
rect 16264 4088 16270 4100
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 15396 4032 15700 4060
rect 14737 4023 14795 4029
rect 15746 4020 15752 4072
rect 15804 4020 15810 4072
rect 15933 4063 15991 4069
rect 15933 4029 15945 4063
rect 15979 4060 15991 4063
rect 16022 4060 16028 4072
rect 15979 4032 16028 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 11977 3995 12035 4001
rect 11977 3961 11989 3995
rect 12023 3992 12035 3995
rect 13722 3992 13728 4004
rect 12023 3964 13728 3992
rect 12023 3961 12035 3964
rect 11977 3955 12035 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 14274 3952 14280 4004
rect 14332 3952 14338 4004
rect 10836 3896 11836 3924
rect 13081 3927 13139 3933
rect 10836 3884 10842 3896
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13262 3924 13268 3936
rect 13127 3896 13268 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13262 3884 13268 3896
rect 13320 3924 13326 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13320 3896 13553 3924
rect 13320 3884 13326 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 14292 3924 14320 3952
rect 16206 3924 16212 3936
rect 14292 3896 16212 3924
rect 13541 3887 13599 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 1104 3834 16836 3856
rect 1104 3782 2916 3834
rect 2968 3782 2980 3834
rect 3032 3782 3044 3834
rect 3096 3782 3108 3834
rect 3160 3782 3172 3834
rect 3224 3782 6849 3834
rect 6901 3782 6913 3834
rect 6965 3782 6977 3834
rect 7029 3782 7041 3834
rect 7093 3782 7105 3834
rect 7157 3782 10782 3834
rect 10834 3782 10846 3834
rect 10898 3782 10910 3834
rect 10962 3782 10974 3834
rect 11026 3782 11038 3834
rect 11090 3782 14715 3834
rect 14767 3782 14779 3834
rect 14831 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 16836 3834
rect 1104 3760 16836 3782
rect 3786 3680 3792 3732
rect 3844 3680 3850 3732
rect 9582 3680 9588 3732
rect 9640 3680 9646 3732
rect 10318 3680 10324 3732
rect 10376 3680 10382 3732
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 13262 3680 13268 3732
rect 13320 3680 13326 3732
rect 14550 3680 14556 3732
rect 14608 3680 14614 3732
rect 15105 3723 15163 3729
rect 15105 3689 15117 3723
rect 15151 3720 15163 3723
rect 15378 3720 15384 3732
rect 15151 3692 15384 3720
rect 15151 3689 15163 3692
rect 15105 3683 15163 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15654 3680 15660 3732
rect 15712 3680 15718 3732
rect 16114 3680 16120 3732
rect 16172 3680 16178 3732
rect 16298 3680 16304 3732
rect 16356 3680 16362 3732
rect 8021 3655 8079 3661
rect 8021 3621 8033 3655
rect 8067 3652 8079 3655
rect 8294 3652 8300 3664
rect 8067 3624 8300 3652
rect 8067 3621 8079 3624
rect 8021 3615 8079 3621
rect 8294 3612 8300 3624
rect 8352 3652 8358 3664
rect 8481 3655 8539 3661
rect 8481 3652 8493 3655
rect 8352 3624 8493 3652
rect 8352 3612 8358 3624
rect 8481 3621 8493 3624
rect 8527 3621 8539 3655
rect 8481 3615 8539 3621
rect 4062 3584 4068 3596
rect 3988 3556 4068 3584
rect 3988 3525 4016 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7239 3556 7573 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 7561 3547 7619 3553
rect 8036 3556 10241 3584
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 6420 3488 6837 3516
rect 6420 3476 6426 3488
rect 6825 3485 6837 3488
rect 6871 3516 6883 3519
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6871 3488 7113 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 8036 3516 8064 3556
rect 10229 3553 10241 3556
rect 10275 3553 10287 3587
rect 10336 3584 10364 3680
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10336 3556 10425 3584
rect 10229 3547 10287 3553
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 10744 3556 11253 3584
rect 10744 3544 10750 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 12986 3584 12992 3596
rect 11572 3556 12992 3584
rect 11572 3544 11578 3556
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13280 3593 13308 3680
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3652 14335 3655
rect 14323 3624 14412 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 13265 3587 13323 3593
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 14384 3541 14412 3624
rect 14458 3612 14464 3664
rect 14516 3652 14522 3664
rect 14516 3624 15424 3652
rect 14516 3612 14522 3624
rect 15396 3593 15424 3624
rect 15381 3587 15439 3593
rect 14568 3556 15332 3584
rect 14369 3535 14427 3541
rect 7423 3488 8064 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7392 3448 7420 3479
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 6972 3420 7420 3448
rect 6972 3408 6978 3420
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 8312 3448 8340 3479
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8720 3488 8953 3516
rect 8720 3476 8726 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11471 3488 12081 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12158 3476 12164 3528
rect 12216 3476 12222 3528
rect 12360 3488 13032 3516
rect 7524 3420 8340 3448
rect 7524 3408 7530 3420
rect 10410 3408 10416 3460
rect 10468 3448 10474 3460
rect 12360 3448 12388 3488
rect 10468 3420 12388 3448
rect 10468 3408 10474 3420
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13004 3448 13032 3488
rect 13078 3476 13084 3528
rect 13136 3476 13142 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13630 3516 13636 3528
rect 13587 3488 13636 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14369 3501 14381 3535
rect 14415 3501 14427 3535
rect 14568 3528 14596 3556
rect 14369 3495 14427 3501
rect 14093 3479 14151 3485
rect 14108 3448 14136 3479
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 15304 3525 15332 3556
rect 15381 3553 15393 3587
rect 15427 3553 15439 3587
rect 15381 3547 15439 3553
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3516 14703 3519
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14691 3488 15025 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 14660 3448 14688 3479
rect 12492 3420 12756 3448
rect 13004 3420 14688 3448
rect 15028 3448 15056 3479
rect 15580 3448 15608 3479
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15896 3488 16037 3516
rect 15896 3476 15902 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16025 3479 16083 3485
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3516 16543 3519
rect 17126 3516 17132 3528
rect 16531 3488 17132 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 15028 3420 15608 3448
rect 12492 3408 12498 3420
rect 7006 3340 7012 3392
rect 7064 3340 7070 3392
rect 11882 3340 11888 3392
rect 11940 3340 11946 3392
rect 12250 3340 12256 3392
rect 12308 3340 12314 3392
rect 12618 3340 12624 3392
rect 12676 3340 12682 3392
rect 12728 3380 12756 3420
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12728 3352 13369 3380
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 14550 3380 14556 3392
rect 13955 3352 14556 3380
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14826 3340 14832 3392
rect 14884 3340 14890 3392
rect 1104 3290 16995 3312
rect 1104 3238 4882 3290
rect 4934 3238 4946 3290
rect 4998 3238 5010 3290
rect 5062 3238 5074 3290
rect 5126 3238 5138 3290
rect 5190 3238 8815 3290
rect 8867 3238 8879 3290
rect 8931 3238 8943 3290
rect 8995 3238 9007 3290
rect 9059 3238 9071 3290
rect 9123 3238 12748 3290
rect 12800 3238 12812 3290
rect 12864 3238 12876 3290
rect 12928 3238 12940 3290
rect 12992 3238 13004 3290
rect 13056 3238 16681 3290
rect 16733 3238 16745 3290
rect 16797 3238 16809 3290
rect 16861 3238 16873 3290
rect 16925 3238 16937 3290
rect 16989 3238 16995 3290
rect 1104 3216 16995 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3234 3176 3240 3188
rect 3007 3148 3240 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 1964 3108 1992 3139
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7466 3136 7472 3188
rect 7524 3136 7530 3188
rect 7653 3179 7711 3185
rect 7653 3145 7665 3179
rect 7699 3176 7711 3179
rect 8110 3176 8116 3188
rect 7699 3148 8116 3176
rect 7699 3145 7711 3148
rect 7653 3139 7711 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8386 3176 8392 3188
rect 8343 3148 8392 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11514 3176 11520 3188
rect 11011 3148 11520 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11609 3179 11667 3185
rect 11609 3145 11621 3179
rect 11655 3176 11667 3179
rect 11882 3176 11888 3188
rect 11655 3148 11888 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12250 3136 12256 3188
rect 12308 3136 12314 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12894 3176 12900 3188
rect 12676 3148 12900 3176
rect 12676 3136 12682 3148
rect 12894 3136 12900 3148
rect 12952 3176 12958 3188
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 12952 3148 13001 3176
rect 12952 3136 12958 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 12989 3139 13047 3145
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 13136 3148 13185 3176
rect 13136 3136 13142 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 13446 3136 13452 3188
rect 13504 3136 13510 3188
rect 13630 3136 13636 3188
rect 13688 3136 13694 3188
rect 13906 3136 13912 3188
rect 13964 3136 13970 3188
rect 15194 3136 15200 3188
rect 15252 3136 15258 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15344 3148 15669 3176
rect 15344 3136 15350 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 15930 3136 15936 3188
rect 15988 3136 15994 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 17218 3176 17224 3188
rect 16347 3148 17224 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 1811 3080 1992 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2148 2972 2176 3003
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 7024 3040 7052 3136
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 8021 3111 8079 3117
rect 8021 3108 8033 3111
rect 7984 3080 8033 3108
rect 7984 3068 7990 3080
rect 8021 3077 8033 3080
rect 8067 3077 8079 3111
rect 11698 3108 11704 3120
rect 8021 3071 8079 3077
rect 8404 3080 11704 3108
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7024 3012 7297 3040
rect 6825 3003 6883 3009
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 2590 2972 2596 2984
rect 2148 2944 2596 2972
rect 2590 2932 2596 2944
rect 2648 2972 2654 2984
rect 6840 2972 6868 3003
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 8404 3049 8432 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11422 3040 11428 3052
rect 11195 3012 11428 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 2648 2944 6868 2972
rect 2648 2932 2654 2944
rect 8128 2904 8156 3003
rect 11072 2972 11100 3003
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 11900 3040 11928 3136
rect 12268 3049 12296 3136
rect 13648 3108 13676 3136
rect 13280 3080 13676 3108
rect 15212 3108 15240 3136
rect 15212 3080 16528 3108
rect 13280 3049 13308 3080
rect 12253 3043 12311 3049
rect 11900 3012 12204 3040
rect 11606 2972 11612 2984
rect 11072 2944 11612 2972
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 12066 2932 12072 2984
rect 12124 2932 12130 2984
rect 12176 2972 12204 3012
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 13354 3000 13360 3052
rect 13412 3000 13418 3052
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14826 3040 14832 3052
rect 14691 3012 14832 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16206 3040 16212 3052
rect 16071 3012 16212 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16206 3000 16212 3012
rect 16264 3000 16270 3052
rect 16500 3049 16528 3080
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3009 16543 3043
rect 16485 3003 16543 3009
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12176 2944 12357 2972
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 12526 2932 12532 2984
rect 12584 2932 12590 2984
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14507 2944 15025 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 14093 2907 14151 2913
rect 14093 2904 14105 2907
rect 8128 2876 14105 2904
rect 14093 2873 14105 2876
rect 14139 2873 14151 2907
rect 14093 2867 14151 2873
rect 14829 2907 14887 2913
rect 14829 2873 14841 2907
rect 14875 2904 14887 2907
rect 15212 2904 15240 2935
rect 14875 2876 15240 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 992 2808 1501 2836
rect 992 2796 998 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 11330 2796 11336 2848
rect 11388 2796 11394 2848
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 15102 2836 15108 2848
rect 11756 2808 15108 2836
rect 11756 2796 11762 2808
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 1104 2746 16836 2768
rect 1104 2694 2916 2746
rect 2968 2694 2980 2746
rect 3032 2694 3044 2746
rect 3096 2694 3108 2746
rect 3160 2694 3172 2746
rect 3224 2694 6849 2746
rect 6901 2694 6913 2746
rect 6965 2694 6977 2746
rect 7029 2694 7041 2746
rect 7093 2694 7105 2746
rect 7157 2694 10782 2746
rect 10834 2694 10846 2746
rect 10898 2694 10910 2746
rect 10962 2694 10974 2746
rect 11026 2694 11038 2746
rect 11090 2694 14715 2746
rect 14767 2694 14779 2746
rect 14831 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 16836 2746
rect 1104 2672 16836 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2774 2632 2780 2644
rect 2179 2604 2780 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 4062 2592 4068 2644
rect 4120 2592 4126 2644
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7558 2632 7564 2644
rect 7055 2604 7564 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9306 2632 9312 2644
rect 8527 2604 9312 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 11422 2592 11428 2644
rect 11480 2592 11486 2644
rect 11606 2592 11612 2644
rect 11664 2592 11670 2644
rect 11793 2635 11851 2641
rect 11793 2601 11805 2635
rect 11839 2632 11851 2635
rect 12066 2632 12072 2644
rect 11839 2604 12072 2632
rect 11839 2601 11851 2604
rect 11793 2595 11851 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12526 2632 12532 2644
rect 12483 2604 12532 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13354 2632 13360 2644
rect 13219 2604 13360 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 14185 2595 14243 2601
rect 14366 2592 14372 2644
rect 14424 2592 14430 2644
rect 14645 2635 14703 2641
rect 14645 2601 14657 2635
rect 14691 2632 14703 2635
rect 15746 2632 15752 2644
rect 14691 2604 15752 2632
rect 14691 2601 14703 2604
rect 14645 2595 14703 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 16022 2592 16028 2644
rect 16080 2592 16086 2644
rect 2590 2524 2596 2576
rect 2648 2524 2654 2576
rect 11057 2567 11115 2573
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 11440 2564 11468 2592
rect 11103 2536 11468 2564
rect 11624 2564 11652 2592
rect 12161 2567 12219 2573
rect 12161 2564 12173 2567
rect 11624 2536 12173 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 12161 2533 12173 2536
rect 12207 2533 12219 2567
rect 12161 2527 12219 2533
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 14384 2564 14412 2592
rect 13679 2536 14412 2564
rect 14829 2567 14887 2573
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 14829 2533 14841 2567
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6696 2468 9628 2496
rect 6696 2456 6702 2468
rect 9600 2440 9628 2468
rect 10060 2468 12296 2496
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 900 2400 1961 2428
rect 900 2388 906 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2406 2388 2412 2440
rect 2464 2388 2470 2440
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 992 2332 1409 2360
rect 992 2320 998 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 10060 2360 10088 2468
rect 10318 2388 10324 2440
rect 10376 2388 10382 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11333 2431 11391 2437
rect 10919 2400 11008 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 1811 2332 10088 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 10980 2304 11008 2400
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 11422 2428 11428 2440
rect 11379 2400 11428 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11572 2400 11621 2428
rect 11572 2388 11578 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 11146 2320 11152 2372
rect 11204 2360 11210 2372
rect 12084 2360 12112 2391
rect 11204 2332 12112 2360
rect 11204 2320 11210 2332
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10686 2292 10692 2304
rect 10551 2264 10692 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 10778 2252 10784 2304
rect 10836 2252 10842 2304
rect 10962 2252 10968 2304
rect 11020 2252 11026 2304
rect 11241 2295 11299 2301
rect 11241 2261 11253 2295
rect 11287 2292 11299 2295
rect 11790 2292 11796 2304
rect 11287 2264 11796 2292
rect 11287 2261 11299 2264
rect 11241 2255 11299 2261
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 12268 2292 12296 2468
rect 12544 2468 13032 2496
rect 12544 2440 12572 2468
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 13004 2437 13032 2468
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13464 2360 13492 2391
rect 13906 2388 13912 2440
rect 13964 2388 13970 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 14148 2400 14381 2428
rect 14148 2388 14154 2400
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2428 14795 2431
rect 14844 2428 14872 2527
rect 15102 2524 15108 2576
rect 15160 2524 15166 2576
rect 16574 2496 16580 2508
rect 15028 2468 16580 2496
rect 15028 2437 15056 2468
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 14783 2400 14872 2428
rect 15013 2431 15071 2437
rect 14783 2397 14795 2400
rect 14737 2391 14795 2397
rect 15013 2397 15025 2431
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 15194 2360 15200 2372
rect 12406 2332 12848 2360
rect 13464 2332 15200 2360
rect 12406 2292 12434 2332
rect 12820 2301 12848 2332
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 15304 2360 15332 2391
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 15838 2388 15844 2440
rect 15896 2388 15902 2440
rect 16114 2388 16120 2440
rect 16172 2388 16178 2440
rect 15304 2332 16344 2360
rect 16316 2304 16344 2332
rect 12268 2264 12434 2292
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13722 2252 13728 2304
rect 13780 2252 13786 2304
rect 15470 2252 15476 2304
rect 15528 2252 15534 2304
rect 16206 2252 16212 2304
rect 16264 2252 16270 2304
rect 16298 2252 16304 2304
rect 16356 2252 16362 2304
rect 1104 2202 16995 2224
rect 1104 2150 4882 2202
rect 4934 2150 4946 2202
rect 4998 2150 5010 2202
rect 5062 2150 5074 2202
rect 5126 2150 5138 2202
rect 5190 2150 8815 2202
rect 8867 2150 8879 2202
rect 8931 2150 8943 2202
rect 8995 2150 9007 2202
rect 9059 2150 9071 2202
rect 9123 2150 12748 2202
rect 12800 2150 12812 2202
rect 12864 2150 12876 2202
rect 12928 2150 12940 2202
rect 12992 2150 13004 2202
rect 13056 2150 16681 2202
rect 16733 2150 16745 2202
rect 16797 2150 16809 2202
rect 16861 2150 16873 2202
rect 16925 2150 16937 2202
rect 16989 2150 16995 2202
rect 1104 2128 16995 2150
rect 10778 2048 10784 2100
rect 10836 2048 10842 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 13722 2088 13728 2100
rect 11020 2060 13728 2088
rect 11020 2048 11026 2060
rect 13722 2048 13728 2060
rect 13780 2048 13786 2100
rect 15470 2048 15476 2100
rect 15528 2048 15534 2100
rect 15838 2048 15844 2100
rect 15896 2048 15902 2100
rect 16114 2048 16120 2100
rect 16172 2048 16178 2100
rect 16206 2048 16212 2100
rect 16264 2048 16270 2100
rect 10686 1912 10692 1964
rect 10744 1912 10750 1964
rect 10796 1952 10824 2048
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 15488 2020 15516 2048
rect 11480 1992 15516 2020
rect 11480 1980 11486 1992
rect 15856 1952 15884 2048
rect 10796 1924 15884 1952
rect 10704 1884 10732 1912
rect 16132 1884 16160 2048
rect 10704 1856 16160 1884
rect 9582 1776 9588 1828
rect 9640 1816 9646 1828
rect 16224 1816 16252 2048
rect 9640 1788 16252 1816
rect 9640 1776 9646 1788
<< via1 >>
rect 2916 15750 2968 15802
rect 2980 15750 3032 15802
rect 3044 15750 3096 15802
rect 3108 15750 3160 15802
rect 3172 15750 3224 15802
rect 6849 15750 6901 15802
rect 6913 15750 6965 15802
rect 6977 15750 7029 15802
rect 7041 15750 7093 15802
rect 7105 15750 7157 15802
rect 10782 15750 10834 15802
rect 10846 15750 10898 15802
rect 10910 15750 10962 15802
rect 10974 15750 11026 15802
rect 11038 15750 11090 15802
rect 14715 15750 14767 15802
rect 14779 15750 14831 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 940 15648 992 15700
rect 16672 15648 16724 15700
rect 16764 15648 16816 15700
rect 11612 15512 11664 15564
rect 13636 15512 13688 15564
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 2872 15444 2924 15496
rect 4344 15487 4396 15496
rect 4344 15453 4353 15487
rect 4353 15453 4387 15487
rect 4387 15453 4396 15487
rect 4344 15444 4396 15453
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 10508 15444 10560 15496
rect 12072 15444 12124 15496
rect 15200 15487 15252 15496
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 3792 15376 3844 15428
rect 15752 15376 15804 15428
rect 15936 15419 15988 15428
rect 15936 15385 15945 15419
rect 15945 15385 15979 15419
rect 15979 15385 15988 15419
rect 15936 15376 15988 15385
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 2780 15308 2832 15360
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 4528 15351 4580 15360
rect 4528 15317 4537 15351
rect 4537 15317 4571 15351
rect 4571 15317 4580 15351
rect 4528 15308 4580 15317
rect 6184 15308 6236 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 13728 15351 13780 15360
rect 13728 15317 13737 15351
rect 13737 15317 13771 15351
rect 13771 15317 13780 15351
rect 13728 15308 13780 15317
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 15108 15308 15160 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 4882 15206 4934 15258
rect 4946 15206 4998 15258
rect 5010 15206 5062 15258
rect 5074 15206 5126 15258
rect 5138 15206 5190 15258
rect 8815 15206 8867 15258
rect 8879 15206 8931 15258
rect 8943 15206 8995 15258
rect 9007 15206 9059 15258
rect 9071 15206 9123 15258
rect 12748 15206 12800 15258
rect 12812 15206 12864 15258
rect 12876 15206 12928 15258
rect 12940 15206 12992 15258
rect 13004 15206 13056 15258
rect 16681 15206 16733 15258
rect 16745 15206 16797 15258
rect 16809 15206 16861 15258
rect 16873 15206 16925 15258
rect 16937 15206 16989 15258
rect 1492 15147 1544 15156
rect 1492 15113 1501 15147
rect 1501 15113 1535 15147
rect 1535 15113 1544 15147
rect 1492 15104 1544 15113
rect 3056 15104 3108 15156
rect 3792 15104 3844 15156
rect 7656 15104 7708 15156
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 11612 15104 11664 15113
rect 13912 15104 13964 15156
rect 15660 15104 15712 15156
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 16488 15104 16540 15156
rect 1124 15036 1176 15088
rect 2872 15036 2924 15088
rect 5724 14968 5776 15020
rect 12164 15036 12216 15088
rect 9956 15011 10008 15020
rect 9956 14977 9965 15011
rect 9965 14977 9999 15011
rect 9999 14977 10008 15011
rect 9956 14968 10008 14977
rect 14004 14968 14056 15020
rect 14740 14968 14792 15020
rect 15016 14968 15068 15020
rect 15476 14968 15528 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 8116 14900 8168 14952
rect 15936 14900 15988 14952
rect 3700 14764 3752 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 14556 14764 14608 14816
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 2916 14662 2968 14714
rect 2980 14662 3032 14714
rect 3044 14662 3096 14714
rect 3108 14662 3160 14714
rect 3172 14662 3224 14714
rect 6849 14662 6901 14714
rect 6913 14662 6965 14714
rect 6977 14662 7029 14714
rect 7041 14662 7093 14714
rect 7105 14662 7157 14714
rect 10782 14662 10834 14714
rect 10846 14662 10898 14714
rect 10910 14662 10962 14714
rect 10974 14662 11026 14714
rect 11038 14662 11090 14714
rect 14715 14662 14767 14714
rect 14779 14662 14831 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 5724 14424 5776 14476
rect 10600 14560 10652 14612
rect 15108 14560 15160 14612
rect 15476 14560 15528 14612
rect 9220 14356 9272 14408
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 11520 14356 11572 14408
rect 12164 14356 12216 14408
rect 13728 14356 13780 14408
rect 940 14288 992 14340
rect 11428 14288 11480 14340
rect 13636 14288 13688 14340
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16488 14331 16540 14340
rect 16488 14297 16497 14331
rect 16497 14297 16531 14331
rect 16531 14297 16540 14331
rect 16488 14288 16540 14297
rect 10048 14220 10100 14272
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 12440 14220 12492 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 15476 14220 15528 14272
rect 15568 14263 15620 14272
rect 15568 14229 15577 14263
rect 15577 14229 15611 14263
rect 15611 14229 15620 14263
rect 15568 14220 15620 14229
rect 15752 14263 15804 14272
rect 15752 14229 15761 14263
rect 15761 14229 15795 14263
rect 15795 14229 15804 14263
rect 15752 14220 15804 14229
rect 4882 14118 4934 14170
rect 4946 14118 4998 14170
rect 5010 14118 5062 14170
rect 5074 14118 5126 14170
rect 5138 14118 5190 14170
rect 8815 14118 8867 14170
rect 8879 14118 8931 14170
rect 8943 14118 8995 14170
rect 9007 14118 9059 14170
rect 9071 14118 9123 14170
rect 12748 14118 12800 14170
rect 12812 14118 12864 14170
rect 12876 14118 12928 14170
rect 12940 14118 12992 14170
rect 13004 14118 13056 14170
rect 16681 14118 16733 14170
rect 16745 14118 16797 14170
rect 16809 14118 16861 14170
rect 16873 14118 16925 14170
rect 16937 14118 16989 14170
rect 9312 14016 9364 14068
rect 6184 13948 6236 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 10324 14016 10376 14068
rect 10508 14016 10560 14068
rect 10784 14016 10836 14068
rect 11428 13812 11480 13864
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14740 14016 14792 14068
rect 15752 14016 15804 14068
rect 12716 13812 12768 13864
rect 15292 13880 15344 13932
rect 16396 13880 16448 13932
rect 16488 13923 16540 13932
rect 16488 13889 16497 13923
rect 16497 13889 16531 13923
rect 16531 13889 16540 13923
rect 16488 13880 16540 13889
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13544 13676 13596 13728
rect 14280 13719 14332 13728
rect 14280 13685 14289 13719
rect 14289 13685 14323 13719
rect 14323 13685 14332 13719
rect 14280 13676 14332 13685
rect 14464 13676 14516 13728
rect 2916 13574 2968 13626
rect 2980 13574 3032 13626
rect 3044 13574 3096 13626
rect 3108 13574 3160 13626
rect 3172 13574 3224 13626
rect 6849 13574 6901 13626
rect 6913 13574 6965 13626
rect 6977 13574 7029 13626
rect 7041 13574 7093 13626
rect 7105 13574 7157 13626
rect 10782 13574 10834 13626
rect 10846 13574 10898 13626
rect 10910 13574 10962 13626
rect 10974 13574 11026 13626
rect 11038 13574 11090 13626
rect 14715 13574 14767 13626
rect 14779 13574 14831 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 9036 13472 9088 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 12992 13472 13044 13524
rect 15660 13515 15712 13524
rect 15660 13481 15669 13515
rect 15669 13481 15703 13515
rect 15703 13481 15712 13515
rect 15660 13472 15712 13481
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 9680 13268 9732 13320
rect 8484 13200 8536 13252
rect 10416 13336 10468 13388
rect 13636 13404 13688 13456
rect 14280 13404 14332 13456
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12808 13336 12860 13388
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 9864 13132 9916 13184
rect 11888 13243 11940 13252
rect 11888 13209 11897 13243
rect 11897 13209 11931 13243
rect 11931 13209 11940 13243
rect 11888 13200 11940 13209
rect 12256 13200 12308 13252
rect 12532 13132 12584 13184
rect 15292 13336 15344 13388
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 15476 13268 15528 13320
rect 16580 13268 16632 13320
rect 13544 13132 13596 13184
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 14464 13132 14516 13184
rect 4882 13030 4934 13082
rect 4946 13030 4998 13082
rect 5010 13030 5062 13082
rect 5074 13030 5126 13082
rect 5138 13030 5190 13082
rect 8815 13030 8867 13082
rect 8879 13030 8931 13082
rect 8943 13030 8995 13082
rect 9007 13030 9059 13082
rect 9071 13030 9123 13082
rect 12748 13030 12800 13082
rect 12812 13030 12864 13082
rect 12876 13030 12928 13082
rect 12940 13030 12992 13082
rect 13004 13030 13056 13082
rect 16681 13030 16733 13082
rect 16745 13030 16797 13082
rect 16809 13030 16861 13082
rect 16873 13030 16925 13082
rect 16937 13030 16989 13082
rect 1768 12928 1820 12980
rect 4528 12928 4580 12980
rect 3332 12792 3384 12844
rect 5356 12860 5408 12912
rect 8484 12928 8536 12980
rect 9220 12928 9272 12980
rect 9680 12928 9732 12980
rect 11888 12928 11940 12980
rect 13820 12928 13872 12980
rect 14372 12928 14424 12980
rect 14648 12928 14700 12980
rect 6184 12792 6236 12844
rect 9680 12792 9732 12844
rect 9864 12835 9916 12844
rect 9864 12801 9898 12835
rect 9898 12801 9916 12835
rect 9864 12792 9916 12801
rect 12164 12860 12216 12912
rect 8484 12724 8536 12776
rect 12624 12792 12676 12844
rect 13636 12792 13688 12844
rect 16120 12860 16172 12912
rect 13544 12767 13596 12776
rect 11520 12656 11572 12708
rect 940 12588 992 12640
rect 12624 12588 12676 12640
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14188 12724 14240 12776
rect 15200 12724 15252 12776
rect 15844 12724 15896 12776
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 2916 12486 2968 12538
rect 2980 12486 3032 12538
rect 3044 12486 3096 12538
rect 3108 12486 3160 12538
rect 3172 12486 3224 12538
rect 6849 12486 6901 12538
rect 6913 12486 6965 12538
rect 6977 12486 7029 12538
rect 7041 12486 7093 12538
rect 7105 12486 7157 12538
rect 10782 12486 10834 12538
rect 10846 12486 10898 12538
rect 10910 12486 10962 12538
rect 10974 12486 11026 12538
rect 11038 12486 11090 12538
rect 14715 12486 14767 12538
rect 14779 12486 14831 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 9312 12384 9364 12436
rect 12532 12384 12584 12436
rect 14372 12384 14424 12436
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 12532 12291 12584 12300
rect 4528 12180 4580 12232
rect 6920 12180 6972 12232
rect 9680 12180 9732 12232
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 15568 12248 15620 12300
rect 940 12112 992 12164
rect 10324 12112 10376 12164
rect 11612 12180 11664 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 15660 12180 15712 12232
rect 7472 12044 7524 12096
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11336 12044 11388 12053
rect 12992 12112 13044 12164
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 14372 12044 14424 12096
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 4882 11942 4934 11994
rect 4946 11942 4998 11994
rect 5010 11942 5062 11994
rect 5074 11942 5126 11994
rect 5138 11942 5190 11994
rect 8815 11942 8867 11994
rect 8879 11942 8931 11994
rect 8943 11942 8995 11994
rect 9007 11942 9059 11994
rect 9071 11942 9123 11994
rect 12748 11942 12800 11994
rect 12812 11942 12864 11994
rect 12876 11942 12928 11994
rect 12940 11942 12992 11994
rect 13004 11942 13056 11994
rect 16681 11942 16733 11994
rect 16745 11942 16797 11994
rect 16809 11942 16861 11994
rect 16873 11942 16925 11994
rect 16937 11942 16989 11994
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 9128 11840 9180 11892
rect 7472 11772 7524 11824
rect 9036 11815 9088 11824
rect 9036 11781 9045 11815
rect 9045 11781 9079 11815
rect 9079 11781 9088 11815
rect 9036 11772 9088 11781
rect 7380 11704 7432 11756
rect 7564 11747 7616 11756
rect 7564 11713 7598 11747
rect 7598 11713 7616 11747
rect 7564 11704 7616 11713
rect 10324 11883 10376 11892
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 10508 11840 10560 11892
rect 11980 11840 12032 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 12532 11704 12584 11756
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 14464 11772 14516 11824
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 6460 11636 6512 11688
rect 10140 11636 10192 11688
rect 10232 11636 10284 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 13268 11636 13320 11688
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 8208 11500 8260 11552
rect 11980 11568 12032 11620
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 15200 11500 15252 11552
rect 15568 11500 15620 11552
rect 2916 11398 2968 11450
rect 2980 11398 3032 11450
rect 3044 11398 3096 11450
rect 3108 11398 3160 11450
rect 3172 11398 3224 11450
rect 6849 11398 6901 11450
rect 6913 11398 6965 11450
rect 6977 11398 7029 11450
rect 7041 11398 7093 11450
rect 7105 11398 7157 11450
rect 10782 11398 10834 11450
rect 10846 11398 10898 11450
rect 10910 11398 10962 11450
rect 10974 11398 11026 11450
rect 11038 11398 11090 11450
rect 14715 11398 14767 11450
rect 14779 11398 14831 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 5632 11296 5684 11348
rect 7472 11339 7524 11348
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 9036 11339 9088 11348
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 9128 11296 9180 11348
rect 10416 11296 10468 11348
rect 11336 11296 11388 11348
rect 11704 11296 11756 11348
rect 15660 11296 15712 11348
rect 6920 11160 6972 11212
rect 2780 11092 2832 11144
rect 4712 11092 4764 11144
rect 1400 11067 1452 11076
rect 1400 11033 1409 11067
rect 1409 11033 1443 11067
rect 1443 11033 1452 11067
rect 1400 11024 1452 11033
rect 7472 11092 7524 11144
rect 8300 11024 8352 11076
rect 9680 11024 9732 11076
rect 9956 11067 10008 11076
rect 9956 11033 9965 11067
rect 9965 11033 9999 11067
rect 9999 11033 10008 11067
rect 9956 11024 10008 11033
rect 4804 10956 4856 11008
rect 7012 10956 7064 11008
rect 9220 10956 9272 11008
rect 10140 11024 10192 11076
rect 10692 11024 10744 11076
rect 13912 11228 13964 11280
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 16120 11296 16172 11348
rect 13084 11092 13136 11144
rect 16212 11160 16264 11212
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 13728 11067 13780 11076
rect 13728 11033 13737 11067
rect 13737 11033 13771 11067
rect 13771 11033 13780 11067
rect 13728 11024 13780 11033
rect 13360 10956 13412 11008
rect 14188 11067 14240 11076
rect 14188 11033 14197 11067
rect 14197 11033 14231 11067
rect 14231 11033 14240 11067
rect 14188 11024 14240 11033
rect 14556 11067 14608 11076
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 15568 11024 15620 11076
rect 13912 10956 13964 11008
rect 14372 10956 14424 11008
rect 4882 10854 4934 10906
rect 4946 10854 4998 10906
rect 5010 10854 5062 10906
rect 5074 10854 5126 10906
rect 5138 10854 5190 10906
rect 8815 10854 8867 10906
rect 8879 10854 8931 10906
rect 8943 10854 8995 10906
rect 9007 10854 9059 10906
rect 9071 10854 9123 10906
rect 12748 10854 12800 10906
rect 12812 10854 12864 10906
rect 12876 10854 12928 10906
rect 12940 10854 12992 10906
rect 13004 10854 13056 10906
rect 16681 10854 16733 10906
rect 16745 10854 16797 10906
rect 16809 10854 16861 10906
rect 16873 10854 16925 10906
rect 16937 10854 16989 10906
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 6920 10752 6972 10804
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 8208 10752 8260 10804
rect 7012 10727 7064 10736
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 940 10412 992 10464
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 6644 10616 6696 10668
rect 8944 10616 8996 10668
rect 9128 10616 9180 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9496 10616 9548 10668
rect 9680 10616 9732 10668
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 13084 10752 13136 10804
rect 16304 10752 16356 10804
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 4528 10412 4580 10464
rect 9864 10548 9916 10600
rect 11980 10548 12032 10600
rect 12256 10616 12308 10668
rect 13820 10684 13872 10736
rect 14372 10684 14424 10736
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13360 10616 13412 10668
rect 15752 10727 15804 10736
rect 15752 10693 15761 10727
rect 15761 10693 15795 10727
rect 15795 10693 15804 10727
rect 15752 10684 15804 10693
rect 13728 10548 13780 10600
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 13544 10480 13596 10532
rect 14372 10480 14424 10532
rect 15936 10548 15988 10600
rect 7380 10412 7432 10464
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9956 10412 10008 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 2916 10310 2968 10362
rect 2980 10310 3032 10362
rect 3044 10310 3096 10362
rect 3108 10310 3160 10362
rect 3172 10310 3224 10362
rect 6849 10310 6901 10362
rect 6913 10310 6965 10362
rect 6977 10310 7029 10362
rect 7041 10310 7093 10362
rect 7105 10310 7157 10362
rect 10782 10310 10834 10362
rect 10846 10310 10898 10362
rect 10910 10310 10962 10362
rect 10974 10310 11026 10362
rect 11038 10310 11090 10362
rect 14715 10310 14767 10362
rect 14779 10310 14831 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 6000 10208 6052 10260
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 9312 10208 9364 10260
rect 6644 10140 6696 10192
rect 6828 10140 6880 10192
rect 4804 10072 4856 10124
rect 6552 10072 6604 10124
rect 9864 10140 9916 10192
rect 12532 10208 12584 10260
rect 14372 10208 14424 10260
rect 2780 10004 2832 10056
rect 4712 10004 4764 10056
rect 5816 10049 5868 10056
rect 5816 10015 5825 10049
rect 5825 10015 5859 10049
rect 5859 10015 5868 10049
rect 5816 10004 5868 10015
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 8116 10072 8168 10124
rect 8392 10004 8444 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 5264 9868 5316 9920
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 6000 9868 6052 9920
rect 8668 9936 8720 9988
rect 9128 9936 9180 9988
rect 10416 9979 10468 9988
rect 10416 9945 10425 9979
rect 10425 9945 10459 9979
rect 10459 9945 10468 9979
rect 10416 9936 10468 9945
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 13544 10004 13596 10056
rect 13820 10072 13872 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 14464 10072 14516 10124
rect 15660 10072 15712 10124
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 13268 9936 13320 9988
rect 15292 9936 15344 9988
rect 16212 9979 16264 9988
rect 16212 9945 16221 9979
rect 16221 9945 16255 9979
rect 16255 9945 16264 9979
rect 16212 9936 16264 9945
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 9772 9868 9824 9920
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 13544 9868 13596 9920
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 4882 9766 4934 9818
rect 4946 9766 4998 9818
rect 5010 9766 5062 9818
rect 5074 9766 5126 9818
rect 5138 9766 5190 9818
rect 8815 9766 8867 9818
rect 8879 9766 8931 9818
rect 8943 9766 8995 9818
rect 9007 9766 9059 9818
rect 9071 9766 9123 9818
rect 12748 9766 12800 9818
rect 12812 9766 12864 9818
rect 12876 9766 12928 9818
rect 12940 9766 12992 9818
rect 13004 9766 13056 9818
rect 16681 9766 16733 9818
rect 16745 9766 16797 9818
rect 16809 9766 16861 9818
rect 16873 9766 16925 9818
rect 16937 9766 16989 9818
rect 4436 9596 4488 9648
rect 5448 9596 5500 9648
rect 5724 9596 5776 9648
rect 6276 9664 6328 9716
rect 7288 9664 7340 9716
rect 4988 9528 5040 9580
rect 2780 9392 2832 9444
rect 5264 9460 5316 9512
rect 6460 9528 6512 9580
rect 7196 9528 7248 9580
rect 7564 9528 7616 9580
rect 8576 9664 8628 9716
rect 8300 9596 8352 9648
rect 7932 9460 7984 9512
rect 8668 9596 8720 9648
rect 5724 9392 5776 9444
rect 9864 9528 9916 9580
rect 13084 9596 13136 9648
rect 13176 9639 13228 9648
rect 15016 9664 15068 9716
rect 16304 9664 16356 9716
rect 13176 9605 13216 9639
rect 13216 9605 13228 9639
rect 13176 9596 13228 9605
rect 13360 9528 13412 9580
rect 13636 9528 13688 9580
rect 14556 9528 14608 9580
rect 15200 9528 15252 9580
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 6000 9324 6052 9376
rect 8392 9324 8444 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9588 9324 9640 9376
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 12348 9324 12400 9376
rect 12716 9324 12768 9376
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 16120 9324 16172 9376
rect 2916 9222 2968 9274
rect 2980 9222 3032 9274
rect 3044 9222 3096 9274
rect 3108 9222 3160 9274
rect 3172 9222 3224 9274
rect 6849 9222 6901 9274
rect 6913 9222 6965 9274
rect 6977 9222 7029 9274
rect 7041 9222 7093 9274
rect 7105 9222 7157 9274
rect 10782 9222 10834 9274
rect 10846 9222 10898 9274
rect 10910 9222 10962 9274
rect 10974 9222 11026 9274
rect 11038 9222 11090 9274
rect 14715 9222 14767 9274
rect 14779 9222 14831 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 3792 9120 3844 9172
rect 4620 9120 4672 9172
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 4988 9120 5040 9172
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 10416 9120 10468 9172
rect 12532 9120 12584 9172
rect 13176 9120 13228 9172
rect 13544 9120 13596 9172
rect 5816 9052 5868 9104
rect 6828 9052 6880 9104
rect 7380 9052 7432 9104
rect 8668 9052 8720 9104
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 5908 8916 5960 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 7196 8916 7248 8968
rect 940 8848 992 8900
rect 5356 8848 5408 8900
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 5540 8891 5592 8900
rect 5540 8857 5549 8891
rect 5549 8857 5583 8891
rect 5583 8857 5592 8891
rect 5540 8848 5592 8857
rect 8484 8916 8536 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12440 9052 12492 9104
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 12624 8916 12676 8968
rect 14556 8984 14608 9036
rect 14188 8916 14240 8968
rect 16120 9120 16172 9172
rect 16764 9120 16816 9172
rect 15292 9095 15344 9104
rect 15292 9061 15301 9095
rect 15301 9061 15335 9095
rect 15335 9061 15344 9095
rect 15292 9052 15344 9061
rect 15476 9052 15528 9104
rect 5816 8780 5868 8832
rect 10692 8780 10744 8832
rect 13820 8780 13872 8832
rect 14004 8780 14056 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 15568 8780 15620 8832
rect 16120 8891 16172 8900
rect 16120 8857 16129 8891
rect 16129 8857 16163 8891
rect 16163 8857 16172 8891
rect 16120 8848 16172 8857
rect 16212 8780 16264 8832
rect 4882 8678 4934 8730
rect 4946 8678 4998 8730
rect 5010 8678 5062 8730
rect 5074 8678 5126 8730
rect 5138 8678 5190 8730
rect 8815 8678 8867 8730
rect 8879 8678 8931 8730
rect 8943 8678 8995 8730
rect 9007 8678 9059 8730
rect 9071 8678 9123 8730
rect 12748 8678 12800 8730
rect 12812 8678 12864 8730
rect 12876 8678 12928 8730
rect 12940 8678 12992 8730
rect 13004 8678 13056 8730
rect 16681 8678 16733 8730
rect 16745 8678 16797 8730
rect 16809 8678 16861 8730
rect 16873 8678 16925 8730
rect 16937 8678 16989 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 2780 8576 2832 8628
rect 4160 8576 4212 8628
rect 5724 8576 5776 8628
rect 6092 8576 6144 8628
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 6276 8508 6328 8560
rect 6828 8508 6880 8560
rect 8484 8619 8536 8628
rect 8484 8585 8493 8619
rect 8493 8585 8527 8619
rect 8527 8585 8536 8619
rect 8484 8576 8536 8585
rect 8576 8576 8628 8628
rect 9680 8576 9732 8628
rect 9864 8576 9916 8628
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 3516 8279 3568 8288
rect 3516 8245 3525 8279
rect 3525 8245 3559 8279
rect 3559 8245 3568 8279
rect 3516 8236 3568 8245
rect 4160 8304 4212 8356
rect 5540 8304 5592 8356
rect 5816 8304 5868 8356
rect 6736 8372 6788 8424
rect 7380 8304 7432 8356
rect 7656 8372 7708 8424
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 9772 8440 9824 8492
rect 9680 8372 9732 8424
rect 10232 8372 10284 8424
rect 11520 8576 11572 8628
rect 12256 8576 12308 8628
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12440 8508 12492 8560
rect 13268 8576 13320 8628
rect 13544 8508 13596 8560
rect 13912 8576 13964 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 15476 8576 15528 8628
rect 16304 8576 16356 8628
rect 16396 8619 16448 8628
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 13820 8508 13872 8560
rect 11336 8304 11388 8356
rect 12532 8440 12584 8492
rect 12900 8483 12952 8492
rect 12440 8372 12492 8424
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14556 8440 14608 8492
rect 15752 8440 15804 8492
rect 13176 8304 13228 8356
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 16488 8372 16540 8424
rect 16120 8304 16172 8356
rect 16396 8304 16448 8356
rect 5724 8236 5776 8288
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 9404 8236 9456 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 13084 8236 13136 8288
rect 13360 8236 13412 8288
rect 14280 8236 14332 8288
rect 2916 8134 2968 8186
rect 2980 8134 3032 8186
rect 3044 8134 3096 8186
rect 3108 8134 3160 8186
rect 3172 8134 3224 8186
rect 6849 8134 6901 8186
rect 6913 8134 6965 8186
rect 6977 8134 7029 8186
rect 7041 8134 7093 8186
rect 7105 8134 7157 8186
rect 10782 8134 10834 8186
rect 10846 8134 10898 8186
rect 10910 8134 10962 8186
rect 10974 8134 11026 8186
rect 11038 8134 11090 8186
rect 14715 8134 14767 8186
rect 14779 8134 14831 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 4252 8032 4304 8084
rect 4988 8032 5040 8084
rect 5264 8032 5316 8084
rect 6460 8032 6512 8084
rect 7288 8032 7340 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 9404 7964 9456 8016
rect 11796 8032 11848 8084
rect 12624 8032 12676 8084
rect 12992 8032 13044 8084
rect 14096 8032 14148 8084
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 13912 7964 13964 8016
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3516 7828 3568 7880
rect 3792 7828 3844 7880
rect 4160 7828 4212 7880
rect 4620 7828 4672 7880
rect 940 7760 992 7812
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 5724 7760 5776 7812
rect 7196 7760 7248 7812
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 10324 7760 10376 7812
rect 10508 7803 10560 7812
rect 10508 7769 10517 7803
rect 10517 7769 10551 7803
rect 10551 7769 10560 7803
rect 10508 7760 10560 7769
rect 11152 7803 11204 7812
rect 11152 7769 11161 7803
rect 11161 7769 11195 7803
rect 11195 7769 11204 7803
rect 11152 7760 11204 7769
rect 11888 7760 11940 7812
rect 12992 7760 13044 7812
rect 13268 7803 13320 7812
rect 13268 7769 13277 7803
rect 13277 7769 13311 7803
rect 13311 7769 13320 7803
rect 13268 7760 13320 7769
rect 13360 7803 13412 7812
rect 13360 7769 13369 7803
rect 13369 7769 13403 7803
rect 13403 7769 13412 7803
rect 13360 7760 13412 7769
rect 13728 7760 13780 7812
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 17224 7828 17276 7880
rect 15568 7760 15620 7812
rect 17132 7760 17184 7812
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 14004 7692 14056 7744
rect 15384 7692 15436 7744
rect 4882 7590 4934 7642
rect 4946 7590 4998 7642
rect 5010 7590 5062 7642
rect 5074 7590 5126 7642
rect 5138 7590 5190 7642
rect 8815 7590 8867 7642
rect 8879 7590 8931 7642
rect 8943 7590 8995 7642
rect 9007 7590 9059 7642
rect 9071 7590 9123 7642
rect 12748 7590 12800 7642
rect 12812 7590 12864 7642
rect 12876 7590 12928 7642
rect 12940 7590 12992 7642
rect 13004 7590 13056 7642
rect 16681 7590 16733 7642
rect 16745 7590 16797 7642
rect 16809 7590 16861 7642
rect 16873 7590 16925 7642
rect 16937 7590 16989 7642
rect 3148 7488 3200 7540
rect 3332 7488 3384 7540
rect 4804 7488 4856 7540
rect 5816 7488 5868 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 3240 7284 3292 7336
rect 4528 7420 4580 7472
rect 5356 7352 5408 7404
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 7288 7488 7340 7540
rect 8116 7488 8168 7540
rect 8668 7488 8720 7540
rect 6736 7420 6788 7472
rect 6460 7352 6512 7404
rect 6644 7395 6696 7404
rect 6644 7361 6678 7395
rect 6678 7361 6696 7395
rect 6644 7352 6696 7361
rect 13268 7488 13320 7540
rect 14096 7488 14148 7540
rect 17040 7488 17092 7540
rect 10508 7463 10560 7472
rect 10508 7429 10517 7463
rect 10517 7429 10551 7463
rect 10551 7429 10560 7463
rect 10508 7420 10560 7429
rect 11152 7420 11204 7472
rect 13176 7420 13228 7472
rect 9128 7352 9180 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13728 7352 13780 7404
rect 15660 7420 15712 7472
rect 14188 7352 14240 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15752 7352 15804 7404
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 10692 7284 10744 7336
rect 11704 7284 11756 7336
rect 11888 7284 11940 7336
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 14096 7284 14148 7336
rect 15200 7284 15252 7336
rect 15568 7284 15620 7336
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 4620 7148 4672 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 6276 7148 6328 7200
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 16212 7284 16264 7336
rect 7840 7148 7892 7200
rect 8392 7148 8444 7200
rect 9680 7148 9732 7200
rect 10508 7148 10560 7200
rect 13544 7148 13596 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 2916 7046 2968 7098
rect 2980 7046 3032 7098
rect 3044 7046 3096 7098
rect 3108 7046 3160 7098
rect 3172 7046 3224 7098
rect 6849 7046 6901 7098
rect 6913 7046 6965 7098
rect 6977 7046 7029 7098
rect 7041 7046 7093 7098
rect 7105 7046 7157 7098
rect 10782 7046 10834 7098
rect 10846 7046 10898 7098
rect 10910 7046 10962 7098
rect 10974 7046 11026 7098
rect 11038 7046 11090 7098
rect 14715 7046 14767 7098
rect 14779 7046 14831 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 1768 6944 1820 6996
rect 5448 6876 5500 6928
rect 6644 6944 6696 6996
rect 8116 6944 8168 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 11152 6944 11204 6996
rect 3700 6808 3752 6860
rect 4620 6808 4672 6860
rect 4252 6740 4304 6792
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 3056 6672 3108 6681
rect 4068 6604 4120 6656
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 8668 6876 8720 6928
rect 11612 6944 11664 6996
rect 13268 6944 13320 6996
rect 13360 6944 13412 6996
rect 14924 6944 14976 6996
rect 4712 6740 4764 6749
rect 5540 6740 5592 6792
rect 6460 6740 6512 6792
rect 9588 6808 9640 6860
rect 7288 6740 7340 6792
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 10508 6808 10560 6860
rect 11428 6876 11480 6928
rect 11336 6808 11388 6860
rect 12348 6808 12400 6860
rect 13544 6808 13596 6860
rect 13636 6808 13688 6860
rect 7840 6672 7892 6724
rect 11152 6672 11204 6724
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 11520 6672 11572 6724
rect 12072 6672 12124 6724
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 13728 6740 13780 6792
rect 14188 6876 14240 6928
rect 14740 6876 14792 6928
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 14372 6808 14424 6860
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 15016 6876 15068 6928
rect 15384 6876 15436 6928
rect 14004 6740 14056 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 13636 6672 13688 6724
rect 4804 6604 4856 6656
rect 5908 6604 5960 6656
rect 9772 6604 9824 6656
rect 11060 6604 11112 6656
rect 12164 6604 12216 6656
rect 12532 6604 12584 6656
rect 12624 6604 12676 6656
rect 14096 6672 14148 6724
rect 15016 6672 15068 6724
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 15568 6604 15620 6656
rect 15660 6604 15712 6656
rect 4882 6502 4934 6554
rect 4946 6502 4998 6554
rect 5010 6502 5062 6554
rect 5074 6502 5126 6554
rect 5138 6502 5190 6554
rect 8815 6502 8867 6554
rect 8879 6502 8931 6554
rect 8943 6502 8995 6554
rect 9007 6502 9059 6554
rect 9071 6502 9123 6554
rect 12748 6502 12800 6554
rect 12812 6502 12864 6554
rect 12876 6502 12928 6554
rect 12940 6502 12992 6554
rect 13004 6502 13056 6554
rect 16681 6502 16733 6554
rect 16745 6502 16797 6554
rect 16809 6502 16861 6554
rect 16873 6502 16925 6554
rect 16937 6502 16989 6554
rect 3056 6400 3108 6452
rect 4620 6400 4672 6452
rect 4804 6400 4856 6452
rect 5080 6332 5132 6384
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 5908 6307 5960 6316
rect 5908 6273 5926 6307
rect 5926 6273 5960 6307
rect 5908 6264 5960 6273
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 6276 6264 6328 6316
rect 7380 6400 7432 6452
rect 7748 6400 7800 6452
rect 7840 6443 7892 6452
rect 7840 6409 7849 6443
rect 7849 6409 7883 6443
rect 7883 6409 7892 6443
rect 7840 6400 7892 6409
rect 8392 6400 8444 6452
rect 10692 6400 10744 6452
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 4436 6196 4488 6248
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 8576 6264 8628 6316
rect 940 6060 992 6112
rect 4712 6060 4764 6112
rect 8208 6128 8260 6180
rect 11060 6332 11112 6384
rect 11612 6400 11664 6452
rect 14832 6400 14884 6452
rect 15476 6400 15528 6452
rect 15844 6400 15896 6452
rect 16580 6400 16632 6452
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 8668 6060 8720 6112
rect 9220 6264 9272 6316
rect 9864 6264 9916 6316
rect 12992 6375 13044 6384
rect 12992 6341 13001 6375
rect 13001 6341 13035 6375
rect 13035 6341 13044 6375
rect 12992 6332 13044 6341
rect 14280 6332 14332 6384
rect 14372 6375 14424 6384
rect 14372 6341 14381 6375
rect 14381 6341 14415 6375
rect 14415 6341 14424 6375
rect 14372 6332 14424 6341
rect 14648 6332 14700 6384
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 11428 6196 11480 6248
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 11244 6128 11296 6180
rect 12900 6128 12952 6180
rect 9772 6060 9824 6112
rect 10048 6060 10100 6112
rect 11152 6060 11204 6112
rect 11888 6060 11940 6112
rect 14004 6196 14056 6248
rect 17040 6332 17092 6384
rect 14372 6196 14424 6248
rect 14556 6196 14608 6248
rect 15752 6264 15804 6316
rect 16120 6264 16172 6316
rect 16212 6196 16264 6248
rect 16580 6196 16632 6248
rect 13820 6128 13872 6180
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 13728 6060 13780 6112
rect 14924 6060 14976 6112
rect 2916 5958 2968 6010
rect 2980 5958 3032 6010
rect 3044 5958 3096 6010
rect 3108 5958 3160 6010
rect 3172 5958 3224 6010
rect 6849 5958 6901 6010
rect 6913 5958 6965 6010
rect 6977 5958 7029 6010
rect 7041 5958 7093 6010
rect 7105 5958 7157 6010
rect 10782 5958 10834 6010
rect 10846 5958 10898 6010
rect 10910 5958 10962 6010
rect 10974 5958 11026 6010
rect 11038 5958 11090 6010
rect 14715 5958 14767 6010
rect 14779 5958 14831 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 5080 5856 5132 5908
rect 5540 5856 5592 5908
rect 8300 5856 8352 5908
rect 5724 5720 5776 5772
rect 7196 5720 7248 5772
rect 7840 5720 7892 5772
rect 8024 5720 8076 5772
rect 8944 5831 8996 5840
rect 8944 5797 8953 5831
rect 8953 5797 8987 5831
rect 8987 5797 8996 5831
rect 8944 5788 8996 5797
rect 9128 5788 9180 5840
rect 9312 5788 9364 5840
rect 10324 5788 10376 5840
rect 8668 5720 8720 5772
rect 10600 5856 10652 5908
rect 11612 5856 11664 5908
rect 11796 5856 11848 5908
rect 11980 5856 12032 5908
rect 12992 5856 13044 5908
rect 13268 5856 13320 5908
rect 13820 5856 13872 5908
rect 12532 5788 12584 5840
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 12072 5720 12124 5772
rect 12164 5720 12216 5772
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 7288 5652 7340 5704
rect 8208 5652 8260 5704
rect 4252 5584 4304 5636
rect 6920 5584 6972 5636
rect 4160 5516 4212 5568
rect 6184 5516 6236 5568
rect 7196 5516 7248 5568
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 10048 5652 10100 5704
rect 9496 5627 9548 5636
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 8484 5516 8536 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 12624 5720 12676 5772
rect 12900 5720 12952 5772
rect 15660 5788 15712 5840
rect 16212 5788 16264 5840
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 14004 5652 14056 5704
rect 14464 5652 14516 5704
rect 15384 5652 15436 5704
rect 13820 5584 13872 5636
rect 15660 5652 15712 5704
rect 16120 5652 16172 5704
rect 11336 5516 11388 5568
rect 15476 5584 15528 5636
rect 16580 5584 16632 5636
rect 14372 5516 14424 5568
rect 4882 5414 4934 5466
rect 4946 5414 4998 5466
rect 5010 5414 5062 5466
rect 5074 5414 5126 5466
rect 5138 5414 5190 5466
rect 8815 5414 8867 5466
rect 8879 5414 8931 5466
rect 8943 5414 8995 5466
rect 9007 5414 9059 5466
rect 9071 5414 9123 5466
rect 12748 5414 12800 5466
rect 12812 5414 12864 5466
rect 12876 5414 12928 5466
rect 12940 5414 12992 5466
rect 13004 5414 13056 5466
rect 16681 5414 16733 5466
rect 16745 5414 16797 5466
rect 16809 5414 16861 5466
rect 16873 5414 16925 5466
rect 16937 5414 16989 5466
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 4620 5312 4672 5364
rect 5080 5312 5132 5364
rect 8484 5312 8536 5364
rect 5448 5287 5500 5296
rect 5448 5253 5457 5287
rect 5457 5253 5491 5287
rect 5491 5253 5500 5287
rect 5448 5244 5500 5253
rect 6920 5244 6972 5296
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4344 5176 4396 5228
rect 5080 5176 5132 5228
rect 5724 5040 5776 5092
rect 6552 5108 6604 5160
rect 6736 5108 6788 5160
rect 7380 5176 7432 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8944 5287 8996 5296
rect 8944 5253 8953 5287
rect 8953 5253 8987 5287
rect 8987 5253 8996 5287
rect 8944 5244 8996 5253
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 12256 5312 12308 5364
rect 8760 5176 8812 5228
rect 9312 5176 9364 5228
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 9680 5176 9732 5228
rect 10324 5176 10376 5228
rect 11520 5176 11572 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12072 5244 12124 5296
rect 13820 5312 13872 5364
rect 14556 5312 14608 5364
rect 16304 5312 16356 5364
rect 16488 5312 16540 5364
rect 12532 5176 12584 5228
rect 8484 5040 8536 5092
rect 8668 5108 8720 5160
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 9128 5040 9180 5092
rect 11428 5040 11480 5092
rect 4344 4972 4396 5024
rect 5540 4972 5592 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 8576 4972 8628 5024
rect 8852 4972 8904 5024
rect 11244 4972 11296 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 13728 5040 13780 5092
rect 14556 5176 14608 5228
rect 15476 5176 15528 5228
rect 15752 5176 15804 5228
rect 15200 5151 15252 5160
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 15292 5108 15344 5160
rect 16120 5108 16172 5160
rect 16396 5176 16448 5228
rect 16580 5108 16632 5160
rect 14188 4972 14240 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 2916 4870 2968 4922
rect 2980 4870 3032 4922
rect 3044 4870 3096 4922
rect 3108 4870 3160 4922
rect 3172 4870 3224 4922
rect 6849 4870 6901 4922
rect 6913 4870 6965 4922
rect 6977 4870 7029 4922
rect 7041 4870 7093 4922
rect 7105 4870 7157 4922
rect 10782 4870 10834 4922
rect 10846 4870 10898 4922
rect 10910 4870 10962 4922
rect 10974 4870 11026 4922
rect 11038 4870 11090 4922
rect 14715 4870 14767 4922
rect 14779 4870 14831 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 6368 4768 6420 4820
rect 8852 4768 8904 4820
rect 5724 4700 5776 4752
rect 8024 4632 8076 4684
rect 9220 4768 9272 4820
rect 10416 4768 10468 4820
rect 13728 4768 13780 4820
rect 15200 4768 15252 4820
rect 14188 4700 14240 4752
rect 14280 4632 14332 4684
rect 14648 4632 14700 4684
rect 4344 4564 4396 4616
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 7104 4564 7156 4616
rect 8300 4564 8352 4616
rect 940 4496 992 4548
rect 5264 4496 5316 4548
rect 5540 4539 5592 4548
rect 5540 4505 5549 4539
rect 5549 4505 5583 4539
rect 5583 4505 5592 4539
rect 5540 4496 5592 4505
rect 4160 4428 4212 4480
rect 8668 4428 8720 4480
rect 12532 4564 12584 4616
rect 13084 4564 13136 4616
rect 13544 4564 13596 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 16028 4632 16080 4684
rect 9588 4496 9640 4548
rect 9312 4428 9364 4480
rect 11428 4428 11480 4480
rect 12072 4496 12124 4548
rect 13360 4428 13412 4480
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 13912 4428 13964 4437
rect 14556 4564 14608 4616
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15384 4564 15436 4616
rect 15752 4564 15804 4616
rect 4882 4326 4934 4378
rect 4946 4326 4998 4378
rect 5010 4326 5062 4378
rect 5074 4326 5126 4378
rect 5138 4326 5190 4378
rect 8815 4326 8867 4378
rect 8879 4326 8931 4378
rect 8943 4326 8995 4378
rect 9007 4326 9059 4378
rect 9071 4326 9123 4378
rect 12748 4326 12800 4378
rect 12812 4326 12864 4378
rect 12876 4326 12928 4378
rect 12940 4326 12992 4378
rect 13004 4326 13056 4378
rect 16681 4326 16733 4378
rect 16745 4326 16797 4378
rect 16809 4326 16861 4378
rect 16873 4326 16925 4378
rect 16937 4326 16989 4378
rect 4160 4224 4212 4276
rect 4344 4224 4396 4276
rect 4804 4224 4856 4276
rect 5264 4267 5316 4276
rect 5264 4233 5273 4267
rect 5273 4233 5307 4267
rect 5307 4233 5316 4267
rect 5264 4224 5316 4233
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7840 4224 7892 4276
rect 3792 4156 3844 4208
rect 4068 4020 4120 4072
rect 5540 4088 5592 4140
rect 6276 4088 6328 4140
rect 6736 4088 6788 4140
rect 7472 4131 7524 4140
rect 7472 4097 7490 4131
rect 7490 4097 7524 4131
rect 8576 4224 8628 4276
rect 12072 4267 12124 4276
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 13084 4224 13136 4276
rect 7472 4088 7524 4097
rect 8024 4088 8076 4140
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8300 4020 8352 4029
rect 11428 4156 11480 4208
rect 10784 4088 10836 4140
rect 11520 4088 11572 4140
rect 12164 4088 12216 4140
rect 14280 4224 14332 4276
rect 14924 4224 14976 4276
rect 15476 4224 15528 4276
rect 6552 3952 6604 4004
rect 9220 4020 9272 4072
rect 9956 4020 10008 4072
rect 11244 4020 11296 4072
rect 11704 4020 11756 4072
rect 13360 4088 13412 4140
rect 13912 4088 13964 4140
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14648 4156 14700 4208
rect 940 3884 992 3936
rect 7472 3884 7524 3936
rect 9496 3884 9548 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 10784 3884 10836 3936
rect 12992 4020 13044 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 14648 4020 14700 4072
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16212 4088 16264 4140
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 15752 4020 15804 4029
rect 16028 4020 16080 4072
rect 13728 3952 13780 4004
rect 14280 3952 14332 4004
rect 13268 3884 13320 3936
rect 16212 3884 16264 3936
rect 2916 3782 2968 3834
rect 2980 3782 3032 3834
rect 3044 3782 3096 3834
rect 3108 3782 3160 3834
rect 3172 3782 3224 3834
rect 6849 3782 6901 3834
rect 6913 3782 6965 3834
rect 6977 3782 7029 3834
rect 7041 3782 7093 3834
rect 7105 3782 7157 3834
rect 10782 3782 10834 3834
rect 10846 3782 10898 3834
rect 10910 3782 10962 3834
rect 10974 3782 11026 3834
rect 11038 3782 11090 3834
rect 14715 3782 14767 3834
rect 14779 3782 14831 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 9588 3723 9640 3732
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 10324 3680 10376 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 13268 3680 13320 3732
rect 14556 3723 14608 3732
rect 14556 3689 14565 3723
rect 14565 3689 14599 3723
rect 14599 3689 14608 3723
rect 14556 3680 14608 3689
rect 15384 3680 15436 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 8300 3612 8352 3664
rect 4068 3544 4120 3596
rect 6368 3476 6420 3528
rect 10692 3544 10744 3596
rect 11520 3544 11572 3596
rect 12992 3544 13044 3596
rect 14464 3612 14516 3664
rect 6920 3408 6972 3460
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 7472 3408 7524 3460
rect 8668 3476 8720 3528
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 10416 3408 10468 3460
rect 12440 3408 12492 3460
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 13636 3476 13688 3528
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 14556 3476 14608 3528
rect 15844 3476 15896 3528
rect 17132 3476 17184 3528
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 12256 3383 12308 3392
rect 12256 3349 12265 3383
rect 12265 3349 12299 3383
rect 12299 3349 12308 3383
rect 12256 3340 12308 3349
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 14556 3340 14608 3392
rect 14832 3383 14884 3392
rect 14832 3349 14841 3383
rect 14841 3349 14875 3383
rect 14875 3349 14884 3383
rect 14832 3340 14884 3349
rect 4882 3238 4934 3290
rect 4946 3238 4998 3290
rect 5010 3238 5062 3290
rect 5074 3238 5126 3290
rect 5138 3238 5190 3290
rect 8815 3238 8867 3290
rect 8879 3238 8931 3290
rect 8943 3238 8995 3290
rect 9007 3238 9059 3290
rect 9071 3238 9123 3290
rect 12748 3238 12800 3290
rect 12812 3238 12864 3290
rect 12876 3238 12928 3290
rect 12940 3238 12992 3290
rect 13004 3238 13056 3290
rect 16681 3238 16733 3290
rect 16745 3238 16797 3290
rect 16809 3238 16861 3290
rect 16873 3238 16925 3290
rect 16937 3238 16989 3290
rect 3240 3136 3292 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 7012 3136 7064 3188
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 8116 3136 8168 3188
rect 8392 3136 8444 3188
rect 11520 3136 11572 3188
rect 11888 3136 11940 3188
rect 12256 3136 12308 3188
rect 12624 3136 12676 3188
rect 12900 3136 12952 3188
rect 13084 3136 13136 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13636 3136 13688 3188
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 15200 3136 15252 3188
rect 15292 3136 15344 3188
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 17224 3136 17276 3188
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 7932 3068 7984 3120
rect 2596 2932 2648 2984
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 11704 3068 11756 3120
rect 11428 3000 11480 3052
rect 11612 2932 11664 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 13360 3043 13412 3052
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 13360 3000 13412 3009
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14832 3000 14884 3052
rect 16212 3000 16264 3052
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 12532 2932 12584 2941
rect 940 2796 992 2848
rect 11336 2839 11388 2848
rect 11336 2805 11345 2839
rect 11345 2805 11379 2839
rect 11379 2805 11388 2839
rect 11336 2796 11388 2805
rect 11704 2796 11756 2848
rect 15108 2796 15160 2848
rect 2916 2694 2968 2746
rect 2980 2694 3032 2746
rect 3044 2694 3096 2746
rect 3108 2694 3160 2746
rect 3172 2694 3224 2746
rect 6849 2694 6901 2746
rect 6913 2694 6965 2746
rect 6977 2694 7029 2746
rect 7041 2694 7093 2746
rect 7105 2694 7157 2746
rect 10782 2694 10834 2746
rect 10846 2694 10898 2746
rect 10910 2694 10962 2746
rect 10974 2694 11026 2746
rect 11038 2694 11090 2746
rect 14715 2694 14767 2746
rect 14779 2694 14831 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 2780 2592 2832 2644
rect 4068 2635 4120 2644
rect 4068 2601 4077 2635
rect 4077 2601 4111 2635
rect 4111 2601 4120 2635
rect 4068 2592 4120 2601
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 7564 2592 7616 2644
rect 9312 2592 9364 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 11428 2592 11480 2644
rect 11612 2592 11664 2644
rect 12072 2592 12124 2644
rect 12532 2592 12584 2644
rect 13360 2592 13412 2644
rect 14004 2592 14056 2644
rect 14372 2592 14424 2644
rect 15752 2592 15804 2644
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 6644 2456 6696 2508
rect 848 2388 900 2440
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9588 2388 9640 2440
rect 9680 2388 9732 2440
rect 940 2320 992 2372
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11428 2388 11480 2440
rect 11520 2388 11572 2440
rect 11152 2320 11204 2372
rect 10692 2252 10744 2304
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 10968 2252 11020 2304
rect 11796 2252 11848 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 12532 2388 12584 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14096 2388 14148 2440
rect 15108 2567 15160 2576
rect 15108 2533 15117 2567
rect 15117 2533 15151 2567
rect 15151 2533 15160 2567
rect 15108 2524 15160 2533
rect 16580 2456 16632 2508
rect 15200 2320 15252 2372
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 16212 2295 16264 2304
rect 16212 2261 16221 2295
rect 16221 2261 16255 2295
rect 16255 2261 16264 2295
rect 16212 2252 16264 2261
rect 16304 2252 16356 2304
rect 4882 2150 4934 2202
rect 4946 2150 4998 2202
rect 5010 2150 5062 2202
rect 5074 2150 5126 2202
rect 5138 2150 5190 2202
rect 8815 2150 8867 2202
rect 8879 2150 8931 2202
rect 8943 2150 8995 2202
rect 9007 2150 9059 2202
rect 9071 2150 9123 2202
rect 12748 2150 12800 2202
rect 12812 2150 12864 2202
rect 12876 2150 12928 2202
rect 12940 2150 12992 2202
rect 13004 2150 13056 2202
rect 16681 2150 16733 2202
rect 16745 2150 16797 2202
rect 16809 2150 16861 2202
rect 16873 2150 16925 2202
rect 16937 2150 16989 2202
rect 10784 2048 10836 2100
rect 10968 2048 11020 2100
rect 13728 2048 13780 2100
rect 15476 2048 15528 2100
rect 15844 2048 15896 2100
rect 16120 2048 16172 2100
rect 16212 2048 16264 2100
rect 10692 1912 10744 1964
rect 11428 1980 11480 2032
rect 9588 1776 9640 1828
<< metal2 >>
rect 1122 17200 1178 18000
rect 2686 17200 2742 18000
rect 4250 17200 4306 18000
rect 5814 17200 5870 18000
rect 7378 17200 7434 18000
rect 8942 17200 8998 18000
rect 10506 17200 10562 18000
rect 12070 17200 12126 18000
rect 13634 17200 13690 18000
rect 14922 17504 14978 17513
rect 14978 17462 15148 17490
rect 14922 17439 14978 17448
rect 938 15872 994 15881
rect 938 15807 994 15816
rect 952 15706 980 15807
rect 940 15700 992 15706
rect 940 15642 992 15648
rect 1136 15094 1164 17200
rect 1490 16688 1546 16697
rect 1490 16623 1546 16632
rect 1504 15162 1532 16623
rect 2700 16574 2728 17200
rect 4264 16574 4292 17200
rect 5828 16574 5856 17200
rect 7392 16574 7420 17200
rect 8956 16574 8984 17200
rect 2700 16546 2820 16574
rect 4264 16546 4384 16574
rect 5828 16546 5948 16574
rect 7392 16546 7512 16574
rect 8956 16546 9076 16574
rect 2792 15502 2820 16546
rect 2916 15804 3224 15813
rect 2916 15802 2922 15804
rect 2978 15802 3002 15804
rect 3058 15802 3082 15804
rect 3138 15802 3162 15804
rect 3218 15802 3224 15804
rect 2978 15750 2980 15802
rect 3160 15750 3162 15802
rect 2916 15748 2922 15750
rect 2978 15748 3002 15750
rect 3058 15748 3082 15750
rect 3138 15748 3162 15750
rect 3218 15748 3224 15750
rect 2916 15739 3224 15748
rect 4356 15502 4384 16546
rect 5920 15502 5948 16546
rect 6849 15804 7157 15813
rect 6849 15802 6855 15804
rect 6911 15802 6935 15804
rect 6991 15802 7015 15804
rect 7071 15802 7095 15804
rect 7151 15802 7157 15804
rect 6911 15750 6913 15802
rect 7093 15750 7095 15802
rect 6849 15748 6855 15750
rect 6911 15748 6935 15750
rect 6991 15748 7015 15750
rect 7071 15748 7095 15750
rect 7151 15748 7157 15750
rect 6849 15739 7157 15748
rect 7484 15502 7512 16546
rect 9048 15502 9076 16546
rect 10520 15502 10548 17200
rect 10782 15804 11090 15813
rect 10782 15802 10788 15804
rect 10844 15802 10868 15804
rect 10924 15802 10948 15804
rect 11004 15802 11028 15804
rect 11084 15802 11090 15804
rect 10844 15750 10846 15802
rect 11026 15750 11028 15802
rect 10782 15748 10788 15750
rect 10844 15748 10868 15750
rect 10924 15748 10948 15750
rect 11004 15748 11028 15750
rect 11084 15748 11090 15750
rect 10782 15739 11090 15748
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2240 15201 2268 15302
rect 2226 15192 2282 15201
rect 1492 15156 1544 15162
rect 2226 15127 2282 15136
rect 1492 15098 1544 15104
rect 1124 15088 1176 15094
rect 1124 15030 1176 15036
rect 940 14340 992 14346
rect 940 14282 992 14288
rect 952 14249 980 14282
rect 938 14240 994 14249
rect 938 14175 994 14184
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13705 1532 13806
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1780 12986 1808 13874
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 940 12640 992 12646
rect 938 12608 940 12617
rect 992 12608 994 12617
rect 938 12543 994 12552
rect 940 12164 992 12170
rect 940 12106 992 12112
rect 952 11801 980 12106
rect 938 11792 994 11801
rect 938 11727 994 11736
rect 2792 11150 2820 15302
rect 2884 15094 2912 15438
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 15162 3096 15302
rect 3804 15162 3832 15370
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 2916 14716 3224 14725
rect 2916 14714 2922 14716
rect 2978 14714 3002 14716
rect 3058 14714 3082 14716
rect 3138 14714 3162 14716
rect 3218 14714 3224 14716
rect 2978 14662 2980 14714
rect 3160 14662 3162 14714
rect 2916 14660 2922 14662
rect 2978 14660 3002 14662
rect 3058 14660 3082 14662
rect 3138 14660 3162 14662
rect 3218 14660 3224 14662
rect 2916 14651 3224 14660
rect 2916 13628 3224 13637
rect 2916 13626 2922 13628
rect 2978 13626 3002 13628
rect 3058 13626 3082 13628
rect 3138 13626 3162 13628
rect 3218 13626 3224 13628
rect 2978 13574 2980 13626
rect 3160 13574 3162 13626
rect 2916 13572 2922 13574
rect 2978 13572 3002 13574
rect 3058 13572 3082 13574
rect 3138 13572 3162 13574
rect 3218 13572 3224 13574
rect 2916 13563 3224 13572
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 2916 12540 3224 12549
rect 2916 12538 2922 12540
rect 2978 12538 3002 12540
rect 3058 12538 3082 12540
rect 3138 12538 3162 12540
rect 3218 12538 3224 12540
rect 2978 12486 2980 12538
rect 3160 12486 3162 12538
rect 2916 12484 2922 12486
rect 2978 12484 3002 12486
rect 3058 12484 3082 12486
rect 3138 12484 3162 12486
rect 3218 12484 3224 12486
rect 2916 12475 3224 12484
rect 2916 11452 3224 11461
rect 2916 11450 2922 11452
rect 2978 11450 3002 11452
rect 3058 11450 3082 11452
rect 3138 11450 3162 11452
rect 3218 11450 3224 11452
rect 2978 11398 2980 11450
rect 3160 11398 3162 11450
rect 2916 11396 2922 11398
rect 2978 11396 3002 11398
rect 3058 11396 3082 11398
rect 3138 11396 3162 11398
rect 3218 11396 3224 11398
rect 2916 11387 3224 11396
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10985 1440 11018
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10169 980 10406
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8537 980 8842
rect 1780 8634 1808 10610
rect 2916 10364 3224 10373
rect 2916 10362 2922 10364
rect 2978 10362 3002 10364
rect 3058 10362 3082 10364
rect 3138 10362 3162 10364
rect 3218 10362 3224 10364
rect 2978 10310 2980 10362
rect 3160 10310 3162 10362
rect 2916 10308 2922 10310
rect 2978 10308 3002 10310
rect 3058 10308 3082 10310
rect 3138 10308 3162 10310
rect 3218 10308 3224 10310
rect 2916 10299 3224 10308
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9450 2820 9998
rect 3344 9625 3372 12786
rect 3330 9616 3386 9625
rect 3330 9551 3386 9560
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 8634 2820 9386
rect 2916 9276 3224 9285
rect 2916 9274 2922 9276
rect 2978 9274 3002 9276
rect 3058 9274 3082 9276
rect 3138 9274 3162 9276
rect 3218 9274 3224 9276
rect 2978 9222 2980 9274
rect 3160 9222 3162 9274
rect 2916 9220 2922 9222
rect 2978 9220 3002 9222
rect 3058 9220 3082 9222
rect 3138 9220 3162 9222
rect 3218 9220 3224 9222
rect 2916 9211 3224 9220
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 2916 8188 3224 8197
rect 2916 8186 2922 8188
rect 2978 8186 3002 8188
rect 3058 8186 3082 8188
rect 3138 8186 3162 8188
rect 3218 8186 3224 8188
rect 2978 8134 2980 8186
rect 3160 8134 3162 8186
rect 2916 8132 2922 8134
rect 2978 8132 3002 8134
rect 3058 8132 3082 8134
rect 3138 8132 3162 8134
rect 3218 8132 3224 8134
rect 2916 8123 3224 8132
rect 3528 7886 3556 8230
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7721 980 7754
rect 938 7712 994 7721
rect 938 7647 994 7656
rect 3160 7546 3188 7822
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3344 7546 3372 7686
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1780 7002 1808 7346
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 2916 7100 3224 7109
rect 2916 7098 2922 7100
rect 2978 7098 3002 7100
rect 3058 7098 3082 7100
rect 3138 7098 3162 7100
rect 3218 7098 3224 7100
rect 2978 7046 2980 7098
rect 3160 7046 3162 7098
rect 2916 7044 2922 7046
rect 2978 7044 3002 7046
rect 3058 7044 3082 7046
rect 3138 7044 3162 7046
rect 3218 7044 3224 7046
rect 2916 7035 3224 7044
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6458 3096 6666
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 940 6112 992 6118
rect 938 6080 940 6089
rect 992 6080 994 6089
rect 938 6015 994 6024
rect 2916 6012 3224 6021
rect 2916 6010 2922 6012
rect 2978 6010 3002 6012
rect 3058 6010 3082 6012
rect 3138 6010 3162 6012
rect 3218 6010 3224 6012
rect 2978 5958 2980 6010
rect 3160 5958 3162 6010
rect 2916 5956 2922 5958
rect 2978 5956 3002 5958
rect 3058 5956 3082 5958
rect 3138 5956 3162 5958
rect 3218 5956 3224 5958
rect 2916 5947 3224 5956
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 2916 4924 3224 4933
rect 2916 4922 2922 4924
rect 2978 4922 3002 4924
rect 3058 4922 3082 4924
rect 3138 4922 3162 4924
rect 3218 4922 3224 4924
rect 2978 4870 2980 4922
rect 3160 4870 3162 4922
rect 2916 4868 2922 4870
rect 2978 4868 3002 4870
rect 3058 4868 3082 4870
rect 3138 4868 3162 4870
rect 3218 4868 3224 4870
rect 2916 4859 3224 4868
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4457 980 4490
rect 938 4448 994 4457
rect 938 4383 994 4392
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 3641 980 3878
rect 2916 3836 3224 3845
rect 2916 3834 2922 3836
rect 2978 3834 3002 3836
rect 3058 3834 3082 3836
rect 3138 3834 3162 3836
rect 3218 3834 3224 3836
rect 2978 3782 2980 3834
rect 3160 3782 3162 3834
rect 2916 3780 2922 3782
rect 2978 3780 3002 3782
rect 3058 3780 3082 3782
rect 3138 3780 3162 3782
rect 3218 3780 3224 3782
rect 2916 3771 3224 3780
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 3252 3194 3280 7278
rect 3712 6866 3740 14758
rect 4540 12986 4568 15302
rect 4882 15260 5190 15269
rect 4882 15258 4888 15260
rect 4944 15258 4968 15260
rect 5024 15258 5048 15260
rect 5104 15258 5128 15260
rect 5184 15258 5190 15260
rect 4944 15206 4946 15258
rect 5126 15206 5128 15258
rect 4882 15204 4888 15206
rect 4944 15204 4968 15206
rect 5024 15204 5048 15206
rect 5104 15204 5128 15206
rect 5184 15204 5190 15206
rect 4882 15195 5190 15204
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5736 14482 5764 14962
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 4882 14172 5190 14181
rect 4882 14170 4888 14172
rect 4944 14170 4968 14172
rect 5024 14170 5048 14172
rect 5104 14170 5128 14172
rect 5184 14170 5190 14172
rect 4944 14118 4946 14170
rect 5126 14118 5128 14170
rect 4882 14116 4888 14118
rect 4944 14116 4968 14118
rect 5024 14116 5048 14118
rect 5104 14116 5128 14118
rect 5184 14116 5190 14118
rect 4882 14107 5190 14116
rect 4882 13084 5190 13093
rect 4882 13082 4888 13084
rect 4944 13082 4968 13084
rect 5024 13082 5048 13084
rect 5104 13082 5128 13084
rect 5184 13082 5190 13084
rect 4944 13030 4946 13082
rect 5126 13030 5128 13082
rect 4882 13028 4888 13030
rect 4944 13028 4968 13030
rect 5024 13028 5048 13030
rect 5104 13028 5128 13030
rect 5184 13028 5190 13030
rect 4882 13019 5190 13028
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4540 12238 4568 12922
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5368 12434 5396 12854
rect 5368 12406 5488 12434
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4882 11996 5190 12005
rect 4882 11994 4888 11996
rect 4944 11994 4968 11996
rect 5024 11994 5048 11996
rect 5104 11994 5128 11996
rect 5184 11994 5190 11996
rect 4944 11942 4946 11994
rect 5126 11942 5128 11994
rect 4882 11940 4888 11942
rect 4944 11940 4968 11942
rect 5024 11940 5048 11942
rect 5104 11940 5128 11942
rect 5184 11940 5190 11942
rect 4882 11931 5190 11940
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10810 4752 11086
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10810 4844 10950
rect 4882 10908 5190 10917
rect 4882 10906 4888 10908
rect 4944 10906 4968 10908
rect 5024 10906 5048 10908
rect 5104 10906 5128 10908
rect 5184 10906 5190 10908
rect 4944 10854 4946 10906
rect 5126 10854 5128 10906
rect 4882 10852 4888 10854
rect 4944 10852 4968 10854
rect 5024 10852 5048 10854
rect 5104 10852 5128 10854
rect 5184 10852 5190 10854
rect 4882 10843 5190 10852
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9654 4476 9862
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3804 8498 3832 9114
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8634 4200 8774
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3804 7886 3832 8434
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 7886 4200 8298
rect 4264 8090 4292 8366
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4540 7478 4568 10406
rect 4816 10130 4844 10746
rect 5460 10606 5488 12406
rect 5736 11762 5764 14418
rect 6196 14006 6224 15302
rect 7668 15162 7696 15302
rect 8815 15260 9123 15269
rect 8815 15258 8821 15260
rect 8877 15258 8901 15260
rect 8957 15258 8981 15260
rect 9037 15258 9061 15260
rect 9117 15258 9123 15260
rect 8877 15206 8879 15258
rect 9059 15206 9061 15258
rect 8815 15204 8821 15206
rect 8877 15204 8901 15206
rect 8957 15204 8981 15206
rect 9037 15204 9061 15206
rect 9117 15204 9123 15206
rect 8815 15195 9123 15204
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 6849 14716 7157 14725
rect 6849 14714 6855 14716
rect 6911 14714 6935 14716
rect 6991 14714 7015 14716
rect 7071 14714 7095 14716
rect 7151 14714 7157 14716
rect 6911 14662 6913 14714
rect 7093 14662 7095 14714
rect 6849 14660 6855 14662
rect 6911 14660 6935 14662
rect 6991 14660 7015 14662
rect 7071 14660 7095 14662
rect 7151 14660 7157 14662
rect 6849 14651 7157 14660
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6196 12850 6224 13942
rect 6849 13628 7157 13637
rect 6849 13626 6855 13628
rect 6911 13626 6935 13628
rect 6991 13626 7015 13628
rect 7071 13626 7095 13628
rect 7151 13626 7157 13628
rect 6911 13574 6913 13626
rect 7093 13574 7095 13626
rect 6849 13572 6855 13574
rect 6911 13572 6935 13574
rect 6991 13572 7015 13574
rect 7071 13572 7095 13574
rect 7151 13572 7157 13574
rect 6849 13563 7157 13572
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6849 12540 7157 12549
rect 6849 12538 6855 12540
rect 6911 12538 6935 12540
rect 6991 12538 7015 12540
rect 7071 12538 7095 12540
rect 7151 12538 7157 12540
rect 6911 12486 6913 12538
rect 7093 12486 7095 12538
rect 6849 12484 6855 12486
rect 6911 12484 6935 12486
rect 6991 12484 7015 12486
rect 7071 12484 7095 12486
rect 7151 12484 7157 12486
rect 6849 12475 7157 12484
rect 7576 12434 7604 14758
rect 7576 12406 7696 12434
rect 7668 12306 7696 12406
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11898 6960 12174
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7484 11830 7512 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11354 5672 11494
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 6012 10266 6040 10610
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 5816 10056 5868 10062
rect 6092 10056 6144 10062
rect 5868 10004 6040 10010
rect 5816 9998 6040 10004
rect 6092 9998 6144 10004
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 4724 9178 4752 9998
rect 5828 9982 6040 9998
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 4882 9820 5190 9829
rect 4882 9818 4888 9820
rect 4944 9818 4968 9820
rect 5024 9818 5048 9820
rect 5104 9818 5128 9820
rect 5184 9818 5190 9820
rect 4944 9766 4946 9818
rect 5126 9766 5128 9818
rect 4882 9764 4888 9766
rect 4944 9764 4968 9766
rect 5024 9764 5048 9766
rect 5104 9764 5128 9766
rect 5184 9764 5190 9766
rect 4882 9755 5190 9764
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9178 5028 9522
rect 5276 9518 5304 9862
rect 5736 9654 5764 9862
rect 5448 9648 5500 9654
rect 5446 9616 5448 9625
rect 5724 9648 5776 9654
rect 5500 9616 5502 9625
rect 5724 9590 5776 9596
rect 5446 9551 5502 9560
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4632 8974 4660 9114
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4882 8732 5190 8741
rect 4882 8730 4888 8732
rect 4944 8730 4968 8732
rect 5024 8730 5048 8732
rect 5104 8730 5128 8732
rect 5184 8730 5190 8732
rect 4944 8678 4946 8730
rect 5126 8678 5128 8730
rect 4882 8676 4888 8678
rect 4944 8676 4968 8678
rect 5024 8676 5048 8678
rect 5104 8676 5128 8678
rect 5184 8676 5190 8678
rect 4882 8667 5190 8676
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4632 7206 4660 7822
rect 4816 7546 4844 8366
rect 5000 8090 5028 8366
rect 5276 8090 5304 9454
rect 5356 8900 5408 8906
rect 5460 8888 5488 9551
rect 5828 9466 5856 9982
rect 6012 9926 6040 9982
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5736 9450 5856 9466
rect 5724 9444 5856 9450
rect 5776 9438 5856 9444
rect 5724 9386 5776 9392
rect 5408 8860 5488 8888
rect 5540 8900 5592 8906
rect 5356 8842 5408 8848
rect 5540 8842 5592 8848
rect 5552 8362 5580 8842
rect 5736 8634 5764 9386
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5828 8838 5856 9046
rect 5920 8974 5948 9862
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 8974 6040 9318
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 6104 8634 6132 9998
rect 6288 9722 6316 9998
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6288 8566 6316 8910
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5736 7818 5764 8230
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 4882 7644 5190 7653
rect 4882 7642 4888 7644
rect 4944 7642 4968 7644
rect 5024 7642 5048 7644
rect 5104 7642 5128 7644
rect 5184 7642 5190 7644
rect 4944 7590 4946 7642
rect 5126 7590 5128 7642
rect 4882 7588 4888 7590
rect 4944 7588 4968 7590
rect 5024 7588 5048 7590
rect 5104 7588 5128 7590
rect 5184 7588 5190 7590
rect 4882 7579 5190 7588
rect 5828 7546 5856 8298
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3344 6225 3372 6258
rect 4080 6254 4108 6598
rect 4068 6248 4120 6254
rect 3330 6216 3386 6225
rect 4068 6190 4120 6196
rect 3330 6151 3386 6160
rect 4264 5760 4292 6734
rect 4632 6458 4660 6802
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4264 5732 4384 5760
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5234 4200 5510
rect 4264 5370 4292 5578
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4356 5234 4384 5732
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4356 5030 4384 5170
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 4622 4384 4966
rect 4448 4826 4476 6190
rect 4632 5370 4660 6394
rect 4724 6118 4752 6734
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 6458 4844 6598
rect 4882 6556 5190 6565
rect 4882 6554 4888 6556
rect 4944 6554 4968 6556
rect 5024 6554 5048 6556
rect 5104 6554 5128 6556
rect 5184 6554 5190 6556
rect 4944 6502 4946 6554
rect 5126 6502 5128 6554
rect 4882 6500 4888 6502
rect 4944 6500 4968 6502
rect 5024 6500 5048 6502
rect 5104 6500 5128 6502
rect 5184 6500 5190 6502
rect 4882 6491 5190 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 5092 5914 5120 6326
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4882 5468 5190 5477
rect 4882 5466 4888 5468
rect 4944 5466 4968 5468
rect 5024 5466 5048 5468
rect 5104 5466 5128 5468
rect 5184 5466 5190 5468
rect 4944 5414 4946 5466
rect 5126 5414 5128 5466
rect 4882 5412 4888 5414
rect 4944 5412 4968 5414
rect 5024 5412 5048 5414
rect 5104 5412 5128 5414
rect 5184 5412 5190 5414
rect 4882 5403 5190 5412
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5234 5120 5306
rect 5276 5250 5304 7142
rect 5368 6780 5396 7346
rect 5460 6934 5488 7346
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5630 6896 5686 6905
rect 5630 6831 5632 6840
rect 5684 6831 5686 6840
rect 5632 6802 5684 6808
rect 5540 6792 5592 6798
rect 5368 6752 5540 6780
rect 5540 6734 5592 6740
rect 5552 5914 5580 6734
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6322 5948 6598
rect 6288 6322 6316 7142
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5448 5296 5500 5302
rect 5276 5244 5448 5250
rect 5276 5238 5500 5244
rect 5080 5228 5132 5234
rect 5276 5222 5488 5238
rect 5080 5170 5132 5176
rect 5736 5098 5764 5714
rect 6196 5574 6224 6258
rect 6380 6254 6408 10542
rect 6472 9586 6500 11630
rect 6849 11452 7157 11461
rect 6849 11450 6855 11452
rect 6911 11450 6935 11452
rect 6991 11450 7015 11452
rect 7071 11450 7095 11452
rect 7151 11450 7157 11452
rect 6911 11398 6913 11450
rect 7093 11398 7095 11450
rect 6849 11396 6855 11398
rect 6911 11396 6935 11398
rect 6991 11396 7015 11398
rect 7071 11396 7095 11398
rect 7151 11396 7157 11398
rect 6849 11387 7157 11396
rect 7392 11234 7420 11698
rect 7484 11354 7512 11766
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11354 7604 11698
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 6920 11212 6972 11218
rect 7392 11206 7512 11234
rect 6920 11154 6972 11160
rect 6932 10810 6960 11154
rect 7484 11150 7512 11206
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7024 10742 7052 10950
rect 7484 10810 7512 11086
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6644 10668 6696 10674
rect 6564 10628 6644 10656
rect 6564 10130 6592 10628
rect 6644 10610 6696 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6849 10364 7157 10373
rect 6849 10362 6855 10364
rect 6911 10362 6935 10364
rect 6991 10362 7015 10364
rect 7071 10362 7095 10364
rect 7151 10362 7157 10364
rect 6911 10310 6913 10362
rect 7093 10310 7095 10362
rect 6849 10308 6855 10310
rect 6911 10308 6935 10310
rect 6991 10308 7015 10310
rect 7071 10308 7095 10310
rect 7151 10308 7157 10310
rect 6849 10299 7157 10308
rect 6644 10192 6696 10198
rect 6828 10192 6880 10198
rect 6696 10140 6828 10146
rect 6644 10134 6880 10140
rect 6552 10124 6604 10130
rect 6656 10118 6868 10134
rect 6552 10066 6604 10072
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6472 8090 6500 9522
rect 6849 9276 7157 9285
rect 6849 9274 6855 9276
rect 6911 9274 6935 9276
rect 6991 9274 7015 9276
rect 7071 9274 7095 9276
rect 7151 9274 7157 9276
rect 6911 9222 6913 9274
rect 7093 9222 7095 9274
rect 6849 9220 6855 9222
rect 6911 9220 6935 9222
rect 6991 9220 7015 9222
rect 7071 9220 7095 9222
rect 7151 9220 7157 9222
rect 6849 9211 7157 9220
rect 7208 9178 7236 9522
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 8566 6868 9046
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6472 7410 6500 8026
rect 6748 7478 6776 8366
rect 6849 8188 7157 8197
rect 6849 8186 6855 8188
rect 6911 8186 6935 8188
rect 6991 8186 7015 8188
rect 7071 8186 7095 8188
rect 7151 8186 7157 8188
rect 6911 8134 6913 8186
rect 7093 8134 7095 8186
rect 6849 8132 6855 8134
rect 6911 8132 6935 8134
rect 6991 8132 7015 8134
rect 7071 8132 7095 8134
rect 7151 8132 7157 8134
rect 6849 8123 7157 8132
rect 7208 7970 7236 8910
rect 7300 8090 7328 9658
rect 7392 9110 7420 10406
rect 8128 10130 8156 14894
rect 9232 14414 9260 15302
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8815 14172 9123 14181
rect 8815 14170 8821 14172
rect 8877 14170 8901 14172
rect 8957 14170 8981 14172
rect 9037 14170 9061 14172
rect 9117 14170 9123 14172
rect 8877 14118 8879 14170
rect 9059 14118 9061 14170
rect 8815 14116 8821 14118
rect 8877 14116 8901 14118
rect 8957 14116 8981 14118
rect 9037 14116 9061 14118
rect 9117 14116 9123 14118
rect 8815 14107 9123 14116
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9048 13530 9076 13874
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9324 13326 9352 14010
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9692 13326 9720 13670
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12986 8524 13194
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8815 13084 9123 13093
rect 8815 13082 8821 13084
rect 8877 13082 8901 13084
rect 8957 13082 8981 13084
rect 9037 13082 9061 13084
rect 9117 13082 9123 13084
rect 8877 13030 8879 13082
rect 9059 13030 9061 13082
rect 8815 13028 8821 13030
rect 8877 13028 8901 13030
rect 8957 13028 8981 13030
rect 9037 13028 9061 13030
rect 9117 13028 9123 13030
rect 8815 13019 9123 13028
rect 9232 12986 9260 13126
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 10810 8248 11494
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9586 7604 9862
rect 8312 9654 8340 11018
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9178 7972 9454
rect 8404 9382 8432 9998
rect 8496 9602 8524 12718
rect 9324 12442 9352 13262
rect 9692 12986 9720 13262
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9876 12850 9904 13126
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9692 12238 9720 12786
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 8815 11996 9123 12005
rect 8815 11994 8821 11996
rect 8877 11994 8901 11996
rect 8957 11994 8981 11996
rect 9037 11994 9061 11996
rect 9117 11994 9123 11996
rect 8877 11942 8879 11994
rect 9059 11942 9061 11994
rect 8815 11940 8821 11942
rect 8877 11940 8901 11942
rect 8957 11940 8981 11942
rect 9037 11940 9061 11942
rect 9117 11940 9123 11942
rect 8815 11931 9123 11940
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9048 11354 9076 11766
rect 9140 11354 9168 11834
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9968 11234 9996 14962
rect 10612 14618 10640 15302
rect 11624 15162 11652 15506
rect 12084 15502 12112 17200
rect 13648 15570 13676 17200
rect 14715 15804 15023 15813
rect 14715 15802 14721 15804
rect 14777 15802 14801 15804
rect 14857 15802 14881 15804
rect 14937 15802 14961 15804
rect 15017 15802 15023 15804
rect 14777 15750 14779 15802
rect 14959 15750 14961 15802
rect 14715 15748 14721 15750
rect 14777 15748 14801 15750
rect 14857 15748 14881 15750
rect 14937 15748 14961 15750
rect 15017 15748 15023 15750
rect 14715 15739 15023 15748
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 12072 15496 12124 15502
rect 15120 15450 15148 17462
rect 15198 17200 15254 18000
rect 16762 17200 16818 18000
rect 15212 15502 15240 17200
rect 16486 16688 16542 16697
rect 16486 16623 16542 16632
rect 12072 15438 12124 15444
rect 15028 15422 15148 15450
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15752 15428 15804 15434
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 12176 15094 12204 15302
rect 12748 15260 13056 15269
rect 12748 15258 12754 15260
rect 12810 15258 12834 15260
rect 12890 15258 12914 15260
rect 12970 15258 12994 15260
rect 13050 15258 13056 15260
rect 12810 15206 12812 15258
rect 12992 15206 12994 15258
rect 12748 15204 12754 15206
rect 12810 15204 12834 15206
rect 12890 15204 12914 15206
rect 12970 15204 12994 15206
rect 13050 15204 13056 15206
rect 12748 15195 13056 15204
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 10782 14716 11090 14725
rect 10782 14714 10788 14716
rect 10844 14714 10868 14716
rect 10924 14714 10948 14716
rect 11004 14714 11028 14716
rect 11084 14714 11090 14716
rect 10844 14662 10846 14714
rect 11026 14662 11028 14714
rect 10782 14660 10788 14662
rect 10844 14660 10868 14662
rect 10924 14660 10948 14662
rect 11004 14660 11028 14662
rect 11084 14660 11090 14662
rect 10782 14651 11090 14660
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 12176 14414 12204 15030
rect 13740 14414 13768 15302
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 12434 10088 14214
rect 10336 14074 10364 14350
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10520 14074 10548 14214
rect 10796 14074 10824 14214
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 11440 13870 11468 14282
rect 11532 13870 11560 14350
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10428 13394 10456 13670
rect 10704 13530 10732 13670
rect 10782 13628 11090 13637
rect 10782 13626 10788 13628
rect 10844 13626 10868 13628
rect 10924 13626 10948 13628
rect 11004 13626 11028 13628
rect 11084 13626 11090 13628
rect 10844 13574 10846 13626
rect 11026 13574 11028 13626
rect 10782 13572 10788 13574
rect 10844 13572 10868 13574
rect 10924 13572 10948 13574
rect 11004 13572 11028 13574
rect 11084 13572 11090 13574
rect 10782 13563 11090 13572
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 11532 12714 11560 13806
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11900 12986 11928 13194
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12176 12918 12204 13670
rect 12268 13258 12296 13670
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 10782 12540 11090 12549
rect 10782 12538 10788 12540
rect 10844 12538 10868 12540
rect 10924 12538 10948 12540
rect 11004 12538 11028 12540
rect 11084 12538 11090 12540
rect 10844 12486 10846 12538
rect 11026 12486 11028 12538
rect 10782 12484 10788 12486
rect 10844 12484 10868 12486
rect 10924 12484 10948 12486
rect 11004 12484 11028 12486
rect 11084 12484 11090 12486
rect 10782 12475 11090 12484
rect 10060 12406 10272 12434
rect 10244 11694 10272 12406
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11898 10364 12106
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10520 11898 10548 12038
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9968 11206 10088 11234
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 8815 10908 9123 10917
rect 8815 10906 8821 10908
rect 8877 10906 8901 10908
rect 8957 10906 8981 10908
rect 9037 10906 9061 10908
rect 9117 10906 9123 10908
rect 8877 10854 8879 10906
rect 9059 10854 9061 10906
rect 8815 10852 8821 10854
rect 8877 10852 8901 10854
rect 8957 10852 8981 10854
rect 9037 10852 9061 10854
rect 9117 10852 9123 10854
rect 8815 10843 9123 10852
rect 9232 10690 9260 10950
rect 9140 10674 9260 10690
rect 9692 10674 9720 11018
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9128 10668 9260 10674
rect 9180 10662 9260 10668
rect 9312 10668 9364 10674
rect 9128 10610 9180 10616
rect 9312 10610 9364 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 8956 10266 8984 10610
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9140 9994 9168 10610
rect 9324 10266 9352 10610
rect 9508 10470 9536 10610
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9876 10198 9904 10542
rect 9968 10470 9996 11018
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 9722 8616 9862
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8680 9654 8708 9930
rect 8815 9820 9123 9829
rect 8815 9818 8821 9820
rect 8877 9818 8901 9820
rect 8957 9818 8981 9820
rect 9037 9818 9061 9820
rect 9117 9818 9123 9820
rect 8877 9766 8879 9818
rect 9059 9766 9061 9818
rect 8815 9764 8821 9766
rect 8877 9764 8901 9766
rect 8957 9764 8981 9766
rect 9037 9764 9061 9766
rect 9117 9764 9123 9766
rect 8815 9755 9123 9764
rect 8668 9648 8720 9654
rect 8496 9574 8616 9602
rect 8668 9590 8720 9596
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 8496 8974 8524 9318
rect 8588 8974 8616 9574
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 9310 9072 9366 9081
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8496 8634 8524 8910
rect 8588 8634 8616 8910
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7208 7942 7328 7970
rect 7300 7886 7328 7942
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6656 7002 6684 7346
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6748 6882 6776 7414
rect 6849 7100 7157 7109
rect 6849 7098 6855 7100
rect 6911 7098 6935 7100
rect 6991 7098 7015 7100
rect 7071 7098 7095 7100
rect 7151 7098 7157 7100
rect 6911 7046 6913 7098
rect 7093 7046 7095 7098
rect 6849 7044 6855 7046
rect 6911 7044 6935 7046
rect 6991 7044 7015 7046
rect 7071 7044 7095 7046
rect 7151 7044 7157 7046
rect 6849 7035 7157 7044
rect 6656 6854 6776 6882
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6361 6500 6734
rect 6458 6352 6514 6361
rect 6458 6287 6514 6296
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6380 5114 6408 6190
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 6288 5086 6408 5114
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4282 4200 4422
rect 4356 4282 4384 4558
rect 4816 4282 4844 4558
rect 5552 4554 5580 4966
rect 5736 4758 5764 5034
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 4882 4380 5190 4389
rect 4882 4378 4888 4380
rect 4944 4378 4968 4380
rect 5024 4378 5048 4380
rect 5104 4378 5128 4380
rect 5184 4378 5190 4380
rect 4944 4326 4946 4378
rect 5126 4326 5128 4378
rect 4882 4324 4888 4326
rect 4944 4324 4968 4326
rect 5024 4324 5048 4326
rect 5104 4324 5128 4326
rect 5184 4324 5190 4326
rect 4882 4315 5190 4324
rect 5276 4282 5304 4490
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3804 3738 3832 4150
rect 6288 4146 6316 5086
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4826 6408 4966
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6380 4282 6408 4558
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 4080 3602 4108 4014
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2596 2984 2648 2990
rect 2884 2938 2912 2994
rect 2596 2926 2648 2932
rect 940 2848 992 2854
rect 938 2816 940 2825
rect 992 2816 994 2825
rect 938 2751 994 2760
rect 2608 2582 2636 2926
rect 2792 2910 2912 2938
rect 2792 2650 2820 2910
rect 2916 2748 3224 2757
rect 2916 2746 2922 2748
rect 2978 2746 3002 2748
rect 3058 2746 3082 2748
rect 3138 2746 3162 2748
rect 3218 2746 3224 2748
rect 2978 2694 2980 2746
rect 3160 2694 3162 2746
rect 2916 2692 2922 2694
rect 2978 2692 3002 2694
rect 3058 2692 3082 2694
rect 3138 2692 3162 2694
rect 3218 2692 3224 2694
rect 2916 2683 3224 2692
rect 4080 2650 4108 3538
rect 4882 3292 5190 3301
rect 4882 3290 4888 3292
rect 4944 3290 4968 3292
rect 5024 3290 5048 3292
rect 5104 3290 5128 3292
rect 5184 3290 5190 3292
rect 4944 3238 4946 3290
rect 5126 3238 5128 3290
rect 4882 3236 4888 3238
rect 4944 3236 4968 3238
rect 5024 3236 5048 3238
rect 5104 3236 5128 3238
rect 5184 3236 5190 3238
rect 4882 3227 5190 3236
rect 5552 2650 5580 4082
rect 6380 3534 6408 4218
rect 6564 4010 6592 5102
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 6656 2514 6684 6854
rect 6849 6012 7157 6021
rect 6849 6010 6855 6012
rect 6911 6010 6935 6012
rect 6991 6010 7015 6012
rect 7071 6010 7095 6012
rect 7151 6010 7157 6012
rect 6911 5958 6913 6010
rect 7093 5958 7095 6010
rect 6849 5956 6855 5958
rect 6911 5956 6935 5958
rect 6991 5956 7015 5958
rect 7071 5956 7095 5958
rect 7151 5956 7157 5958
rect 6849 5947 7157 5956
rect 7208 5778 7236 7754
rect 7300 7546 7328 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7300 5710 7328 6734
rect 7392 6458 7420 8298
rect 7668 8294 7696 8366
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 8090 7696 8230
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8680 7886 8708 9046
rect 9310 9007 9366 9016
rect 9324 8974 9352 9007
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8815 8732 9123 8741
rect 8815 8730 8821 8732
rect 8877 8730 8901 8732
rect 8957 8730 8981 8732
rect 9037 8730 9061 8732
rect 9117 8730 9123 8732
rect 8877 8678 8879 8730
rect 9059 8678 9061 8730
rect 8815 8676 8821 8678
rect 8877 8676 8901 8678
rect 8957 8676 8981 8678
rect 9037 8676 9061 8678
rect 9117 8676 9123 8678
rect 8815 8667 9123 8676
rect 9600 8498 9628 9318
rect 9692 8634 9720 9998
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9784 8498 9812 9862
rect 9876 9586 9904 10134
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8634 9904 9318
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 8022 9444 8230
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8128 7546 8156 7822
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6458 7788 6734
rect 7852 6730 7880 7142
rect 8128 7002 8156 7482
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 6458 7880 6666
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7838 5808 7894 5817
rect 7838 5743 7840 5752
rect 7892 5743 7894 5752
rect 7840 5714 7892 5720
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7838 5672 7894 5681
rect 6920 5636 6972 5642
rect 7838 5607 7894 5616
rect 6920 5578 6972 5584
rect 6932 5302 6960 5578
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 4146 6776 5102
rect 6849 4924 7157 4933
rect 6849 4922 6855 4924
rect 6911 4922 6935 4924
rect 6991 4922 7015 4924
rect 7071 4922 7095 4924
rect 7151 4922 7157 4924
rect 6911 4870 6913 4922
rect 7093 4870 7095 4922
rect 6849 4868 6855 4870
rect 6911 4868 6935 4870
rect 6991 4868 7015 4870
rect 7071 4868 7095 4870
rect 7151 4868 7157 4870
rect 6849 4859 7157 4868
rect 7208 4706 7236 5510
rect 7378 5264 7434 5273
rect 7378 5199 7380 5208
rect 7432 5199 7434 5208
rect 7380 5170 7432 5176
rect 7116 4678 7236 4706
rect 7116 4622 7144 4678
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7852 4282 7880 5607
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3942 7512 4082
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 6849 3836 7157 3845
rect 6849 3834 6855 3836
rect 6911 3834 6935 3836
rect 6991 3834 7015 3836
rect 7071 3834 7095 3836
rect 7151 3834 7157 3836
rect 6911 3782 6913 3834
rect 7093 3782 7095 3834
rect 6849 3780 6855 3782
rect 6911 3780 6935 3782
rect 6991 3780 7015 3782
rect 7071 3780 7095 3782
rect 7151 3780 7157 3782
rect 6849 3771 7157 3780
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 6932 3194 6960 3402
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3194 7052 3334
rect 7484 3194 7512 3402
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7944 3126 7972 6734
rect 8022 6216 8078 6225
rect 8220 6186 8248 6734
rect 8022 6151 8078 6160
rect 8208 6180 8260 6186
rect 8036 5778 8064 6151
rect 8208 6122 8260 6128
rect 8312 5914 8340 7278
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 6458 8432 7142
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 6322 8524 7278
rect 8588 6322 8616 7686
rect 8680 7546 8708 7822
rect 8815 7644 9123 7653
rect 8815 7642 8821 7644
rect 8877 7642 8901 7644
rect 8957 7642 8981 7644
rect 9037 7642 9061 7644
rect 9117 7642 9123 7644
rect 8877 7590 8879 7642
rect 9059 7590 9061 7642
rect 8815 7588 8821 7590
rect 8877 7588 8901 7590
rect 8957 7588 8981 7590
rect 9037 7588 9061 7590
rect 9117 7588 9123 7590
rect 8815 7579 9123 7588
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 9128 7404 9180 7410
rect 9180 7364 9260 7392
rect 9128 7346 9180 7352
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8036 5234 8064 5714
rect 8208 5704 8260 5710
rect 8496 5658 8524 6258
rect 8680 6118 8708 6870
rect 8815 6556 9123 6565
rect 8815 6554 8821 6556
rect 8877 6554 8901 6556
rect 8957 6554 8981 6556
rect 9037 6554 9061 6556
rect 9117 6554 9123 6556
rect 8877 6502 8879 6554
rect 9059 6502 9061 6554
rect 8815 6500 8821 6502
rect 8877 6500 8901 6502
rect 8957 6500 8981 6502
rect 9037 6500 9061 6502
rect 9117 6500 9123 6502
rect 8815 6491 9123 6500
rect 8758 6352 8814 6361
rect 9232 6322 9260 7364
rect 8758 6287 8760 6296
rect 8812 6287 8814 6296
rect 9220 6316 9272 6322
rect 8760 6258 8812 6264
rect 9220 6258 9272 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8260 5652 8340 5658
rect 8208 5646 8340 5652
rect 8220 5630 8340 5646
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4146 8064 4626
rect 8312 4622 8340 5630
rect 8404 5630 8524 5658
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8312 3670 8340 4014
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3194 8156 3470
rect 8404 3194 8432 5630
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5370 8524 5510
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8588 5114 8616 6054
rect 8944 5840 8996 5846
rect 8666 5808 8722 5817
rect 8944 5782 8996 5788
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 8666 5743 8668 5752
rect 8720 5743 8722 5752
rect 8668 5714 8720 5720
rect 8956 5681 8984 5782
rect 9140 5710 9168 5782
rect 9128 5704 9180 5710
rect 8942 5672 8998 5681
rect 9128 5646 9180 5652
rect 8942 5607 8998 5616
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5166 8708 5510
rect 8815 5468 9123 5477
rect 8815 5466 8821 5468
rect 8877 5466 8901 5468
rect 8957 5466 8981 5468
rect 9037 5466 9061 5468
rect 9117 5466 9123 5468
rect 8877 5414 8879 5466
rect 9059 5414 9061 5466
rect 8815 5412 8821 5414
rect 8877 5412 8901 5414
rect 8957 5412 8981 5414
rect 9037 5412 9061 5414
rect 9117 5412 9123 5414
rect 8815 5403 9123 5412
rect 8944 5296 8996 5302
rect 8942 5264 8944 5273
rect 8996 5264 8998 5273
rect 8760 5228 8812 5234
rect 8942 5199 8998 5208
rect 8760 5170 8812 5176
rect 8496 5098 8616 5114
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8484 5092 8616 5098
rect 8536 5086 8616 5092
rect 8484 5034 8536 5040
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4282 8616 4966
rect 8668 4480 8720 4486
rect 8772 4468 8800 5170
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4826 8892 4966
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 9140 4570 9168 5034
rect 9232 4826 9260 6258
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9324 5234 9352 5782
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9140 4542 9260 4570
rect 8720 4440 8800 4468
rect 8668 4422 8720 4428
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8680 3534 8708 4422
rect 8815 4380 9123 4389
rect 8815 4378 8821 4380
rect 8877 4378 8901 4380
rect 8957 4378 8981 4380
rect 9037 4378 9061 4380
rect 9117 4378 9123 4380
rect 8877 4326 8879 4378
rect 9059 4326 9061 4378
rect 8815 4324 8821 4326
rect 8877 4324 8901 4326
rect 8957 4324 8981 4326
rect 9037 4324 9061 4326
rect 9117 4324 9123 4326
rect 8815 4315 9123 4324
rect 9232 4078 9260 4542
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8815 3292 9123 3301
rect 8815 3290 8821 3292
rect 8877 3290 8901 3292
rect 8957 3290 8981 3292
rect 9037 3290 9061 3292
rect 9117 3290 9123 3292
rect 8877 3238 8879 3290
rect 9059 3238 9061 3290
rect 8815 3236 8821 3238
rect 8877 3236 8901 3238
rect 8957 3236 8981 3238
rect 9037 3236 9061 3238
rect 9117 3236 9123 3238
rect 8815 3227 9123 3236
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 6849 2748 7157 2757
rect 6849 2746 6855 2748
rect 6911 2746 6935 2748
rect 6991 2746 7015 2748
rect 7071 2746 7095 2748
rect 7151 2746 7157 2748
rect 6911 2694 6913 2746
rect 7093 2694 7095 2746
rect 6849 2692 6855 2694
rect 6911 2692 6935 2694
rect 6991 2692 7015 2694
rect 7071 2692 7095 2694
rect 7151 2692 7157 2694
rect 6849 2683 7157 2692
rect 7576 2650 7604 2994
rect 9324 2650 9352 4422
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9416 2553 9444 7958
rect 9600 7018 9628 8434
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 7206 9720 8366
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9600 6990 9720 7018
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 3942 9536 5578
rect 9600 5234 9628 6802
rect 9692 5234 9720 6990
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6118 9812 6598
rect 10060 6338 10088 11206
rect 10152 11082 10180 11630
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10244 8430 10272 11630
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11354 10456 11494
rect 10782 11452 11090 11461
rect 10782 11450 10788 11452
rect 10844 11450 10868 11452
rect 10924 11450 10948 11452
rect 11004 11450 11028 11452
rect 11084 11450 11090 11452
rect 10844 11398 10846 11450
rect 11026 11398 11028 11450
rect 10782 11396 10788 11398
rect 10844 11396 10868 11398
rect 10924 11396 10948 11398
rect 11004 11396 11028 11398
rect 11084 11396 11090 11398
rect 10782 11387 11090 11396
rect 11348 11354 11376 12038
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11532 11121 11560 11630
rect 11518 11112 11574 11121
rect 10692 11076 10744 11082
rect 11518 11047 11574 11056
rect 10692 11018 10744 11024
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10428 9178 10456 9930
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10336 7002 10364 7754
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9968 6310 10088 6338
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9600 3738 9628 4490
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9784 2650 9812 6054
rect 9876 5370 9904 6258
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9968 4078 9996 6310
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5710 10088 6054
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10336 5234 10364 5782
rect 10428 5710 10456 9114
rect 10704 8838 10732 11018
rect 10782 10364 11090 10373
rect 10782 10362 10788 10364
rect 10844 10362 10868 10364
rect 10924 10362 10948 10364
rect 11004 10362 11028 10364
rect 11084 10362 11090 10364
rect 10844 10310 10846 10362
rect 11026 10310 11028 10362
rect 10782 10308 10788 10310
rect 10844 10308 10868 10310
rect 10924 10308 10948 10310
rect 11004 10308 11028 10310
rect 11084 10308 11090 10310
rect 10782 10299 11090 10308
rect 10782 9276 11090 9285
rect 10782 9274 10788 9276
rect 10844 9274 10868 9276
rect 10924 9274 10948 9276
rect 11004 9274 11028 9276
rect 11084 9274 11090 9276
rect 10844 9222 10846 9274
rect 11026 9222 11028 9274
rect 10782 9220 10788 9222
rect 10844 9220 10868 9222
rect 10924 9220 10948 9222
rect 11004 9220 11028 9222
rect 11084 9220 11090 9222
rect 10782 9211 11090 9220
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 11532 8634 11560 8910
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 10782 8188 11090 8197
rect 10782 8186 10788 8188
rect 10844 8186 10868 8188
rect 10924 8186 10948 8188
rect 11004 8186 11028 8188
rect 11084 8186 11090 8188
rect 10844 8134 10846 8186
rect 11026 8134 11028 8186
rect 10782 8132 10788 8134
rect 10844 8132 10868 8134
rect 10924 8132 10948 8134
rect 11004 8132 11028 8134
rect 11084 8132 11090 8134
rect 10782 8123 11090 8132
rect 11164 7818 11192 8230
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 10520 7478 10548 7754
rect 11164 7562 11192 7754
rect 11164 7534 11284 7562
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 6866 10548 7142
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10704 6458 10732 7278
rect 10782 7100 11090 7109
rect 10782 7098 10788 7100
rect 10844 7098 10868 7100
rect 10924 7098 10948 7100
rect 11004 7098 11028 7100
rect 11084 7098 11090 7100
rect 10844 7046 10846 7098
rect 11026 7046 11028 7098
rect 10782 7044 10788 7046
rect 10844 7044 10868 7046
rect 10924 7044 10948 7046
rect 11004 7044 11028 7046
rect 11084 7044 11090 7046
rect 10782 7035 11090 7044
rect 11164 7002 11192 7414
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4826 10456 5102
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3738 10364 3878
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10428 3466 10456 4762
rect 10612 4162 10640 5850
rect 10704 5370 10732 6394
rect 11072 6390 11100 6598
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11164 6118 11192 6666
rect 11256 6186 11284 7534
rect 11348 6866 11376 8298
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 6934 11468 7686
rect 11624 7002 11652 12174
rect 11992 11898 12020 12174
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11716 11354 11744 11630
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11992 11218 12020 11562
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10810 12112 11018
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10169 12020 10542
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 12268 10033 12296 10610
rect 12254 10024 12310 10033
rect 12254 9959 12310 9968
rect 12268 9926 12296 9959
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8634 12296 8910
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11716 7342 11744 8434
rect 12360 8412 12388 9318
rect 12452 9194 12480 14214
rect 12748 14172 13056 14181
rect 12748 14170 12754 14172
rect 12810 14170 12834 14172
rect 12890 14170 12914 14172
rect 12970 14170 12994 14172
rect 13050 14170 13056 14172
rect 12810 14118 12812 14170
rect 12992 14118 12994 14170
rect 12748 14116 12754 14118
rect 12810 14116 12834 14118
rect 12890 14116 12914 14118
rect 12970 14116 12994 14118
rect 13050 14116 13056 14118
rect 12748 14107 13056 14116
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12442 12572 13126
rect 12636 12850 12664 13670
rect 12728 13394 12756 13806
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13394 12848 13670
rect 13004 13530 13032 13874
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 13556 13190 13584 13670
rect 13648 13462 13676 14282
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 12748 13084 13056 13093
rect 12748 13082 12754 13084
rect 12810 13082 12834 13084
rect 12890 13082 12914 13084
rect 12970 13082 12994 13084
rect 13050 13082 13056 13084
rect 12810 13030 12812 13082
rect 12992 13030 12994 13082
rect 12748 13028 12754 13030
rect 12810 13028 12834 13030
rect 12890 13028 12914 13030
rect 12970 13028 12994 13030
rect 13050 13028 13056 13030
rect 12748 13019 13056 13028
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 13556 12782 13584 13126
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12544 11762 12572 12242
rect 12636 11880 12664 12582
rect 13004 12170 13032 12582
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12748 11996 13056 12005
rect 12748 11994 12754 11996
rect 12810 11994 12834 11996
rect 12890 11994 12914 11996
rect 12970 11994 12994 11996
rect 13050 11994 13056 11996
rect 12810 11942 12812 11994
rect 12992 11942 12994 11994
rect 12748 11940 12754 11942
rect 12810 11940 12834 11942
rect 12890 11940 12914 11942
rect 12970 11940 12994 11942
rect 13050 11940 13056 11942
rect 12748 11931 13056 11940
rect 12636 11852 12756 11880
rect 12728 11762 12756 11852
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12544 10266 12572 11698
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12748 10908 13056 10917
rect 12748 10906 12754 10908
rect 12810 10906 12834 10908
rect 12890 10906 12914 10908
rect 12970 10906 12994 10908
rect 13050 10906 13056 10908
rect 12810 10854 12812 10906
rect 12992 10854 12994 10906
rect 12748 10852 12754 10854
rect 12810 10852 12834 10854
rect 12890 10852 12914 10854
rect 12970 10852 12994 10854
rect 13050 10852 13056 10854
rect 12748 10843 13056 10852
rect 13096 10810 13124 11086
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13280 10674 13308 11630
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10674 13400 10950
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 13556 10062 13584 10474
rect 13648 10282 13676 12786
rect 13924 11286 13952 15098
rect 14752 15026 14780 15302
rect 15028 15026 15056 15422
rect 15752 15370 15804 15376
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13740 10606 13768 11018
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13648 10254 13768 10282
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13268 9988 13320 9994
rect 13320 9948 13492 9976
rect 13268 9930 13320 9936
rect 13464 9908 13492 9948
rect 13544 9920 13596 9926
rect 13464 9880 13544 9908
rect 13544 9862 13596 9868
rect 12748 9820 13056 9829
rect 12748 9818 12754 9820
rect 12810 9818 12834 9820
rect 12890 9818 12914 9820
rect 12970 9818 12994 9820
rect 13050 9818 13056 9820
rect 12810 9766 12812 9818
rect 12992 9766 12994 9818
rect 12748 9764 12754 9766
rect 12810 9764 12834 9766
rect 12890 9764 12914 9766
rect 12970 9764 12994 9766
rect 13050 9764 13056 9766
rect 12748 9755 13056 9764
rect 13084 9648 13136 9654
rect 13176 9648 13228 9654
rect 13084 9590 13136 9596
rect 13174 9616 13176 9625
rect 13228 9616 13230 9625
rect 12716 9376 12768 9382
rect 12636 9336 12716 9364
rect 12452 9178 12572 9194
rect 12452 9172 12584 9178
rect 12452 9166 12532 9172
rect 12532 9114 12584 9120
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12452 8566 12480 9046
rect 12636 8974 12664 9336
rect 12716 9318 12768 9324
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12440 8424 12492 8430
rect 12360 8384 12440 8412
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11440 6338 11468 6870
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11348 6310 11468 6338
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10782 6012 11090 6021
rect 10782 6010 10788 6012
rect 10844 6010 10868 6012
rect 10924 6010 10948 6012
rect 11004 6010 11028 6012
rect 11084 6010 11090 6012
rect 10844 5958 10846 6010
rect 11026 5958 11028 6010
rect 10782 5956 10788 5958
rect 10844 5956 10868 5958
rect 10924 5956 10948 5958
rect 11004 5956 11028 5958
rect 11084 5956 11090 5958
rect 10782 5947 11090 5956
rect 11348 5574 11376 6310
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11336 5568 11388 5574
rect 11242 5536 11298 5545
rect 11336 5510 11388 5516
rect 11242 5471 11298 5480
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 11256 5030 11284 5471
rect 11440 5098 11468 6190
rect 11532 5234 11560 6666
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11624 5914 11652 6394
rect 11808 5914 11836 8026
rect 11900 7818 11928 8230
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11900 6798 11928 7278
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10782 4924 11090 4933
rect 10782 4922 10788 4924
rect 10844 4922 10868 4924
rect 10924 4922 10948 4924
rect 11004 4922 11028 4924
rect 11084 4922 11090 4924
rect 10844 4870 10846 4922
rect 11026 4870 11028 4922
rect 10782 4868 10788 4870
rect 10844 4868 10868 4870
rect 10924 4868 10948 4870
rect 11004 4868 11028 4870
rect 11084 4868 11090 4870
rect 10782 4859 11090 4868
rect 10520 4134 10640 4162
rect 10784 4140 10836 4146
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10520 2774 10548 4134
rect 10784 4082 10836 4088
rect 10796 4026 10824 4082
rect 11256 4078 11284 4966
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11440 4214 11468 4422
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 10428 2746 10548 2774
rect 10612 3998 10824 4026
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9402 2544 9458 2553
rect 6644 2508 6696 2514
rect 9402 2479 9458 2488
rect 6644 2450 6696 2456
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6828 2440 6880 2446
rect 8300 2440 8352 2446
rect 6828 2382 6880 2388
rect 8220 2400 8300 2428
rect 860 800 888 2382
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2009 980 2314
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 2424 1306 2452 2382
rect 3896 1306 3924 2382
rect 4882 2204 5190 2213
rect 4882 2202 4888 2204
rect 4944 2202 4968 2204
rect 5024 2202 5048 2204
rect 5104 2202 5128 2204
rect 5184 2202 5190 2204
rect 4944 2150 4946 2202
rect 5126 2150 5128 2202
rect 4882 2148 4888 2150
rect 4944 2148 4968 2150
rect 5024 2148 5048 2150
rect 5104 2148 5128 2150
rect 5184 2148 5190 2150
rect 4882 2139 5190 2148
rect 5368 1306 5396 2382
rect 2332 1278 2452 1306
rect 3804 1278 3924 1306
rect 5276 1278 5396 1306
rect 2332 800 2360 1278
rect 3804 800 3832 1278
rect 5276 800 5304 1278
rect 6840 1034 6868 2382
rect 6748 1006 6868 1034
rect 6748 800 6776 1006
rect 8220 800 8248 2400
rect 8300 2382 8352 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10324 2440 10376 2446
rect 10428 2428 10456 2746
rect 10612 2446 10640 3998
rect 10796 3942 10824 3998
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10704 3738 10732 3878
rect 10782 3836 11090 3845
rect 10782 3834 10788 3836
rect 10844 3834 10868 3836
rect 10924 3834 10948 3836
rect 11004 3834 11028 3836
rect 11084 3834 11090 3836
rect 10844 3782 10846 3834
rect 11026 3782 11028 3834
rect 10782 3780 10788 3782
rect 10844 3780 10868 3782
rect 10924 3780 10948 3782
rect 11004 3780 11028 3782
rect 11084 3780 11090 3782
rect 10782 3771 11090 3780
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10704 3602 10732 3674
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 11440 3058 11468 4150
rect 11532 4146 11560 4966
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11716 4078 11744 5170
rect 11900 4468 11928 6054
rect 11992 5914 12020 6190
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12084 5778 12112 6666
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 5778 12204 6598
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12084 5302 12112 5714
rect 12268 5370 12296 7278
rect 12360 6866 12388 8384
rect 12440 8366 12492 8372
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7410 12480 8230
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12544 6662 12572 8434
rect 12636 8090 12664 8910
rect 12748 8732 13056 8741
rect 12748 8730 12754 8732
rect 12810 8730 12834 8732
rect 12890 8730 12914 8732
rect 12970 8730 12994 8732
rect 13050 8730 13056 8732
rect 12810 8678 12812 8730
rect 12992 8678 12994 8730
rect 12748 8676 12754 8678
rect 12810 8676 12834 8678
rect 12890 8676 12914 8678
rect 12970 8676 12994 8678
rect 13050 8676 13056 8678
rect 12748 8667 13056 8676
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12912 7886 12940 8434
rect 13096 8294 13124 9590
rect 13648 9586 13676 10066
rect 13174 9551 13230 9560
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13188 8362 13216 9114
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12900 7880 12952 7886
rect 12898 7848 12900 7857
rect 12952 7848 12954 7857
rect 13004 7818 13032 8026
rect 12898 7783 12954 7792
rect 12992 7812 13044 7818
rect 12992 7754 13044 7760
rect 12748 7644 13056 7653
rect 12748 7642 12754 7644
rect 12810 7642 12834 7644
rect 12890 7642 12914 7644
rect 12970 7642 12994 7644
rect 13050 7642 13056 7644
rect 12810 7590 12812 7642
rect 12992 7590 12994 7642
rect 12748 7588 12754 7590
rect 12810 7588 12834 7590
rect 12890 7588 12914 7590
rect 12970 7588 12994 7590
rect 13050 7588 13056 7590
rect 12748 7579 13056 7588
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12544 5234 12572 5782
rect 12636 5778 12664 6598
rect 12748 6556 13056 6565
rect 12748 6554 12754 6556
rect 12810 6554 12834 6556
rect 12890 6554 12914 6556
rect 12970 6554 12994 6556
rect 13050 6554 13056 6556
rect 12810 6502 12812 6554
rect 12992 6502 12994 6554
rect 12748 6500 12754 6502
rect 12810 6500 12834 6502
rect 12890 6500 12914 6502
rect 12970 6500 12994 6502
rect 13050 6500 13056 6502
rect 12748 6491 13056 6500
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12912 5778 12940 6122
rect 13004 5914 13032 6326
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12992 5704 13044 5710
rect 13096 5692 13124 8230
rect 13280 7970 13308 8570
rect 13372 8294 13400 9522
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9178 13584 9318
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13188 7942 13308 7970
rect 13188 7478 13216 7942
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13280 7546 13308 7754
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13280 7002 13308 7482
rect 13372 7002 13400 7754
rect 13556 7290 13584 8502
rect 13740 7818 13768 10254
rect 13832 10130 13860 10678
rect 13924 10470 13952 10950
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14016 8922 14044 14962
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14292 13462 14320 13670
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12434 14228 12718
rect 14292 12714 14320 13398
rect 14476 13190 14504 13670
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14384 12986 14412 13126
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14476 12866 14504 13126
rect 14384 12838 14504 12866
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14384 12442 14412 12838
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14108 12406 14228 12434
rect 14372 12436 14424 12442
rect 14108 12102 14136 12406
rect 14372 12378 14424 12384
rect 14384 12102 14412 12378
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14476 11830 14504 12582
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14568 11200 14596 14758
rect 14715 14716 15023 14725
rect 14715 14714 14721 14716
rect 14777 14714 14801 14716
rect 14857 14714 14881 14716
rect 14937 14714 14961 14716
rect 15017 14714 15023 14716
rect 14777 14662 14779 14714
rect 14959 14662 14961 14714
rect 14715 14660 14721 14662
rect 14777 14660 14801 14662
rect 14857 14660 14881 14662
rect 14937 14660 14961 14662
rect 15017 14660 15023 14662
rect 14715 14651 15023 14660
rect 15120 14618 15148 15302
rect 15580 15065 15608 15302
rect 15764 15162 15792 15370
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15566 15056 15622 15065
rect 15476 15020 15528 15026
rect 15672 15026 15700 15098
rect 15566 14991 15622 15000
rect 15660 15020 15712 15026
rect 15476 14962 15528 14968
rect 15660 14962 15712 14968
rect 15488 14906 15516 14962
rect 15948 14958 15976 15370
rect 16500 15162 16528 16623
rect 16670 15872 16726 15881
rect 16670 15807 16726 15816
rect 16684 15706 16712 15807
rect 16776 15706 16804 17200
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16681 15260 16989 15269
rect 16681 15258 16687 15260
rect 16743 15258 16767 15260
rect 16823 15258 16847 15260
rect 16903 15258 16927 15260
rect 16983 15258 16989 15260
rect 16743 15206 16745 15258
rect 16925 15206 16927 15258
rect 16681 15204 16687 15206
rect 16743 15204 16767 15206
rect 16823 15204 16847 15206
rect 16903 15204 16927 15206
rect 16983 15204 16989 15206
rect 16681 15195 16989 15204
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 15936 14952 15988 14958
rect 15488 14878 15884 14906
rect 15936 14894 15988 14900
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14618 15516 14758
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 14074 14780 14214
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 14715 13628 15023 13637
rect 14715 13626 14721 13628
rect 14777 13626 14801 13628
rect 14857 13626 14881 13628
rect 14937 13626 14961 13628
rect 15017 13626 15023 13628
rect 14777 13574 14779 13626
rect 14959 13574 14961 13626
rect 14715 13572 14721 13574
rect 14777 13572 14801 13574
rect 14857 13572 14881 13574
rect 14937 13572 14961 13574
rect 15017 13572 15023 13574
rect 14715 13563 15023 13572
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12986 14688 13262
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14715 12540 15023 12549
rect 14715 12538 14721 12540
rect 14777 12538 14801 12540
rect 14857 12538 14881 12540
rect 14937 12538 14961 12540
rect 15017 12538 15023 12540
rect 14777 12486 14779 12538
rect 14959 12486 14961 12538
rect 14715 12484 14721 12486
rect 14777 12484 14801 12486
rect 14857 12484 14881 12486
rect 14937 12484 14961 12486
rect 15017 12484 15023 12486
rect 14715 12475 15023 12484
rect 15120 11801 15148 13806
rect 15304 13394 15332 13874
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 15212 11558 15240 12718
rect 15396 11898 15424 14350
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15488 13326 15516 14214
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15580 12306 15608 14214
rect 15672 13530 15700 14350
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 14074 15792 14214
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 14715 11452 15023 11461
rect 14715 11450 14721 11452
rect 14777 11450 14801 11452
rect 14857 11450 14881 11452
rect 14937 11450 14961 11452
rect 15017 11450 15023 11452
rect 14777 11398 14779 11450
rect 14959 11398 14961 11450
rect 14715 11396 14721 11398
rect 14777 11396 14801 11398
rect 14857 11396 14881 11398
rect 14937 11396 14961 11398
rect 15017 11396 15023 11398
rect 14715 11387 15023 11396
rect 14292 11172 14596 11200
rect 14186 11112 14242 11121
rect 14186 11047 14188 11056
rect 14240 11047 14242 11056
rect 14188 11018 14240 11024
rect 14292 10146 14320 11172
rect 14554 11112 14610 11121
rect 15580 11082 15608 11494
rect 15672 11354 15700 12174
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 14554 11047 14556 11056
rect 14608 11047 14610 11056
rect 15568 11076 15620 11082
rect 14556 11018 14608 11024
rect 15568 11018 15620 11024
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10742 14412 10950
rect 15764 10742 15792 13806
rect 15856 12782 15884 14878
rect 16486 14376 16542 14385
rect 16486 14311 16488 14320
rect 16540 14311 16542 14320
rect 16488 14282 16540 14288
rect 16681 14172 16989 14181
rect 16681 14170 16687 14172
rect 16743 14170 16767 14172
rect 16823 14170 16847 14172
rect 16903 14170 16927 14172
rect 16983 14170 16989 14172
rect 16743 14118 16745 14170
rect 16925 14118 16927 14170
rect 16681 14116 16687 14118
rect 16743 14116 16767 14118
rect 16823 14116 16847 14118
rect 16903 14116 16927 14118
rect 16983 14116 16989 14118
rect 16681 14107 16989 14116
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 15844 12776 15896 12782
rect 15896 12736 15976 12764
rect 15844 12718 15896 12724
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15948 10606 15976 12736
rect 16132 11354 16160 12854
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16224 11218 16252 11698
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16316 10810 16344 12038
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 14832 10600 14884 10606
rect 14830 10568 14832 10577
rect 15936 10600 15988 10606
rect 14884 10568 14886 10577
rect 14372 10532 14424 10538
rect 15936 10542 15988 10548
rect 14830 10503 14886 10512
rect 14372 10474 14424 10480
rect 14384 10266 14412 10474
rect 14715 10364 15023 10373
rect 14715 10362 14721 10364
rect 14777 10362 14801 10364
rect 14857 10362 14881 10364
rect 14937 10362 14961 10364
rect 15017 10362 15023 10364
rect 14777 10310 14779 10362
rect 14959 10310 14961 10362
rect 14715 10308 14721 10310
rect 14777 10308 14801 10310
rect 14857 10308 14881 10310
rect 14937 10308 14961 10310
rect 15017 10308 15023 10310
rect 14715 10299 15023 10308
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 16302 10160 16358 10169
rect 14096 10124 14148 10130
rect 14292 10118 14412 10146
rect 14096 10066 14148 10072
rect 14108 9625 14136 10066
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 13924 8894 14044 8922
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8566 13860 8774
rect 13924 8634 13952 8894
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13924 8022 13952 8570
rect 14016 8498 14044 8774
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14108 8090 14136 8774
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 14200 7857 14228 8910
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7886 14320 8230
rect 14384 7970 14412 10118
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 15660 10124 15712 10130
rect 16302 10095 16358 10104
rect 15660 10066 15712 10072
rect 14476 8634 14504 10066
rect 14648 10056 14700 10062
rect 14646 10024 14648 10033
rect 15016 10056 15068 10062
rect 14700 10024 14702 10033
rect 15016 9998 15068 10004
rect 14646 9959 14702 9968
rect 15028 9722 15056 9998
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 14568 9042 14596 9522
rect 14715 9276 15023 9285
rect 14715 9274 14721 9276
rect 14777 9274 14801 9276
rect 14857 9274 14881 9276
rect 14937 9274 14961 9276
rect 15017 9274 15023 9276
rect 14777 9222 14779 9274
rect 14959 9222 14961 9274
rect 14715 9220 14721 9222
rect 14777 9220 14801 9222
rect 14857 9220 14881 9222
rect 14937 9220 14961 9222
rect 15017 9220 15023 9222
rect 14715 9211 15023 9220
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14476 8090 14504 8570
rect 14568 8498 14596 8978
rect 15212 8634 15240 9522
rect 15304 9110 15332 9930
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 9110 15516 9862
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15488 8634 15516 9046
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15106 8528 15162 8537
rect 14556 8492 14608 8498
rect 15106 8463 15162 8472
rect 14556 8434 14608 8440
rect 14715 8188 15023 8197
rect 14715 8186 14721 8188
rect 14777 8186 14801 8188
rect 14857 8186 14881 8188
rect 14937 8186 14961 8188
rect 15017 8186 15023 8188
rect 14777 8134 14779 8186
rect 14959 8134 14961 8186
rect 14715 8132 14721 8134
rect 14777 8132 14801 8134
rect 14857 8132 14881 8134
rect 14937 8132 14961 8134
rect 15017 8132 15023 8134
rect 14715 8123 15023 8132
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14384 7942 14596 7970
rect 14280 7880 14332 7886
rect 14186 7848 14242 7857
rect 13728 7812 13780 7818
rect 14280 7822 14332 7828
rect 14186 7783 14242 7792
rect 13728 7754 13780 7760
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13556 7262 13676 7290
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13556 6866 13584 7142
rect 13648 6866 13676 7262
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13740 6798 13768 7346
rect 14016 6798 14044 7686
rect 14096 7540 14148 7546
rect 14200 7528 14228 7783
rect 14148 7500 14228 7528
rect 14096 7482 14148 7488
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 6866 14136 7278
rect 14200 6934 14228 7346
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13280 5914 13308 6258
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13044 5664 13124 5692
rect 12992 5646 13044 5652
rect 12748 5468 13056 5477
rect 12748 5466 12754 5468
rect 12810 5466 12834 5468
rect 12890 5466 12914 5468
rect 12970 5466 12994 5468
rect 13050 5466 13056 5468
rect 12810 5414 12812 5466
rect 12992 5414 12994 5466
rect 12748 5412 12754 5414
rect 12810 5412 12834 5414
rect 12890 5412 12914 5414
rect 12970 5412 12994 5414
rect 13050 5412 13056 5414
rect 12748 5403 13056 5412
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12544 4622 12572 5170
rect 12532 4616 12584 4622
rect 12438 4584 12494 4593
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 12360 4542 12438 4570
rect 11808 4440 11928 4468
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11532 3194 11560 3538
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11336 2848 11388 2854
rect 11388 2796 11560 2802
rect 11336 2790 11560 2796
rect 11348 2774 11560 2790
rect 10782 2748 11090 2757
rect 10782 2746 10788 2748
rect 10844 2746 10868 2748
rect 10924 2746 10948 2748
rect 11004 2746 11028 2748
rect 11084 2746 11090 2748
rect 10844 2694 10846 2746
rect 11026 2694 11028 2746
rect 10782 2692 10788 2694
rect 10844 2692 10868 2694
rect 10924 2692 10948 2694
rect 11004 2692 11028 2694
rect 11084 2692 11090 2694
rect 10782 2683 11090 2692
rect 11426 2680 11482 2689
rect 11426 2615 11428 2624
rect 11480 2615 11482 2624
rect 11428 2586 11480 2592
rect 11532 2446 11560 2774
rect 11624 2650 11652 2926
rect 11716 2854 11744 3062
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 10376 2400 10456 2428
rect 10600 2440 10652 2446
rect 10324 2382 10376 2388
rect 10600 2382 10652 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 8815 2204 9123 2213
rect 8815 2202 8821 2204
rect 8877 2202 8901 2204
rect 8957 2202 8981 2204
rect 9037 2202 9061 2204
rect 9117 2202 9123 2204
rect 8877 2150 8879 2202
rect 9059 2150 9061 2202
rect 8815 2148 8821 2150
rect 8877 2148 8901 2150
rect 8957 2148 8981 2150
rect 9037 2148 9061 2150
rect 9117 2148 9123 2150
rect 8815 2139 9123 2148
rect 9600 1834 9628 2382
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 9692 800 9720 2382
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10704 1970 10732 2246
rect 10796 2106 10824 2246
rect 10980 2106 11008 2246
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 10692 1964 10744 1970
rect 10692 1906 10744 1912
rect 11164 800 11192 2314
rect 11440 2038 11468 2382
rect 11808 2310 11836 4440
rect 12084 4282 12112 4490
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12176 3534 12204 4082
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11900 3194 11928 3334
rect 12268 3194 12296 3334
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2650 12112 2926
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11886 2544 11942 2553
rect 11886 2479 11942 2488
rect 11900 2310 11928 2479
rect 12360 2446 12388 4542
rect 12532 4558 12584 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 12438 4519 12494 4528
rect 12748 4380 13056 4389
rect 12748 4378 12754 4380
rect 12810 4378 12834 4380
rect 12890 4378 12914 4380
rect 12970 4378 12994 4380
rect 13050 4378 13056 4380
rect 12810 4326 12812 4378
rect 12992 4326 12994 4378
rect 12748 4324 12754 4326
rect 12810 4324 12834 4326
rect 12890 4324 12914 4326
rect 12970 4324 12994 4326
rect 13050 4324 13056 4326
rect 12748 4315 13056 4324
rect 13096 4282 13124 4558
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13372 4146 13400 4422
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13004 3602 13032 4014
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3738 13308 3878
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12452 2530 12480 3402
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 3194 12664 3334
rect 12748 3292 13056 3301
rect 12748 3290 12754 3292
rect 12810 3290 12834 3292
rect 12890 3290 12914 3292
rect 12970 3290 12994 3292
rect 13050 3290 13056 3292
rect 12810 3238 12812 3290
rect 12992 3238 12994 3290
rect 12748 3236 12754 3238
rect 12810 3236 12834 3238
rect 12890 3236 12914 3238
rect 12970 3236 12994 3238
rect 13050 3236 13056 3238
rect 12748 3227 13056 3236
rect 13096 3194 13124 3470
rect 13464 3194 13492 6734
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 13648 6497 13676 6666
rect 13634 6488 13690 6497
rect 13634 6423 13690 6432
rect 14108 6322 14136 6666
rect 14292 6390 14320 7346
rect 14568 6882 14596 7942
rect 14715 7100 15023 7109
rect 14715 7098 14721 7100
rect 14777 7098 14801 7100
rect 14857 7098 14881 7100
rect 14937 7098 14961 7100
rect 15017 7098 15023 7100
rect 14777 7046 14779 7098
rect 14959 7046 14961 7098
rect 14715 7044 14721 7046
rect 14777 7044 14801 7046
rect 14857 7044 14881 7046
rect 14937 7044 14961 7046
rect 15017 7044 15023 7046
rect 14715 7035 15023 7044
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14740 6928 14792 6934
rect 14568 6876 14740 6882
rect 14568 6870 14792 6876
rect 14830 6896 14886 6905
rect 14372 6860 14424 6866
rect 14568 6854 14780 6870
rect 14830 6831 14832 6840
rect 14372 6802 14424 6808
rect 14884 6831 14886 6840
rect 14832 6802 14884 6808
rect 14384 6390 14412 6802
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14108 6202 14136 6258
rect 14372 6248 14424 6254
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13556 4622 13584 6054
rect 13740 5710 13768 6054
rect 13832 5914 13860 6122
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 14016 5710 14044 6190
rect 14108 6174 14320 6202
rect 14556 6248 14608 6254
rect 14372 6190 14424 6196
rect 14476 6208 14556 6236
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5370 13860 5578
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13818 5264 13874 5273
rect 13818 5199 13874 5208
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13740 4826 13768 5034
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13740 4706 13768 4762
rect 13648 4678 13768 4706
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13648 3534 13676 4678
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 4010 13768 4558
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13832 3890 13860 5199
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4758 14228 4966
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 4146 13952 4422
rect 14200 4146 14228 4694
rect 14292 4690 14320 6174
rect 14384 5574 14412 6190
rect 14476 5710 14504 6208
rect 14556 6190 14608 6196
rect 14660 6066 14688 6326
rect 14844 6225 14872 6394
rect 14830 6216 14886 6225
rect 14830 6151 14886 6160
rect 14936 6118 14964 6938
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15028 6730 15056 6870
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 14568 6038 14688 6066
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14292 4282 14320 4626
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14292 4146 14320 4218
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 13910 4040 13966 4049
rect 14292 4010 14320 4082
rect 13910 3975 13966 3984
rect 14280 4004 14332 4010
rect 13740 3862 13860 3890
rect 13740 3534 13768 3862
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13648 3194 13676 3470
rect 13924 3194 13952 3975
rect 14280 3946 14332 3952
rect 14476 3670 14504 5646
rect 14568 5370 14596 6038
rect 14715 6012 15023 6021
rect 14715 6010 14721 6012
rect 14777 6010 14801 6012
rect 14857 6010 14881 6012
rect 14937 6010 14961 6012
rect 15017 6010 15023 6012
rect 14777 5958 14779 6010
rect 14959 5958 14961 6010
rect 14715 5956 14721 5958
rect 14777 5956 14801 5958
rect 14857 5956 14881 5958
rect 14937 5956 14961 5958
rect 15017 5956 15023 5958
rect 14715 5947 15023 5956
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14568 4706 14596 5170
rect 14715 4924 15023 4933
rect 14715 4922 14721 4924
rect 14777 4922 14801 4924
rect 14857 4922 14881 4924
rect 14937 4922 14961 4924
rect 15017 4922 15023 4924
rect 14777 4870 14779 4922
rect 14959 4870 14961 4922
rect 14715 4868 14721 4870
rect 14777 4868 14801 4870
rect 14857 4868 14881 4870
rect 14937 4868 14961 4870
rect 15017 4868 15023 4870
rect 14715 4859 15023 4868
rect 14568 4690 14688 4706
rect 14568 4684 14700 4690
rect 14568 4678 14648 4684
rect 14648 4626 14700 4632
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4078 14596 4558
rect 14660 4214 14688 4626
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14936 4282 14964 4558
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14660 3890 14688 4014
rect 14568 3862 14688 3890
rect 14568 3738 14596 3862
rect 14715 3836 15023 3845
rect 14715 3834 14721 3836
rect 14777 3834 14801 3836
rect 14857 3834 14881 3836
rect 14937 3834 14961 3836
rect 15017 3834 15023 3836
rect 14777 3782 14779 3834
rect 14959 3782 14961 3834
rect 14715 3780 14721 3782
rect 14777 3780 14801 3782
rect 14857 3780 14881 3782
rect 14937 3780 14961 3782
rect 15017 3780 15023 3782
rect 14715 3771 15023 3780
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14464 3664 14516 3670
rect 14370 3632 14426 3641
rect 14292 3590 14370 3618
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12544 2650 12572 2926
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12452 2502 12664 2530
rect 12636 2446 12664 2502
rect 12912 2446 12940 3130
rect 14292 3058 14320 3590
rect 14464 3606 14516 3612
rect 14370 3567 14426 3576
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 3398 14596 3470
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3058 14872 3334
rect 15120 3176 15148 8463
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15212 5250 15240 7278
rect 15304 5914 15332 8366
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 6934 15424 7686
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15396 5710 15424 6666
rect 15488 6458 15516 8366
rect 15580 7818 15608 8774
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15672 7478 15700 10066
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16224 9761 16252 9930
rect 16210 9752 16266 9761
rect 16316 9722 16344 10095
rect 16210 9687 16266 9696
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9178 16160 9318
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16132 8906 16160 9114
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15764 7410 15792 8434
rect 16132 8362 16160 8842
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16224 7698 16252 8774
rect 16316 8634 16344 9522
rect 16408 8634 16436 13874
rect 16500 13433 16528 13874
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12594 16620 13262
rect 16681 13084 16989 13093
rect 16681 13082 16687 13084
rect 16743 13082 16767 13084
rect 16823 13082 16847 13084
rect 16903 13082 16927 13084
rect 16983 13082 16989 13084
rect 16743 13030 16745 13082
rect 16925 13030 16927 13082
rect 16681 13028 16687 13030
rect 16743 13028 16767 13030
rect 16823 13028 16847 13030
rect 16903 13028 16927 13030
rect 16983 13028 16989 13030
rect 16681 13019 16989 13028
rect 16762 12608 16818 12617
rect 16592 12566 16762 12594
rect 16762 12543 16818 12552
rect 16681 11996 16989 12005
rect 16681 11994 16687 11996
rect 16743 11994 16767 11996
rect 16823 11994 16847 11996
rect 16903 11994 16927 11996
rect 16983 11994 16989 11996
rect 16743 11942 16745 11994
rect 16925 11942 16927 11994
rect 16681 11940 16687 11942
rect 16743 11940 16767 11942
rect 16823 11940 16847 11942
rect 16903 11940 16927 11942
rect 16983 11940 16989 11942
rect 16681 11931 16989 11940
rect 16681 10908 16989 10917
rect 16681 10906 16687 10908
rect 16743 10906 16767 10908
rect 16823 10906 16847 10908
rect 16903 10906 16927 10908
rect 16983 10906 16989 10908
rect 16743 10854 16745 10906
rect 16925 10854 16927 10906
rect 16681 10852 16687 10854
rect 16743 10852 16767 10854
rect 16823 10852 16847 10854
rect 16903 10852 16927 10854
rect 16983 10852 16989 10854
rect 16681 10843 16989 10852
rect 16486 10160 16542 10169
rect 16486 10095 16542 10104
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8430 16528 10095
rect 16681 9820 16989 9829
rect 16681 9818 16687 9820
rect 16743 9818 16767 9820
rect 16823 9818 16847 9820
rect 16903 9818 16927 9820
rect 16983 9818 16989 9820
rect 16743 9766 16745 9818
rect 16925 9766 16927 9818
rect 16681 9764 16687 9766
rect 16743 9764 16767 9766
rect 16823 9764 16847 9766
rect 16903 9764 16927 9766
rect 16983 9764 16989 9766
rect 16681 9755 16989 9764
rect 16762 9344 16818 9353
rect 16762 9279 16818 9288
rect 16776 9178 16804 9279
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16681 8732 16989 8741
rect 16681 8730 16687 8732
rect 16743 8730 16767 8732
rect 16823 8730 16847 8732
rect 16903 8730 16927 8732
rect 16983 8730 16989 8732
rect 16743 8678 16745 8730
rect 16925 8678 16927 8730
rect 16681 8676 16687 8678
rect 16743 8676 16767 8678
rect 16823 8676 16847 8678
rect 16903 8676 16927 8678
rect 16983 8676 16989 8678
rect 16681 8667 16989 8676
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16224 7670 16344 7698
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 15580 6662 15608 7278
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15212 5222 15332 5250
rect 15488 5234 15516 5578
rect 15304 5166 15332 5222
rect 15476 5228 15528 5234
rect 15396 5188 15476 5216
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15212 4826 15240 5102
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15396 4706 15424 5188
rect 15476 5170 15528 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15304 4678 15424 4706
rect 15304 3194 15332 4678
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 3738 15424 4558
rect 15488 4282 15516 4966
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15580 4146 15608 6598
rect 15672 5846 15700 6598
rect 15750 6488 15806 6497
rect 15750 6423 15806 6432
rect 15844 6452 15896 6458
rect 15764 6322 15792 6423
rect 15844 6394 15896 6400
rect 15856 6361 15884 6394
rect 15842 6352 15898 6361
rect 15752 6316 15804 6322
rect 15842 6287 15898 6296
rect 15752 6258 15804 6264
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15672 3738 15700 5646
rect 15764 5234 15792 6258
rect 15842 6216 15898 6225
rect 15842 6151 15898 6160
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15764 4078 15792 4558
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15200 3188 15252 3194
rect 15120 3148 15200 3176
rect 15200 3130 15252 3136
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 13372 2650 13400 2994
rect 14016 2650 14044 2994
rect 14384 2650 14412 2994
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15658 2816 15714 2825
rect 14715 2748 15023 2757
rect 14715 2746 14721 2748
rect 14777 2746 14801 2748
rect 14857 2746 14881 2748
rect 14937 2746 14961 2748
rect 15017 2746 15023 2748
rect 14777 2694 14779 2746
rect 14959 2694 14961 2746
rect 14715 2692 14721 2694
rect 14777 2692 14801 2694
rect 14857 2692 14881 2694
rect 14937 2692 14961 2694
rect 15017 2692 15023 2694
rect 14715 2683 15023 2692
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 15120 2582 15148 2790
rect 15658 2751 15714 2760
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15672 2446 15700 2751
rect 15764 2650 15792 4014
rect 15856 3534 15884 6151
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15948 3194 15976 6734
rect 16040 4690 16068 7278
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6322 16160 7142
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16224 6254 16252 7278
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 5166 16160 5646
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16040 2650 16068 4014
rect 16132 3738 16160 5102
rect 16224 4146 16252 5782
rect 16316 5370 16344 7670
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16408 5234 16436 8298
rect 17224 7880 17276 7886
rect 16486 7848 16542 7857
rect 17224 7822 17276 7828
rect 16486 7783 16542 7792
rect 17132 7812 17184 7818
rect 16500 5370 16528 7783
rect 17132 7754 17184 7760
rect 16681 7644 16989 7653
rect 16681 7642 16687 7644
rect 16743 7642 16767 7644
rect 16823 7642 16847 7644
rect 16903 7642 16927 7644
rect 16983 7642 16989 7644
rect 16743 7590 16745 7642
rect 16925 7590 16927 7642
rect 16681 7588 16687 7590
rect 16743 7588 16767 7590
rect 16823 7588 16847 7590
rect 16903 7588 16927 7590
rect 16983 7588 16989 7590
rect 16681 7579 16989 7588
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16592 6458 16620 6831
rect 16681 6556 16989 6565
rect 16681 6554 16687 6556
rect 16743 6554 16767 6556
rect 16823 6554 16847 6556
rect 16903 6554 16927 6556
rect 16983 6554 16989 6556
rect 16743 6502 16745 6554
rect 16925 6502 16927 6554
rect 16681 6500 16687 6502
rect 16743 6500 16767 6502
rect 16823 6500 16847 6502
rect 16903 6500 16927 6502
rect 16983 6500 16989 6502
rect 16681 6491 16989 6500
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 17052 6390 17080 7482
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5642 16620 6190
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16592 5166 16620 5578
rect 16681 5468 16989 5477
rect 16681 5466 16687 5468
rect 16743 5466 16767 5468
rect 16823 5466 16847 5468
rect 16903 5466 16927 5468
rect 16983 5466 16989 5468
rect 16743 5414 16745 5466
rect 16925 5414 16927 5466
rect 16681 5412 16687 5414
rect 16743 5412 16767 5414
rect 16823 5412 16847 5414
rect 16903 5412 16927 5414
rect 16983 5412 16989 5414
rect 16681 5403 16989 5412
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16681 4380 16989 4389
rect 16681 4378 16687 4380
rect 16743 4378 16767 4380
rect 16823 4378 16847 4380
rect 16903 4378 16927 4380
rect 16983 4378 16989 4380
rect 16743 4326 16745 4378
rect 16925 4326 16927 4378
rect 16681 4324 16687 4326
rect 16743 4324 16767 4326
rect 16823 4324 16847 4326
rect 16903 4324 16927 4326
rect 16983 4324 16989 4326
rect 16681 4315 16989 4324
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16302 4040 16358 4049
rect 16302 3975 16358 3984
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16224 3058 16252 3878
rect 16316 3738 16344 3975
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 17144 3534 17172 7754
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16681 3292 16989 3301
rect 16681 3290 16687 3292
rect 16743 3290 16767 3292
rect 16823 3290 16847 3292
rect 16903 3290 16927 3292
rect 16983 3290 16989 3292
rect 16743 3238 16745 3290
rect 16925 3238 16927 3290
rect 16681 3236 16687 3238
rect 16743 3236 16767 3238
rect 16823 3236 16847 3238
rect 16903 3236 16927 3238
rect 16983 3236 16989 3238
rect 16681 3227 16989 3236
rect 17236 3194 17264 7822
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 12544 1306 12572 2382
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 12748 2204 13056 2213
rect 12748 2202 12754 2204
rect 12810 2202 12834 2204
rect 12890 2202 12914 2204
rect 12970 2202 12994 2204
rect 13050 2202 13056 2204
rect 12810 2150 12812 2202
rect 12992 2150 12994 2202
rect 12748 2148 12754 2150
rect 12810 2148 12834 2150
rect 12890 2148 12914 2150
rect 12970 2148 12994 2150
rect 13050 2148 13056 2150
rect 12748 2139 13056 2148
rect 13740 2106 13768 2246
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 12544 1278 12664 1306
rect 12636 800 12664 1278
rect 846 0 902 800
rect 2318 0 2374 800
rect 3790 0 3846 800
rect 5262 0 5318 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 13818 368 13874 377
rect 13924 354 13952 2382
rect 14108 800 14136 2382
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 13874 326 13952 354
rect 13818 303 13874 312
rect 14094 0 14150 800
rect 15212 762 15240 2314
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 2106 15516 2246
rect 15856 2106 15884 2382
rect 16132 2106 16160 2382
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16224 2106 16252 2246
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 15844 2100 15896 2106
rect 15844 2042 15896 2048
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16316 1193 16344 2246
rect 16592 2009 16620 2450
rect 16681 2204 16989 2213
rect 16681 2202 16687 2204
rect 16743 2202 16767 2204
rect 16823 2202 16847 2204
rect 16903 2202 16927 2204
rect 16983 2202 16989 2204
rect 16743 2150 16745 2202
rect 16925 2150 16927 2202
rect 16681 2148 16687 2150
rect 16743 2148 16767 2150
rect 16823 2148 16847 2150
rect 16903 2148 16927 2150
rect 16983 2148 16989 2150
rect 16681 2139 16989 2148
rect 16578 2000 16634 2009
rect 16578 1935 16634 1944
rect 16302 1184 16358 1193
rect 16302 1119 16358 1128
rect 15488 870 15608 898
rect 15488 762 15516 870
rect 15580 800 15608 870
rect 15212 734 15516 762
rect 15566 0 15622 800
<< via2 >>
rect 14922 17448 14978 17504
rect 938 15816 994 15872
rect 1490 16632 1546 16688
rect 2922 15802 2978 15804
rect 3002 15802 3058 15804
rect 3082 15802 3138 15804
rect 3162 15802 3218 15804
rect 2922 15750 2968 15802
rect 2968 15750 2978 15802
rect 3002 15750 3032 15802
rect 3032 15750 3044 15802
rect 3044 15750 3058 15802
rect 3082 15750 3096 15802
rect 3096 15750 3108 15802
rect 3108 15750 3138 15802
rect 3162 15750 3172 15802
rect 3172 15750 3218 15802
rect 2922 15748 2978 15750
rect 3002 15748 3058 15750
rect 3082 15748 3138 15750
rect 3162 15748 3218 15750
rect 6855 15802 6911 15804
rect 6935 15802 6991 15804
rect 7015 15802 7071 15804
rect 7095 15802 7151 15804
rect 6855 15750 6901 15802
rect 6901 15750 6911 15802
rect 6935 15750 6965 15802
rect 6965 15750 6977 15802
rect 6977 15750 6991 15802
rect 7015 15750 7029 15802
rect 7029 15750 7041 15802
rect 7041 15750 7071 15802
rect 7095 15750 7105 15802
rect 7105 15750 7151 15802
rect 6855 15748 6911 15750
rect 6935 15748 6991 15750
rect 7015 15748 7071 15750
rect 7095 15748 7151 15750
rect 10788 15802 10844 15804
rect 10868 15802 10924 15804
rect 10948 15802 11004 15804
rect 11028 15802 11084 15804
rect 10788 15750 10834 15802
rect 10834 15750 10844 15802
rect 10868 15750 10898 15802
rect 10898 15750 10910 15802
rect 10910 15750 10924 15802
rect 10948 15750 10962 15802
rect 10962 15750 10974 15802
rect 10974 15750 11004 15802
rect 11028 15750 11038 15802
rect 11038 15750 11084 15802
rect 10788 15748 10844 15750
rect 10868 15748 10924 15750
rect 10948 15748 11004 15750
rect 11028 15748 11084 15750
rect 2226 15136 2282 15192
rect 938 14184 994 14240
rect 1490 13640 1546 13696
rect 938 12588 940 12608
rect 940 12588 992 12608
rect 992 12588 994 12608
rect 938 12552 994 12588
rect 938 11736 994 11792
rect 2922 14714 2978 14716
rect 3002 14714 3058 14716
rect 3082 14714 3138 14716
rect 3162 14714 3218 14716
rect 2922 14662 2968 14714
rect 2968 14662 2978 14714
rect 3002 14662 3032 14714
rect 3032 14662 3044 14714
rect 3044 14662 3058 14714
rect 3082 14662 3096 14714
rect 3096 14662 3108 14714
rect 3108 14662 3138 14714
rect 3162 14662 3172 14714
rect 3172 14662 3218 14714
rect 2922 14660 2978 14662
rect 3002 14660 3058 14662
rect 3082 14660 3138 14662
rect 3162 14660 3218 14662
rect 2922 13626 2978 13628
rect 3002 13626 3058 13628
rect 3082 13626 3138 13628
rect 3162 13626 3218 13628
rect 2922 13574 2968 13626
rect 2968 13574 2978 13626
rect 3002 13574 3032 13626
rect 3032 13574 3044 13626
rect 3044 13574 3058 13626
rect 3082 13574 3096 13626
rect 3096 13574 3108 13626
rect 3108 13574 3138 13626
rect 3162 13574 3172 13626
rect 3172 13574 3218 13626
rect 2922 13572 2978 13574
rect 3002 13572 3058 13574
rect 3082 13572 3138 13574
rect 3162 13572 3218 13574
rect 2922 12538 2978 12540
rect 3002 12538 3058 12540
rect 3082 12538 3138 12540
rect 3162 12538 3218 12540
rect 2922 12486 2968 12538
rect 2968 12486 2978 12538
rect 3002 12486 3032 12538
rect 3032 12486 3044 12538
rect 3044 12486 3058 12538
rect 3082 12486 3096 12538
rect 3096 12486 3108 12538
rect 3108 12486 3138 12538
rect 3162 12486 3172 12538
rect 3172 12486 3218 12538
rect 2922 12484 2978 12486
rect 3002 12484 3058 12486
rect 3082 12484 3138 12486
rect 3162 12484 3218 12486
rect 2922 11450 2978 11452
rect 3002 11450 3058 11452
rect 3082 11450 3138 11452
rect 3162 11450 3218 11452
rect 2922 11398 2968 11450
rect 2968 11398 2978 11450
rect 3002 11398 3032 11450
rect 3032 11398 3044 11450
rect 3044 11398 3058 11450
rect 3082 11398 3096 11450
rect 3096 11398 3108 11450
rect 3108 11398 3138 11450
rect 3162 11398 3172 11450
rect 3172 11398 3218 11450
rect 2922 11396 2978 11398
rect 3002 11396 3058 11398
rect 3082 11396 3138 11398
rect 3162 11396 3218 11398
rect 1398 10920 1454 10976
rect 938 10104 994 10160
rect 2922 10362 2978 10364
rect 3002 10362 3058 10364
rect 3082 10362 3138 10364
rect 3162 10362 3218 10364
rect 2922 10310 2968 10362
rect 2968 10310 2978 10362
rect 3002 10310 3032 10362
rect 3032 10310 3044 10362
rect 3044 10310 3058 10362
rect 3082 10310 3096 10362
rect 3096 10310 3108 10362
rect 3108 10310 3138 10362
rect 3162 10310 3172 10362
rect 3172 10310 3218 10362
rect 2922 10308 2978 10310
rect 3002 10308 3058 10310
rect 3082 10308 3138 10310
rect 3162 10308 3218 10310
rect 3330 9560 3386 9616
rect 2922 9274 2978 9276
rect 3002 9274 3058 9276
rect 3082 9274 3138 9276
rect 3162 9274 3218 9276
rect 2922 9222 2968 9274
rect 2968 9222 2978 9274
rect 3002 9222 3032 9274
rect 3032 9222 3044 9274
rect 3044 9222 3058 9274
rect 3082 9222 3096 9274
rect 3096 9222 3108 9274
rect 3108 9222 3138 9274
rect 3162 9222 3172 9274
rect 3172 9222 3218 9274
rect 2922 9220 2978 9222
rect 3002 9220 3058 9222
rect 3082 9220 3138 9222
rect 3162 9220 3218 9222
rect 938 8472 994 8528
rect 2922 8186 2978 8188
rect 3002 8186 3058 8188
rect 3082 8186 3138 8188
rect 3162 8186 3218 8188
rect 2922 8134 2968 8186
rect 2968 8134 2978 8186
rect 3002 8134 3032 8186
rect 3032 8134 3044 8186
rect 3044 8134 3058 8186
rect 3082 8134 3096 8186
rect 3096 8134 3108 8186
rect 3108 8134 3138 8186
rect 3162 8134 3172 8186
rect 3172 8134 3218 8186
rect 2922 8132 2978 8134
rect 3002 8132 3058 8134
rect 3082 8132 3138 8134
rect 3162 8132 3218 8134
rect 938 7656 994 7712
rect 2922 7098 2978 7100
rect 3002 7098 3058 7100
rect 3082 7098 3138 7100
rect 3162 7098 3218 7100
rect 2922 7046 2968 7098
rect 2968 7046 2978 7098
rect 3002 7046 3032 7098
rect 3032 7046 3044 7098
rect 3044 7046 3058 7098
rect 3082 7046 3096 7098
rect 3096 7046 3108 7098
rect 3108 7046 3138 7098
rect 3162 7046 3172 7098
rect 3172 7046 3218 7098
rect 2922 7044 2978 7046
rect 3002 7044 3058 7046
rect 3082 7044 3138 7046
rect 3162 7044 3218 7046
rect 1490 6840 1546 6896
rect 938 6060 940 6080
rect 940 6060 992 6080
rect 992 6060 994 6080
rect 938 6024 994 6060
rect 2922 6010 2978 6012
rect 3002 6010 3058 6012
rect 3082 6010 3138 6012
rect 3162 6010 3218 6012
rect 2922 5958 2968 6010
rect 2968 5958 2978 6010
rect 3002 5958 3032 6010
rect 3032 5958 3044 6010
rect 3044 5958 3058 6010
rect 3082 5958 3096 6010
rect 3096 5958 3108 6010
rect 3108 5958 3138 6010
rect 3162 5958 3172 6010
rect 3172 5958 3218 6010
rect 2922 5956 2978 5958
rect 3002 5956 3058 5958
rect 3082 5956 3138 5958
rect 3162 5956 3218 5958
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 2922 4922 2978 4924
rect 3002 4922 3058 4924
rect 3082 4922 3138 4924
rect 3162 4922 3218 4924
rect 2922 4870 2968 4922
rect 2968 4870 2978 4922
rect 3002 4870 3032 4922
rect 3032 4870 3044 4922
rect 3044 4870 3058 4922
rect 3082 4870 3096 4922
rect 3096 4870 3108 4922
rect 3108 4870 3138 4922
rect 3162 4870 3172 4922
rect 3172 4870 3218 4922
rect 2922 4868 2978 4870
rect 3002 4868 3058 4870
rect 3082 4868 3138 4870
rect 3162 4868 3218 4870
rect 938 4392 994 4448
rect 2922 3834 2978 3836
rect 3002 3834 3058 3836
rect 3082 3834 3138 3836
rect 3162 3834 3218 3836
rect 2922 3782 2968 3834
rect 2968 3782 2978 3834
rect 3002 3782 3032 3834
rect 3032 3782 3044 3834
rect 3044 3782 3058 3834
rect 3082 3782 3096 3834
rect 3096 3782 3108 3834
rect 3108 3782 3138 3834
rect 3162 3782 3172 3834
rect 3172 3782 3218 3834
rect 2922 3780 2978 3782
rect 3002 3780 3058 3782
rect 3082 3780 3138 3782
rect 3162 3780 3218 3782
rect 938 3576 994 3632
rect 4888 15258 4944 15260
rect 4968 15258 5024 15260
rect 5048 15258 5104 15260
rect 5128 15258 5184 15260
rect 4888 15206 4934 15258
rect 4934 15206 4944 15258
rect 4968 15206 4998 15258
rect 4998 15206 5010 15258
rect 5010 15206 5024 15258
rect 5048 15206 5062 15258
rect 5062 15206 5074 15258
rect 5074 15206 5104 15258
rect 5128 15206 5138 15258
rect 5138 15206 5184 15258
rect 4888 15204 4944 15206
rect 4968 15204 5024 15206
rect 5048 15204 5104 15206
rect 5128 15204 5184 15206
rect 4888 14170 4944 14172
rect 4968 14170 5024 14172
rect 5048 14170 5104 14172
rect 5128 14170 5184 14172
rect 4888 14118 4934 14170
rect 4934 14118 4944 14170
rect 4968 14118 4998 14170
rect 4998 14118 5010 14170
rect 5010 14118 5024 14170
rect 5048 14118 5062 14170
rect 5062 14118 5074 14170
rect 5074 14118 5104 14170
rect 5128 14118 5138 14170
rect 5138 14118 5184 14170
rect 4888 14116 4944 14118
rect 4968 14116 5024 14118
rect 5048 14116 5104 14118
rect 5128 14116 5184 14118
rect 4888 13082 4944 13084
rect 4968 13082 5024 13084
rect 5048 13082 5104 13084
rect 5128 13082 5184 13084
rect 4888 13030 4934 13082
rect 4934 13030 4944 13082
rect 4968 13030 4998 13082
rect 4998 13030 5010 13082
rect 5010 13030 5024 13082
rect 5048 13030 5062 13082
rect 5062 13030 5074 13082
rect 5074 13030 5104 13082
rect 5128 13030 5138 13082
rect 5138 13030 5184 13082
rect 4888 13028 4944 13030
rect 4968 13028 5024 13030
rect 5048 13028 5104 13030
rect 5128 13028 5184 13030
rect 4888 11994 4944 11996
rect 4968 11994 5024 11996
rect 5048 11994 5104 11996
rect 5128 11994 5184 11996
rect 4888 11942 4934 11994
rect 4934 11942 4944 11994
rect 4968 11942 4998 11994
rect 4998 11942 5010 11994
rect 5010 11942 5024 11994
rect 5048 11942 5062 11994
rect 5062 11942 5074 11994
rect 5074 11942 5104 11994
rect 5128 11942 5138 11994
rect 5138 11942 5184 11994
rect 4888 11940 4944 11942
rect 4968 11940 5024 11942
rect 5048 11940 5104 11942
rect 5128 11940 5184 11942
rect 4888 10906 4944 10908
rect 4968 10906 5024 10908
rect 5048 10906 5104 10908
rect 5128 10906 5184 10908
rect 4888 10854 4934 10906
rect 4934 10854 4944 10906
rect 4968 10854 4998 10906
rect 4998 10854 5010 10906
rect 5010 10854 5024 10906
rect 5048 10854 5062 10906
rect 5062 10854 5074 10906
rect 5074 10854 5104 10906
rect 5128 10854 5138 10906
rect 5138 10854 5184 10906
rect 4888 10852 4944 10854
rect 4968 10852 5024 10854
rect 5048 10852 5104 10854
rect 5128 10852 5184 10854
rect 8821 15258 8877 15260
rect 8901 15258 8957 15260
rect 8981 15258 9037 15260
rect 9061 15258 9117 15260
rect 8821 15206 8867 15258
rect 8867 15206 8877 15258
rect 8901 15206 8931 15258
rect 8931 15206 8943 15258
rect 8943 15206 8957 15258
rect 8981 15206 8995 15258
rect 8995 15206 9007 15258
rect 9007 15206 9037 15258
rect 9061 15206 9071 15258
rect 9071 15206 9117 15258
rect 8821 15204 8877 15206
rect 8901 15204 8957 15206
rect 8981 15204 9037 15206
rect 9061 15204 9117 15206
rect 6855 14714 6911 14716
rect 6935 14714 6991 14716
rect 7015 14714 7071 14716
rect 7095 14714 7151 14716
rect 6855 14662 6901 14714
rect 6901 14662 6911 14714
rect 6935 14662 6965 14714
rect 6965 14662 6977 14714
rect 6977 14662 6991 14714
rect 7015 14662 7029 14714
rect 7029 14662 7041 14714
rect 7041 14662 7071 14714
rect 7095 14662 7105 14714
rect 7105 14662 7151 14714
rect 6855 14660 6911 14662
rect 6935 14660 6991 14662
rect 7015 14660 7071 14662
rect 7095 14660 7151 14662
rect 6855 13626 6911 13628
rect 6935 13626 6991 13628
rect 7015 13626 7071 13628
rect 7095 13626 7151 13628
rect 6855 13574 6901 13626
rect 6901 13574 6911 13626
rect 6935 13574 6965 13626
rect 6965 13574 6977 13626
rect 6977 13574 6991 13626
rect 7015 13574 7029 13626
rect 7029 13574 7041 13626
rect 7041 13574 7071 13626
rect 7095 13574 7105 13626
rect 7105 13574 7151 13626
rect 6855 13572 6911 13574
rect 6935 13572 6991 13574
rect 7015 13572 7071 13574
rect 7095 13572 7151 13574
rect 6855 12538 6911 12540
rect 6935 12538 6991 12540
rect 7015 12538 7071 12540
rect 7095 12538 7151 12540
rect 6855 12486 6901 12538
rect 6901 12486 6911 12538
rect 6935 12486 6965 12538
rect 6965 12486 6977 12538
rect 6977 12486 6991 12538
rect 7015 12486 7029 12538
rect 7029 12486 7041 12538
rect 7041 12486 7071 12538
rect 7095 12486 7105 12538
rect 7105 12486 7151 12538
rect 6855 12484 6911 12486
rect 6935 12484 6991 12486
rect 7015 12484 7071 12486
rect 7095 12484 7151 12486
rect 4888 9818 4944 9820
rect 4968 9818 5024 9820
rect 5048 9818 5104 9820
rect 5128 9818 5184 9820
rect 4888 9766 4934 9818
rect 4934 9766 4944 9818
rect 4968 9766 4998 9818
rect 4998 9766 5010 9818
rect 5010 9766 5024 9818
rect 5048 9766 5062 9818
rect 5062 9766 5074 9818
rect 5074 9766 5104 9818
rect 5128 9766 5138 9818
rect 5138 9766 5184 9818
rect 4888 9764 4944 9766
rect 4968 9764 5024 9766
rect 5048 9764 5104 9766
rect 5128 9764 5184 9766
rect 5446 9596 5448 9616
rect 5448 9596 5500 9616
rect 5500 9596 5502 9616
rect 5446 9560 5502 9596
rect 4888 8730 4944 8732
rect 4968 8730 5024 8732
rect 5048 8730 5104 8732
rect 5128 8730 5184 8732
rect 4888 8678 4934 8730
rect 4934 8678 4944 8730
rect 4968 8678 4998 8730
rect 4998 8678 5010 8730
rect 5010 8678 5024 8730
rect 5048 8678 5062 8730
rect 5062 8678 5074 8730
rect 5074 8678 5104 8730
rect 5128 8678 5138 8730
rect 5138 8678 5184 8730
rect 4888 8676 4944 8678
rect 4968 8676 5024 8678
rect 5048 8676 5104 8678
rect 5128 8676 5184 8678
rect 4888 7642 4944 7644
rect 4968 7642 5024 7644
rect 5048 7642 5104 7644
rect 5128 7642 5184 7644
rect 4888 7590 4934 7642
rect 4934 7590 4944 7642
rect 4968 7590 4998 7642
rect 4998 7590 5010 7642
rect 5010 7590 5024 7642
rect 5048 7590 5062 7642
rect 5062 7590 5074 7642
rect 5074 7590 5104 7642
rect 5128 7590 5138 7642
rect 5138 7590 5184 7642
rect 4888 7588 4944 7590
rect 4968 7588 5024 7590
rect 5048 7588 5104 7590
rect 5128 7588 5184 7590
rect 3330 6160 3386 6216
rect 4888 6554 4944 6556
rect 4968 6554 5024 6556
rect 5048 6554 5104 6556
rect 5128 6554 5184 6556
rect 4888 6502 4934 6554
rect 4934 6502 4944 6554
rect 4968 6502 4998 6554
rect 4998 6502 5010 6554
rect 5010 6502 5024 6554
rect 5048 6502 5062 6554
rect 5062 6502 5074 6554
rect 5074 6502 5104 6554
rect 5128 6502 5138 6554
rect 5138 6502 5184 6554
rect 4888 6500 4944 6502
rect 4968 6500 5024 6502
rect 5048 6500 5104 6502
rect 5128 6500 5184 6502
rect 4888 5466 4944 5468
rect 4968 5466 5024 5468
rect 5048 5466 5104 5468
rect 5128 5466 5184 5468
rect 4888 5414 4934 5466
rect 4934 5414 4944 5466
rect 4968 5414 4998 5466
rect 4998 5414 5010 5466
rect 5010 5414 5024 5466
rect 5048 5414 5062 5466
rect 5062 5414 5074 5466
rect 5074 5414 5104 5466
rect 5128 5414 5138 5466
rect 5138 5414 5184 5466
rect 4888 5412 4944 5414
rect 4968 5412 5024 5414
rect 5048 5412 5104 5414
rect 5128 5412 5184 5414
rect 5630 6860 5686 6896
rect 5630 6840 5632 6860
rect 5632 6840 5684 6860
rect 5684 6840 5686 6860
rect 6855 11450 6911 11452
rect 6935 11450 6991 11452
rect 7015 11450 7071 11452
rect 7095 11450 7151 11452
rect 6855 11398 6901 11450
rect 6901 11398 6911 11450
rect 6935 11398 6965 11450
rect 6965 11398 6977 11450
rect 6977 11398 6991 11450
rect 7015 11398 7029 11450
rect 7029 11398 7041 11450
rect 7041 11398 7071 11450
rect 7095 11398 7105 11450
rect 7105 11398 7151 11450
rect 6855 11396 6911 11398
rect 6935 11396 6991 11398
rect 7015 11396 7071 11398
rect 7095 11396 7151 11398
rect 6855 10362 6911 10364
rect 6935 10362 6991 10364
rect 7015 10362 7071 10364
rect 7095 10362 7151 10364
rect 6855 10310 6901 10362
rect 6901 10310 6911 10362
rect 6935 10310 6965 10362
rect 6965 10310 6977 10362
rect 6977 10310 6991 10362
rect 7015 10310 7029 10362
rect 7029 10310 7041 10362
rect 7041 10310 7071 10362
rect 7095 10310 7105 10362
rect 7105 10310 7151 10362
rect 6855 10308 6911 10310
rect 6935 10308 6991 10310
rect 7015 10308 7071 10310
rect 7095 10308 7151 10310
rect 6855 9274 6911 9276
rect 6935 9274 6991 9276
rect 7015 9274 7071 9276
rect 7095 9274 7151 9276
rect 6855 9222 6901 9274
rect 6901 9222 6911 9274
rect 6935 9222 6965 9274
rect 6965 9222 6977 9274
rect 6977 9222 6991 9274
rect 7015 9222 7029 9274
rect 7029 9222 7041 9274
rect 7041 9222 7071 9274
rect 7095 9222 7105 9274
rect 7105 9222 7151 9274
rect 6855 9220 6911 9222
rect 6935 9220 6991 9222
rect 7015 9220 7071 9222
rect 7095 9220 7151 9222
rect 6855 8186 6911 8188
rect 6935 8186 6991 8188
rect 7015 8186 7071 8188
rect 7095 8186 7151 8188
rect 6855 8134 6901 8186
rect 6901 8134 6911 8186
rect 6935 8134 6965 8186
rect 6965 8134 6977 8186
rect 6977 8134 6991 8186
rect 7015 8134 7029 8186
rect 7029 8134 7041 8186
rect 7041 8134 7071 8186
rect 7095 8134 7105 8186
rect 7105 8134 7151 8186
rect 6855 8132 6911 8134
rect 6935 8132 6991 8134
rect 7015 8132 7071 8134
rect 7095 8132 7151 8134
rect 8821 14170 8877 14172
rect 8901 14170 8957 14172
rect 8981 14170 9037 14172
rect 9061 14170 9117 14172
rect 8821 14118 8867 14170
rect 8867 14118 8877 14170
rect 8901 14118 8931 14170
rect 8931 14118 8943 14170
rect 8943 14118 8957 14170
rect 8981 14118 8995 14170
rect 8995 14118 9007 14170
rect 9007 14118 9037 14170
rect 9061 14118 9071 14170
rect 9071 14118 9117 14170
rect 8821 14116 8877 14118
rect 8901 14116 8957 14118
rect 8981 14116 9037 14118
rect 9061 14116 9117 14118
rect 8821 13082 8877 13084
rect 8901 13082 8957 13084
rect 8981 13082 9037 13084
rect 9061 13082 9117 13084
rect 8821 13030 8867 13082
rect 8867 13030 8877 13082
rect 8901 13030 8931 13082
rect 8931 13030 8943 13082
rect 8943 13030 8957 13082
rect 8981 13030 8995 13082
rect 8995 13030 9007 13082
rect 9007 13030 9037 13082
rect 9061 13030 9071 13082
rect 9071 13030 9117 13082
rect 8821 13028 8877 13030
rect 8901 13028 8957 13030
rect 8981 13028 9037 13030
rect 9061 13028 9117 13030
rect 8821 11994 8877 11996
rect 8901 11994 8957 11996
rect 8981 11994 9037 11996
rect 9061 11994 9117 11996
rect 8821 11942 8867 11994
rect 8867 11942 8877 11994
rect 8901 11942 8931 11994
rect 8931 11942 8943 11994
rect 8943 11942 8957 11994
rect 8981 11942 8995 11994
rect 8995 11942 9007 11994
rect 9007 11942 9037 11994
rect 9061 11942 9071 11994
rect 9071 11942 9117 11994
rect 8821 11940 8877 11942
rect 8901 11940 8957 11942
rect 8981 11940 9037 11942
rect 9061 11940 9117 11942
rect 14721 15802 14777 15804
rect 14801 15802 14857 15804
rect 14881 15802 14937 15804
rect 14961 15802 15017 15804
rect 14721 15750 14767 15802
rect 14767 15750 14777 15802
rect 14801 15750 14831 15802
rect 14831 15750 14843 15802
rect 14843 15750 14857 15802
rect 14881 15750 14895 15802
rect 14895 15750 14907 15802
rect 14907 15750 14937 15802
rect 14961 15750 14971 15802
rect 14971 15750 15017 15802
rect 14721 15748 14777 15750
rect 14801 15748 14857 15750
rect 14881 15748 14937 15750
rect 14961 15748 15017 15750
rect 16486 16632 16542 16688
rect 12754 15258 12810 15260
rect 12834 15258 12890 15260
rect 12914 15258 12970 15260
rect 12994 15258 13050 15260
rect 12754 15206 12800 15258
rect 12800 15206 12810 15258
rect 12834 15206 12864 15258
rect 12864 15206 12876 15258
rect 12876 15206 12890 15258
rect 12914 15206 12928 15258
rect 12928 15206 12940 15258
rect 12940 15206 12970 15258
rect 12994 15206 13004 15258
rect 13004 15206 13050 15258
rect 12754 15204 12810 15206
rect 12834 15204 12890 15206
rect 12914 15204 12970 15206
rect 12994 15204 13050 15206
rect 10788 14714 10844 14716
rect 10868 14714 10924 14716
rect 10948 14714 11004 14716
rect 11028 14714 11084 14716
rect 10788 14662 10834 14714
rect 10834 14662 10844 14714
rect 10868 14662 10898 14714
rect 10898 14662 10910 14714
rect 10910 14662 10924 14714
rect 10948 14662 10962 14714
rect 10962 14662 10974 14714
rect 10974 14662 11004 14714
rect 11028 14662 11038 14714
rect 11038 14662 11084 14714
rect 10788 14660 10844 14662
rect 10868 14660 10924 14662
rect 10948 14660 11004 14662
rect 11028 14660 11084 14662
rect 10788 13626 10844 13628
rect 10868 13626 10924 13628
rect 10948 13626 11004 13628
rect 11028 13626 11084 13628
rect 10788 13574 10834 13626
rect 10834 13574 10844 13626
rect 10868 13574 10898 13626
rect 10898 13574 10910 13626
rect 10910 13574 10924 13626
rect 10948 13574 10962 13626
rect 10962 13574 10974 13626
rect 10974 13574 11004 13626
rect 11028 13574 11038 13626
rect 11038 13574 11084 13626
rect 10788 13572 10844 13574
rect 10868 13572 10924 13574
rect 10948 13572 11004 13574
rect 11028 13572 11084 13574
rect 10788 12538 10844 12540
rect 10868 12538 10924 12540
rect 10948 12538 11004 12540
rect 11028 12538 11084 12540
rect 10788 12486 10834 12538
rect 10834 12486 10844 12538
rect 10868 12486 10898 12538
rect 10898 12486 10910 12538
rect 10910 12486 10924 12538
rect 10948 12486 10962 12538
rect 10962 12486 10974 12538
rect 10974 12486 11004 12538
rect 11028 12486 11038 12538
rect 11038 12486 11084 12538
rect 10788 12484 10844 12486
rect 10868 12484 10924 12486
rect 10948 12484 11004 12486
rect 11028 12484 11084 12486
rect 8821 10906 8877 10908
rect 8901 10906 8957 10908
rect 8981 10906 9037 10908
rect 9061 10906 9117 10908
rect 8821 10854 8867 10906
rect 8867 10854 8877 10906
rect 8901 10854 8931 10906
rect 8931 10854 8943 10906
rect 8943 10854 8957 10906
rect 8981 10854 8995 10906
rect 8995 10854 9007 10906
rect 9007 10854 9037 10906
rect 9061 10854 9071 10906
rect 9071 10854 9117 10906
rect 8821 10852 8877 10854
rect 8901 10852 8957 10854
rect 8981 10852 9037 10854
rect 9061 10852 9117 10854
rect 8821 9818 8877 9820
rect 8901 9818 8957 9820
rect 8981 9818 9037 9820
rect 9061 9818 9117 9820
rect 8821 9766 8867 9818
rect 8867 9766 8877 9818
rect 8901 9766 8931 9818
rect 8931 9766 8943 9818
rect 8943 9766 8957 9818
rect 8981 9766 8995 9818
rect 8995 9766 9007 9818
rect 9007 9766 9037 9818
rect 9061 9766 9071 9818
rect 9071 9766 9117 9818
rect 8821 9764 8877 9766
rect 8901 9764 8957 9766
rect 8981 9764 9037 9766
rect 9061 9764 9117 9766
rect 6855 7098 6911 7100
rect 6935 7098 6991 7100
rect 7015 7098 7071 7100
rect 7095 7098 7151 7100
rect 6855 7046 6901 7098
rect 6901 7046 6911 7098
rect 6935 7046 6965 7098
rect 6965 7046 6977 7098
rect 6977 7046 6991 7098
rect 7015 7046 7029 7098
rect 7029 7046 7041 7098
rect 7041 7046 7071 7098
rect 7095 7046 7105 7098
rect 7105 7046 7151 7098
rect 6855 7044 6911 7046
rect 6935 7044 6991 7046
rect 7015 7044 7071 7046
rect 7095 7044 7151 7046
rect 6458 6296 6514 6352
rect 4888 4378 4944 4380
rect 4968 4378 5024 4380
rect 5048 4378 5104 4380
rect 5128 4378 5184 4380
rect 4888 4326 4934 4378
rect 4934 4326 4944 4378
rect 4968 4326 4998 4378
rect 4998 4326 5010 4378
rect 5010 4326 5024 4378
rect 5048 4326 5062 4378
rect 5062 4326 5074 4378
rect 5074 4326 5104 4378
rect 5128 4326 5138 4378
rect 5138 4326 5184 4378
rect 4888 4324 4944 4326
rect 4968 4324 5024 4326
rect 5048 4324 5104 4326
rect 5128 4324 5184 4326
rect 938 2796 940 2816
rect 940 2796 992 2816
rect 992 2796 994 2816
rect 938 2760 994 2796
rect 2922 2746 2978 2748
rect 3002 2746 3058 2748
rect 3082 2746 3138 2748
rect 3162 2746 3218 2748
rect 2922 2694 2968 2746
rect 2968 2694 2978 2746
rect 3002 2694 3032 2746
rect 3032 2694 3044 2746
rect 3044 2694 3058 2746
rect 3082 2694 3096 2746
rect 3096 2694 3108 2746
rect 3108 2694 3138 2746
rect 3162 2694 3172 2746
rect 3172 2694 3218 2746
rect 2922 2692 2978 2694
rect 3002 2692 3058 2694
rect 3082 2692 3138 2694
rect 3162 2692 3218 2694
rect 4888 3290 4944 3292
rect 4968 3290 5024 3292
rect 5048 3290 5104 3292
rect 5128 3290 5184 3292
rect 4888 3238 4934 3290
rect 4934 3238 4944 3290
rect 4968 3238 4998 3290
rect 4998 3238 5010 3290
rect 5010 3238 5024 3290
rect 5048 3238 5062 3290
rect 5062 3238 5074 3290
rect 5074 3238 5104 3290
rect 5128 3238 5138 3290
rect 5138 3238 5184 3290
rect 4888 3236 4944 3238
rect 4968 3236 5024 3238
rect 5048 3236 5104 3238
rect 5128 3236 5184 3238
rect 6855 6010 6911 6012
rect 6935 6010 6991 6012
rect 7015 6010 7071 6012
rect 7095 6010 7151 6012
rect 6855 5958 6901 6010
rect 6901 5958 6911 6010
rect 6935 5958 6965 6010
rect 6965 5958 6977 6010
rect 6977 5958 6991 6010
rect 7015 5958 7029 6010
rect 7029 5958 7041 6010
rect 7041 5958 7071 6010
rect 7095 5958 7105 6010
rect 7105 5958 7151 6010
rect 6855 5956 6911 5958
rect 6935 5956 6991 5958
rect 7015 5956 7071 5958
rect 7095 5956 7151 5958
rect 9310 9016 9366 9072
rect 8821 8730 8877 8732
rect 8901 8730 8957 8732
rect 8981 8730 9037 8732
rect 9061 8730 9117 8732
rect 8821 8678 8867 8730
rect 8867 8678 8877 8730
rect 8901 8678 8931 8730
rect 8931 8678 8943 8730
rect 8943 8678 8957 8730
rect 8981 8678 8995 8730
rect 8995 8678 9007 8730
rect 9007 8678 9037 8730
rect 9061 8678 9071 8730
rect 9071 8678 9117 8730
rect 8821 8676 8877 8678
rect 8901 8676 8957 8678
rect 8981 8676 9037 8678
rect 9061 8676 9117 8678
rect 7838 5772 7894 5808
rect 7838 5752 7840 5772
rect 7840 5752 7892 5772
rect 7892 5752 7894 5772
rect 7838 5616 7894 5672
rect 6855 4922 6911 4924
rect 6935 4922 6991 4924
rect 7015 4922 7071 4924
rect 7095 4922 7151 4924
rect 6855 4870 6901 4922
rect 6901 4870 6911 4922
rect 6935 4870 6965 4922
rect 6965 4870 6977 4922
rect 6977 4870 6991 4922
rect 7015 4870 7029 4922
rect 7029 4870 7041 4922
rect 7041 4870 7071 4922
rect 7095 4870 7105 4922
rect 7105 4870 7151 4922
rect 6855 4868 6911 4870
rect 6935 4868 6991 4870
rect 7015 4868 7071 4870
rect 7095 4868 7151 4870
rect 7378 5228 7434 5264
rect 7378 5208 7380 5228
rect 7380 5208 7432 5228
rect 7432 5208 7434 5228
rect 6855 3834 6911 3836
rect 6935 3834 6991 3836
rect 7015 3834 7071 3836
rect 7095 3834 7151 3836
rect 6855 3782 6901 3834
rect 6901 3782 6911 3834
rect 6935 3782 6965 3834
rect 6965 3782 6977 3834
rect 6977 3782 6991 3834
rect 7015 3782 7029 3834
rect 7029 3782 7041 3834
rect 7041 3782 7071 3834
rect 7095 3782 7105 3834
rect 7105 3782 7151 3834
rect 6855 3780 6911 3782
rect 6935 3780 6991 3782
rect 7015 3780 7071 3782
rect 7095 3780 7151 3782
rect 8022 6160 8078 6216
rect 8821 7642 8877 7644
rect 8901 7642 8957 7644
rect 8981 7642 9037 7644
rect 9061 7642 9117 7644
rect 8821 7590 8867 7642
rect 8867 7590 8877 7642
rect 8901 7590 8931 7642
rect 8931 7590 8943 7642
rect 8943 7590 8957 7642
rect 8981 7590 8995 7642
rect 8995 7590 9007 7642
rect 9007 7590 9037 7642
rect 9061 7590 9071 7642
rect 9071 7590 9117 7642
rect 8821 7588 8877 7590
rect 8901 7588 8957 7590
rect 8981 7588 9037 7590
rect 9061 7588 9117 7590
rect 8821 6554 8877 6556
rect 8901 6554 8957 6556
rect 8981 6554 9037 6556
rect 9061 6554 9117 6556
rect 8821 6502 8867 6554
rect 8867 6502 8877 6554
rect 8901 6502 8931 6554
rect 8931 6502 8943 6554
rect 8943 6502 8957 6554
rect 8981 6502 8995 6554
rect 8995 6502 9007 6554
rect 9007 6502 9037 6554
rect 9061 6502 9071 6554
rect 9071 6502 9117 6554
rect 8821 6500 8877 6502
rect 8901 6500 8957 6502
rect 8981 6500 9037 6502
rect 9061 6500 9117 6502
rect 8758 6316 8814 6352
rect 8758 6296 8760 6316
rect 8760 6296 8812 6316
rect 8812 6296 8814 6316
rect 8666 5772 8722 5808
rect 8666 5752 8668 5772
rect 8668 5752 8720 5772
rect 8720 5752 8722 5772
rect 8942 5616 8998 5672
rect 8821 5466 8877 5468
rect 8901 5466 8957 5468
rect 8981 5466 9037 5468
rect 9061 5466 9117 5468
rect 8821 5414 8867 5466
rect 8867 5414 8877 5466
rect 8901 5414 8931 5466
rect 8931 5414 8943 5466
rect 8943 5414 8957 5466
rect 8981 5414 8995 5466
rect 8995 5414 9007 5466
rect 9007 5414 9037 5466
rect 9061 5414 9071 5466
rect 9071 5414 9117 5466
rect 8821 5412 8877 5414
rect 8901 5412 8957 5414
rect 8981 5412 9037 5414
rect 9061 5412 9117 5414
rect 8942 5244 8944 5264
rect 8944 5244 8996 5264
rect 8996 5244 8998 5264
rect 8942 5208 8998 5244
rect 8821 4378 8877 4380
rect 8901 4378 8957 4380
rect 8981 4378 9037 4380
rect 9061 4378 9117 4380
rect 8821 4326 8867 4378
rect 8867 4326 8877 4378
rect 8901 4326 8931 4378
rect 8931 4326 8943 4378
rect 8943 4326 8957 4378
rect 8981 4326 8995 4378
rect 8995 4326 9007 4378
rect 9007 4326 9037 4378
rect 9061 4326 9071 4378
rect 9071 4326 9117 4378
rect 8821 4324 8877 4326
rect 8901 4324 8957 4326
rect 8981 4324 9037 4326
rect 9061 4324 9117 4326
rect 8821 3290 8877 3292
rect 8901 3290 8957 3292
rect 8981 3290 9037 3292
rect 9061 3290 9117 3292
rect 8821 3238 8867 3290
rect 8867 3238 8877 3290
rect 8901 3238 8931 3290
rect 8931 3238 8943 3290
rect 8943 3238 8957 3290
rect 8981 3238 8995 3290
rect 8995 3238 9007 3290
rect 9007 3238 9037 3290
rect 9061 3238 9071 3290
rect 9071 3238 9117 3290
rect 8821 3236 8877 3238
rect 8901 3236 8957 3238
rect 8981 3236 9037 3238
rect 9061 3236 9117 3238
rect 6855 2746 6911 2748
rect 6935 2746 6991 2748
rect 7015 2746 7071 2748
rect 7095 2746 7151 2748
rect 6855 2694 6901 2746
rect 6901 2694 6911 2746
rect 6935 2694 6965 2746
rect 6965 2694 6977 2746
rect 6977 2694 6991 2746
rect 7015 2694 7029 2746
rect 7029 2694 7041 2746
rect 7041 2694 7071 2746
rect 7095 2694 7105 2746
rect 7105 2694 7151 2746
rect 6855 2692 6911 2694
rect 6935 2692 6991 2694
rect 7015 2692 7071 2694
rect 7095 2692 7151 2694
rect 10788 11450 10844 11452
rect 10868 11450 10924 11452
rect 10948 11450 11004 11452
rect 11028 11450 11084 11452
rect 10788 11398 10834 11450
rect 10834 11398 10844 11450
rect 10868 11398 10898 11450
rect 10898 11398 10910 11450
rect 10910 11398 10924 11450
rect 10948 11398 10962 11450
rect 10962 11398 10974 11450
rect 10974 11398 11004 11450
rect 11028 11398 11038 11450
rect 11038 11398 11084 11450
rect 10788 11396 10844 11398
rect 10868 11396 10924 11398
rect 10948 11396 11004 11398
rect 11028 11396 11084 11398
rect 11518 11056 11574 11112
rect 10788 10362 10844 10364
rect 10868 10362 10924 10364
rect 10948 10362 11004 10364
rect 11028 10362 11084 10364
rect 10788 10310 10834 10362
rect 10834 10310 10844 10362
rect 10868 10310 10898 10362
rect 10898 10310 10910 10362
rect 10910 10310 10924 10362
rect 10948 10310 10962 10362
rect 10962 10310 10974 10362
rect 10974 10310 11004 10362
rect 11028 10310 11038 10362
rect 11038 10310 11084 10362
rect 10788 10308 10844 10310
rect 10868 10308 10924 10310
rect 10948 10308 11004 10310
rect 11028 10308 11084 10310
rect 10788 9274 10844 9276
rect 10868 9274 10924 9276
rect 10948 9274 11004 9276
rect 11028 9274 11084 9276
rect 10788 9222 10834 9274
rect 10834 9222 10844 9274
rect 10868 9222 10898 9274
rect 10898 9222 10910 9274
rect 10910 9222 10924 9274
rect 10948 9222 10962 9274
rect 10962 9222 10974 9274
rect 10974 9222 11004 9274
rect 11028 9222 11038 9274
rect 11038 9222 11084 9274
rect 10788 9220 10844 9222
rect 10868 9220 10924 9222
rect 10948 9220 11004 9222
rect 11028 9220 11084 9222
rect 10788 8186 10844 8188
rect 10868 8186 10924 8188
rect 10948 8186 11004 8188
rect 11028 8186 11084 8188
rect 10788 8134 10834 8186
rect 10834 8134 10844 8186
rect 10868 8134 10898 8186
rect 10898 8134 10910 8186
rect 10910 8134 10924 8186
rect 10948 8134 10962 8186
rect 10962 8134 10974 8186
rect 10974 8134 11004 8186
rect 11028 8134 11038 8186
rect 11038 8134 11084 8186
rect 10788 8132 10844 8134
rect 10868 8132 10924 8134
rect 10948 8132 11004 8134
rect 11028 8132 11084 8134
rect 10788 7098 10844 7100
rect 10868 7098 10924 7100
rect 10948 7098 11004 7100
rect 11028 7098 11084 7100
rect 10788 7046 10834 7098
rect 10834 7046 10844 7098
rect 10868 7046 10898 7098
rect 10898 7046 10910 7098
rect 10910 7046 10924 7098
rect 10948 7046 10962 7098
rect 10962 7046 10974 7098
rect 10974 7046 11004 7098
rect 11028 7046 11038 7098
rect 11038 7046 11084 7098
rect 10788 7044 10844 7046
rect 10868 7044 10924 7046
rect 10948 7044 11004 7046
rect 11028 7044 11084 7046
rect 11978 10104 12034 10160
rect 12254 9968 12310 10024
rect 12754 14170 12810 14172
rect 12834 14170 12890 14172
rect 12914 14170 12970 14172
rect 12994 14170 13050 14172
rect 12754 14118 12800 14170
rect 12800 14118 12810 14170
rect 12834 14118 12864 14170
rect 12864 14118 12876 14170
rect 12876 14118 12890 14170
rect 12914 14118 12928 14170
rect 12928 14118 12940 14170
rect 12940 14118 12970 14170
rect 12994 14118 13004 14170
rect 13004 14118 13050 14170
rect 12754 14116 12810 14118
rect 12834 14116 12890 14118
rect 12914 14116 12970 14118
rect 12994 14116 13050 14118
rect 12754 13082 12810 13084
rect 12834 13082 12890 13084
rect 12914 13082 12970 13084
rect 12994 13082 13050 13084
rect 12754 13030 12800 13082
rect 12800 13030 12810 13082
rect 12834 13030 12864 13082
rect 12864 13030 12876 13082
rect 12876 13030 12890 13082
rect 12914 13030 12928 13082
rect 12928 13030 12940 13082
rect 12940 13030 12970 13082
rect 12994 13030 13004 13082
rect 13004 13030 13050 13082
rect 12754 13028 12810 13030
rect 12834 13028 12890 13030
rect 12914 13028 12970 13030
rect 12994 13028 13050 13030
rect 12754 11994 12810 11996
rect 12834 11994 12890 11996
rect 12914 11994 12970 11996
rect 12994 11994 13050 11996
rect 12754 11942 12800 11994
rect 12800 11942 12810 11994
rect 12834 11942 12864 11994
rect 12864 11942 12876 11994
rect 12876 11942 12890 11994
rect 12914 11942 12928 11994
rect 12928 11942 12940 11994
rect 12940 11942 12970 11994
rect 12994 11942 13004 11994
rect 13004 11942 13050 11994
rect 12754 11940 12810 11942
rect 12834 11940 12890 11942
rect 12914 11940 12970 11942
rect 12994 11940 13050 11942
rect 12754 10906 12810 10908
rect 12834 10906 12890 10908
rect 12914 10906 12970 10908
rect 12994 10906 13050 10908
rect 12754 10854 12800 10906
rect 12800 10854 12810 10906
rect 12834 10854 12864 10906
rect 12864 10854 12876 10906
rect 12876 10854 12890 10906
rect 12914 10854 12928 10906
rect 12928 10854 12940 10906
rect 12940 10854 12970 10906
rect 12994 10854 13004 10906
rect 13004 10854 13050 10906
rect 12754 10852 12810 10854
rect 12834 10852 12890 10854
rect 12914 10852 12970 10854
rect 12994 10852 13050 10854
rect 12754 9818 12810 9820
rect 12834 9818 12890 9820
rect 12914 9818 12970 9820
rect 12994 9818 13050 9820
rect 12754 9766 12800 9818
rect 12800 9766 12810 9818
rect 12834 9766 12864 9818
rect 12864 9766 12876 9818
rect 12876 9766 12890 9818
rect 12914 9766 12928 9818
rect 12928 9766 12940 9818
rect 12940 9766 12970 9818
rect 12994 9766 13004 9818
rect 13004 9766 13050 9818
rect 12754 9764 12810 9766
rect 12834 9764 12890 9766
rect 12914 9764 12970 9766
rect 12994 9764 13050 9766
rect 13174 9596 13176 9616
rect 13176 9596 13228 9616
rect 13228 9596 13230 9616
rect 10788 6010 10844 6012
rect 10868 6010 10924 6012
rect 10948 6010 11004 6012
rect 11028 6010 11084 6012
rect 10788 5958 10834 6010
rect 10834 5958 10844 6010
rect 10868 5958 10898 6010
rect 10898 5958 10910 6010
rect 10910 5958 10924 6010
rect 10948 5958 10962 6010
rect 10962 5958 10974 6010
rect 10974 5958 11004 6010
rect 11028 5958 11038 6010
rect 11038 5958 11084 6010
rect 10788 5956 10844 5958
rect 10868 5956 10924 5958
rect 10948 5956 11004 5958
rect 11028 5956 11084 5958
rect 11242 5480 11298 5536
rect 10788 4922 10844 4924
rect 10868 4922 10924 4924
rect 10948 4922 11004 4924
rect 11028 4922 11084 4924
rect 10788 4870 10834 4922
rect 10834 4870 10844 4922
rect 10868 4870 10898 4922
rect 10898 4870 10910 4922
rect 10910 4870 10924 4922
rect 10948 4870 10962 4922
rect 10962 4870 10974 4922
rect 10974 4870 11004 4922
rect 11028 4870 11038 4922
rect 11038 4870 11084 4922
rect 10788 4868 10844 4870
rect 10868 4868 10924 4870
rect 10948 4868 11004 4870
rect 11028 4868 11084 4870
rect 9402 2488 9458 2544
rect 938 1944 994 2000
rect 4888 2202 4944 2204
rect 4968 2202 5024 2204
rect 5048 2202 5104 2204
rect 5128 2202 5184 2204
rect 4888 2150 4934 2202
rect 4934 2150 4944 2202
rect 4968 2150 4998 2202
rect 4998 2150 5010 2202
rect 5010 2150 5024 2202
rect 5048 2150 5062 2202
rect 5062 2150 5074 2202
rect 5074 2150 5104 2202
rect 5128 2150 5138 2202
rect 5138 2150 5184 2202
rect 4888 2148 4944 2150
rect 4968 2148 5024 2150
rect 5048 2148 5104 2150
rect 5128 2148 5184 2150
rect 10788 3834 10844 3836
rect 10868 3834 10924 3836
rect 10948 3834 11004 3836
rect 11028 3834 11084 3836
rect 10788 3782 10834 3834
rect 10834 3782 10844 3834
rect 10868 3782 10898 3834
rect 10898 3782 10910 3834
rect 10910 3782 10924 3834
rect 10948 3782 10962 3834
rect 10962 3782 10974 3834
rect 10974 3782 11004 3834
rect 11028 3782 11038 3834
rect 11038 3782 11084 3834
rect 10788 3780 10844 3782
rect 10868 3780 10924 3782
rect 10948 3780 11004 3782
rect 11028 3780 11084 3782
rect 12754 8730 12810 8732
rect 12834 8730 12890 8732
rect 12914 8730 12970 8732
rect 12994 8730 13050 8732
rect 12754 8678 12800 8730
rect 12800 8678 12810 8730
rect 12834 8678 12864 8730
rect 12864 8678 12876 8730
rect 12876 8678 12890 8730
rect 12914 8678 12928 8730
rect 12928 8678 12940 8730
rect 12940 8678 12970 8730
rect 12994 8678 13004 8730
rect 13004 8678 13050 8730
rect 12754 8676 12810 8678
rect 12834 8676 12890 8678
rect 12914 8676 12970 8678
rect 12994 8676 13050 8678
rect 13174 9560 13230 9596
rect 12898 7828 12900 7848
rect 12900 7828 12952 7848
rect 12952 7828 12954 7848
rect 12898 7792 12954 7828
rect 12754 7642 12810 7644
rect 12834 7642 12890 7644
rect 12914 7642 12970 7644
rect 12994 7642 13050 7644
rect 12754 7590 12800 7642
rect 12800 7590 12810 7642
rect 12834 7590 12864 7642
rect 12864 7590 12876 7642
rect 12876 7590 12890 7642
rect 12914 7590 12928 7642
rect 12928 7590 12940 7642
rect 12940 7590 12970 7642
rect 12994 7590 13004 7642
rect 13004 7590 13050 7642
rect 12754 7588 12810 7590
rect 12834 7588 12890 7590
rect 12914 7588 12970 7590
rect 12994 7588 13050 7590
rect 12754 6554 12810 6556
rect 12834 6554 12890 6556
rect 12914 6554 12970 6556
rect 12994 6554 13050 6556
rect 12754 6502 12800 6554
rect 12800 6502 12810 6554
rect 12834 6502 12864 6554
rect 12864 6502 12876 6554
rect 12876 6502 12890 6554
rect 12914 6502 12928 6554
rect 12928 6502 12940 6554
rect 12940 6502 12970 6554
rect 12994 6502 13004 6554
rect 13004 6502 13050 6554
rect 12754 6500 12810 6502
rect 12834 6500 12890 6502
rect 12914 6500 12970 6502
rect 12994 6500 13050 6502
rect 14721 14714 14777 14716
rect 14801 14714 14857 14716
rect 14881 14714 14937 14716
rect 14961 14714 15017 14716
rect 14721 14662 14767 14714
rect 14767 14662 14777 14714
rect 14801 14662 14831 14714
rect 14831 14662 14843 14714
rect 14843 14662 14857 14714
rect 14881 14662 14895 14714
rect 14895 14662 14907 14714
rect 14907 14662 14937 14714
rect 14961 14662 14971 14714
rect 14971 14662 15017 14714
rect 14721 14660 14777 14662
rect 14801 14660 14857 14662
rect 14881 14660 14937 14662
rect 14961 14660 15017 14662
rect 15566 15000 15622 15056
rect 16670 15816 16726 15872
rect 16687 15258 16743 15260
rect 16767 15258 16823 15260
rect 16847 15258 16903 15260
rect 16927 15258 16983 15260
rect 16687 15206 16733 15258
rect 16733 15206 16743 15258
rect 16767 15206 16797 15258
rect 16797 15206 16809 15258
rect 16809 15206 16823 15258
rect 16847 15206 16861 15258
rect 16861 15206 16873 15258
rect 16873 15206 16903 15258
rect 16927 15206 16937 15258
rect 16937 15206 16983 15258
rect 16687 15204 16743 15206
rect 16767 15204 16823 15206
rect 16847 15204 16903 15206
rect 16927 15204 16983 15206
rect 14721 13626 14777 13628
rect 14801 13626 14857 13628
rect 14881 13626 14937 13628
rect 14961 13626 15017 13628
rect 14721 13574 14767 13626
rect 14767 13574 14777 13626
rect 14801 13574 14831 13626
rect 14831 13574 14843 13626
rect 14843 13574 14857 13626
rect 14881 13574 14895 13626
rect 14895 13574 14907 13626
rect 14907 13574 14937 13626
rect 14961 13574 14971 13626
rect 14971 13574 15017 13626
rect 14721 13572 14777 13574
rect 14801 13572 14857 13574
rect 14881 13572 14937 13574
rect 14961 13572 15017 13574
rect 14721 12538 14777 12540
rect 14801 12538 14857 12540
rect 14881 12538 14937 12540
rect 14961 12538 15017 12540
rect 14721 12486 14767 12538
rect 14767 12486 14777 12538
rect 14801 12486 14831 12538
rect 14831 12486 14843 12538
rect 14843 12486 14857 12538
rect 14881 12486 14895 12538
rect 14895 12486 14907 12538
rect 14907 12486 14937 12538
rect 14961 12486 14971 12538
rect 14971 12486 15017 12538
rect 14721 12484 14777 12486
rect 14801 12484 14857 12486
rect 14881 12484 14937 12486
rect 14961 12484 15017 12486
rect 15106 11736 15162 11792
rect 14721 11450 14777 11452
rect 14801 11450 14857 11452
rect 14881 11450 14937 11452
rect 14961 11450 15017 11452
rect 14721 11398 14767 11450
rect 14767 11398 14777 11450
rect 14801 11398 14831 11450
rect 14831 11398 14843 11450
rect 14843 11398 14857 11450
rect 14881 11398 14895 11450
rect 14895 11398 14907 11450
rect 14907 11398 14937 11450
rect 14961 11398 14971 11450
rect 14971 11398 15017 11450
rect 14721 11396 14777 11398
rect 14801 11396 14857 11398
rect 14881 11396 14937 11398
rect 14961 11396 15017 11398
rect 14186 11076 14242 11112
rect 14186 11056 14188 11076
rect 14188 11056 14240 11076
rect 14240 11056 14242 11076
rect 14554 11076 14610 11112
rect 14554 11056 14556 11076
rect 14556 11056 14608 11076
rect 14608 11056 14610 11076
rect 16486 14340 16542 14376
rect 16486 14320 16488 14340
rect 16488 14320 16540 14340
rect 16540 14320 16542 14340
rect 16687 14170 16743 14172
rect 16767 14170 16823 14172
rect 16847 14170 16903 14172
rect 16927 14170 16983 14172
rect 16687 14118 16733 14170
rect 16733 14118 16743 14170
rect 16767 14118 16797 14170
rect 16797 14118 16809 14170
rect 16809 14118 16823 14170
rect 16847 14118 16861 14170
rect 16861 14118 16873 14170
rect 16873 14118 16903 14170
rect 16927 14118 16937 14170
rect 16937 14118 16983 14170
rect 16687 14116 16743 14118
rect 16767 14116 16823 14118
rect 16847 14116 16903 14118
rect 16927 14116 16983 14118
rect 14830 10548 14832 10568
rect 14832 10548 14884 10568
rect 14884 10548 14886 10568
rect 14830 10512 14886 10548
rect 14721 10362 14777 10364
rect 14801 10362 14857 10364
rect 14881 10362 14937 10364
rect 14961 10362 15017 10364
rect 14721 10310 14767 10362
rect 14767 10310 14777 10362
rect 14801 10310 14831 10362
rect 14831 10310 14843 10362
rect 14843 10310 14857 10362
rect 14881 10310 14895 10362
rect 14895 10310 14907 10362
rect 14907 10310 14937 10362
rect 14961 10310 14971 10362
rect 14971 10310 15017 10362
rect 14721 10308 14777 10310
rect 14801 10308 14857 10310
rect 14881 10308 14937 10310
rect 14961 10308 15017 10310
rect 14094 9560 14150 9616
rect 16302 10104 16358 10160
rect 14646 10004 14648 10024
rect 14648 10004 14700 10024
rect 14700 10004 14702 10024
rect 14646 9968 14702 10004
rect 14721 9274 14777 9276
rect 14801 9274 14857 9276
rect 14881 9274 14937 9276
rect 14961 9274 15017 9276
rect 14721 9222 14767 9274
rect 14767 9222 14777 9274
rect 14801 9222 14831 9274
rect 14831 9222 14843 9274
rect 14843 9222 14857 9274
rect 14881 9222 14895 9274
rect 14895 9222 14907 9274
rect 14907 9222 14937 9274
rect 14961 9222 14971 9274
rect 14971 9222 15017 9274
rect 14721 9220 14777 9222
rect 14801 9220 14857 9222
rect 14881 9220 14937 9222
rect 14961 9220 15017 9222
rect 15106 8472 15162 8528
rect 14721 8186 14777 8188
rect 14801 8186 14857 8188
rect 14881 8186 14937 8188
rect 14961 8186 15017 8188
rect 14721 8134 14767 8186
rect 14767 8134 14777 8186
rect 14801 8134 14831 8186
rect 14831 8134 14843 8186
rect 14843 8134 14857 8186
rect 14881 8134 14895 8186
rect 14895 8134 14907 8186
rect 14907 8134 14937 8186
rect 14961 8134 14971 8186
rect 14971 8134 15017 8186
rect 14721 8132 14777 8134
rect 14801 8132 14857 8134
rect 14881 8132 14937 8134
rect 14961 8132 15017 8134
rect 14186 7792 14242 7848
rect 12754 5466 12810 5468
rect 12834 5466 12890 5468
rect 12914 5466 12970 5468
rect 12994 5466 13050 5468
rect 12754 5414 12800 5466
rect 12800 5414 12810 5466
rect 12834 5414 12864 5466
rect 12864 5414 12876 5466
rect 12876 5414 12890 5466
rect 12914 5414 12928 5466
rect 12928 5414 12940 5466
rect 12940 5414 12970 5466
rect 12994 5414 13004 5466
rect 13004 5414 13050 5466
rect 12754 5412 12810 5414
rect 12834 5412 12890 5414
rect 12914 5412 12970 5414
rect 12994 5412 13050 5414
rect 10788 2746 10844 2748
rect 10868 2746 10924 2748
rect 10948 2746 11004 2748
rect 11028 2746 11084 2748
rect 10788 2694 10834 2746
rect 10834 2694 10844 2746
rect 10868 2694 10898 2746
rect 10898 2694 10910 2746
rect 10910 2694 10924 2746
rect 10948 2694 10962 2746
rect 10962 2694 10974 2746
rect 10974 2694 11004 2746
rect 11028 2694 11038 2746
rect 11038 2694 11084 2746
rect 10788 2692 10844 2694
rect 10868 2692 10924 2694
rect 10948 2692 11004 2694
rect 11028 2692 11084 2694
rect 11426 2644 11482 2680
rect 11426 2624 11428 2644
rect 11428 2624 11480 2644
rect 11480 2624 11482 2644
rect 8821 2202 8877 2204
rect 8901 2202 8957 2204
rect 8981 2202 9037 2204
rect 9061 2202 9117 2204
rect 8821 2150 8867 2202
rect 8867 2150 8877 2202
rect 8901 2150 8931 2202
rect 8931 2150 8943 2202
rect 8943 2150 8957 2202
rect 8981 2150 8995 2202
rect 8995 2150 9007 2202
rect 9007 2150 9037 2202
rect 9061 2150 9071 2202
rect 9071 2150 9117 2202
rect 8821 2148 8877 2150
rect 8901 2148 8957 2150
rect 8981 2148 9037 2150
rect 9061 2148 9117 2150
rect 11886 2488 11942 2544
rect 12438 4528 12494 4584
rect 12754 4378 12810 4380
rect 12834 4378 12890 4380
rect 12914 4378 12970 4380
rect 12994 4378 13050 4380
rect 12754 4326 12800 4378
rect 12800 4326 12810 4378
rect 12834 4326 12864 4378
rect 12864 4326 12876 4378
rect 12876 4326 12890 4378
rect 12914 4326 12928 4378
rect 12928 4326 12940 4378
rect 12940 4326 12970 4378
rect 12994 4326 13004 4378
rect 13004 4326 13050 4378
rect 12754 4324 12810 4326
rect 12834 4324 12890 4326
rect 12914 4324 12970 4326
rect 12994 4324 13050 4326
rect 12754 3290 12810 3292
rect 12834 3290 12890 3292
rect 12914 3290 12970 3292
rect 12994 3290 13050 3292
rect 12754 3238 12800 3290
rect 12800 3238 12810 3290
rect 12834 3238 12864 3290
rect 12864 3238 12876 3290
rect 12876 3238 12890 3290
rect 12914 3238 12928 3290
rect 12928 3238 12940 3290
rect 12940 3238 12970 3290
rect 12994 3238 13004 3290
rect 13004 3238 13050 3290
rect 12754 3236 12810 3238
rect 12834 3236 12890 3238
rect 12914 3236 12970 3238
rect 12994 3236 13050 3238
rect 13634 6432 13690 6488
rect 14721 7098 14777 7100
rect 14801 7098 14857 7100
rect 14881 7098 14937 7100
rect 14961 7098 15017 7100
rect 14721 7046 14767 7098
rect 14767 7046 14777 7098
rect 14801 7046 14831 7098
rect 14831 7046 14843 7098
rect 14843 7046 14857 7098
rect 14881 7046 14895 7098
rect 14895 7046 14907 7098
rect 14907 7046 14937 7098
rect 14961 7046 14971 7098
rect 14971 7046 15017 7098
rect 14721 7044 14777 7046
rect 14801 7044 14857 7046
rect 14881 7044 14937 7046
rect 14961 7044 15017 7046
rect 14830 6860 14886 6896
rect 14830 6840 14832 6860
rect 14832 6840 14884 6860
rect 14884 6840 14886 6860
rect 13818 5208 13874 5264
rect 14830 6160 14886 6216
rect 13910 3984 13966 4040
rect 14721 6010 14777 6012
rect 14801 6010 14857 6012
rect 14881 6010 14937 6012
rect 14961 6010 15017 6012
rect 14721 5958 14767 6010
rect 14767 5958 14777 6010
rect 14801 5958 14831 6010
rect 14831 5958 14843 6010
rect 14843 5958 14857 6010
rect 14881 5958 14895 6010
rect 14895 5958 14907 6010
rect 14907 5958 14937 6010
rect 14961 5958 14971 6010
rect 14971 5958 15017 6010
rect 14721 5956 14777 5958
rect 14801 5956 14857 5958
rect 14881 5956 14937 5958
rect 14961 5956 15017 5958
rect 14721 4922 14777 4924
rect 14801 4922 14857 4924
rect 14881 4922 14937 4924
rect 14961 4922 15017 4924
rect 14721 4870 14767 4922
rect 14767 4870 14777 4922
rect 14801 4870 14831 4922
rect 14831 4870 14843 4922
rect 14843 4870 14857 4922
rect 14881 4870 14895 4922
rect 14895 4870 14907 4922
rect 14907 4870 14937 4922
rect 14961 4870 14971 4922
rect 14971 4870 15017 4922
rect 14721 4868 14777 4870
rect 14801 4868 14857 4870
rect 14881 4868 14937 4870
rect 14961 4868 15017 4870
rect 14721 3834 14777 3836
rect 14801 3834 14857 3836
rect 14881 3834 14937 3836
rect 14961 3834 15017 3836
rect 14721 3782 14767 3834
rect 14767 3782 14777 3834
rect 14801 3782 14831 3834
rect 14831 3782 14843 3834
rect 14843 3782 14857 3834
rect 14881 3782 14895 3834
rect 14895 3782 14907 3834
rect 14907 3782 14937 3834
rect 14961 3782 14971 3834
rect 14971 3782 15017 3834
rect 14721 3780 14777 3782
rect 14801 3780 14857 3782
rect 14881 3780 14937 3782
rect 14961 3780 15017 3782
rect 14370 3576 14426 3632
rect 16210 9696 16266 9752
rect 16486 13368 16542 13424
rect 16687 13082 16743 13084
rect 16767 13082 16823 13084
rect 16847 13082 16903 13084
rect 16927 13082 16983 13084
rect 16687 13030 16733 13082
rect 16733 13030 16743 13082
rect 16767 13030 16797 13082
rect 16797 13030 16809 13082
rect 16809 13030 16823 13082
rect 16847 13030 16861 13082
rect 16861 13030 16873 13082
rect 16873 13030 16903 13082
rect 16927 13030 16937 13082
rect 16937 13030 16983 13082
rect 16687 13028 16743 13030
rect 16767 13028 16823 13030
rect 16847 13028 16903 13030
rect 16927 13028 16983 13030
rect 16762 12552 16818 12608
rect 16687 11994 16743 11996
rect 16767 11994 16823 11996
rect 16847 11994 16903 11996
rect 16927 11994 16983 11996
rect 16687 11942 16733 11994
rect 16733 11942 16743 11994
rect 16767 11942 16797 11994
rect 16797 11942 16809 11994
rect 16809 11942 16823 11994
rect 16847 11942 16861 11994
rect 16861 11942 16873 11994
rect 16873 11942 16903 11994
rect 16927 11942 16937 11994
rect 16937 11942 16983 11994
rect 16687 11940 16743 11942
rect 16767 11940 16823 11942
rect 16847 11940 16903 11942
rect 16927 11940 16983 11942
rect 16687 10906 16743 10908
rect 16767 10906 16823 10908
rect 16847 10906 16903 10908
rect 16927 10906 16983 10908
rect 16687 10854 16733 10906
rect 16733 10854 16743 10906
rect 16767 10854 16797 10906
rect 16797 10854 16809 10906
rect 16809 10854 16823 10906
rect 16847 10854 16861 10906
rect 16861 10854 16873 10906
rect 16873 10854 16903 10906
rect 16927 10854 16937 10906
rect 16937 10854 16983 10906
rect 16687 10852 16743 10854
rect 16767 10852 16823 10854
rect 16847 10852 16903 10854
rect 16927 10852 16983 10854
rect 16486 10104 16542 10160
rect 16687 9818 16743 9820
rect 16767 9818 16823 9820
rect 16847 9818 16903 9820
rect 16927 9818 16983 9820
rect 16687 9766 16733 9818
rect 16733 9766 16743 9818
rect 16767 9766 16797 9818
rect 16797 9766 16809 9818
rect 16809 9766 16823 9818
rect 16847 9766 16861 9818
rect 16861 9766 16873 9818
rect 16873 9766 16903 9818
rect 16927 9766 16937 9818
rect 16937 9766 16983 9818
rect 16687 9764 16743 9766
rect 16767 9764 16823 9766
rect 16847 9764 16903 9766
rect 16927 9764 16983 9766
rect 16762 9288 16818 9344
rect 16687 8730 16743 8732
rect 16767 8730 16823 8732
rect 16847 8730 16903 8732
rect 16927 8730 16983 8732
rect 16687 8678 16733 8730
rect 16733 8678 16743 8730
rect 16767 8678 16797 8730
rect 16797 8678 16809 8730
rect 16809 8678 16823 8730
rect 16847 8678 16861 8730
rect 16861 8678 16873 8730
rect 16873 8678 16903 8730
rect 16927 8678 16937 8730
rect 16937 8678 16983 8730
rect 16687 8676 16743 8678
rect 16767 8676 16823 8678
rect 16847 8676 16903 8678
rect 16927 8676 16983 8678
rect 15750 6432 15806 6488
rect 15842 6296 15898 6352
rect 15842 6160 15898 6216
rect 14721 2746 14777 2748
rect 14801 2746 14857 2748
rect 14881 2746 14937 2748
rect 14961 2746 15017 2748
rect 14721 2694 14767 2746
rect 14767 2694 14777 2746
rect 14801 2694 14831 2746
rect 14831 2694 14843 2746
rect 14843 2694 14857 2746
rect 14881 2694 14895 2746
rect 14895 2694 14907 2746
rect 14907 2694 14937 2746
rect 14961 2694 14971 2746
rect 14971 2694 15017 2746
rect 14721 2692 14777 2694
rect 14801 2692 14857 2694
rect 14881 2692 14937 2694
rect 14961 2692 15017 2694
rect 15658 2760 15714 2816
rect 16486 7792 16542 7848
rect 16687 7642 16743 7644
rect 16767 7642 16823 7644
rect 16847 7642 16903 7644
rect 16927 7642 16983 7644
rect 16687 7590 16733 7642
rect 16733 7590 16743 7642
rect 16767 7590 16797 7642
rect 16797 7590 16809 7642
rect 16809 7590 16823 7642
rect 16847 7590 16861 7642
rect 16861 7590 16873 7642
rect 16873 7590 16903 7642
rect 16927 7590 16937 7642
rect 16937 7590 16983 7642
rect 16687 7588 16743 7590
rect 16767 7588 16823 7590
rect 16847 7588 16903 7590
rect 16927 7588 16983 7590
rect 16578 6840 16634 6896
rect 16687 6554 16743 6556
rect 16767 6554 16823 6556
rect 16847 6554 16903 6556
rect 16927 6554 16983 6556
rect 16687 6502 16733 6554
rect 16733 6502 16743 6554
rect 16767 6502 16797 6554
rect 16797 6502 16809 6554
rect 16809 6502 16823 6554
rect 16847 6502 16861 6554
rect 16861 6502 16873 6554
rect 16873 6502 16903 6554
rect 16927 6502 16937 6554
rect 16937 6502 16983 6554
rect 16687 6500 16743 6502
rect 16767 6500 16823 6502
rect 16847 6500 16903 6502
rect 16927 6500 16983 6502
rect 16687 5466 16743 5468
rect 16767 5466 16823 5468
rect 16847 5466 16903 5468
rect 16927 5466 16983 5468
rect 16687 5414 16733 5466
rect 16733 5414 16743 5466
rect 16767 5414 16797 5466
rect 16797 5414 16809 5466
rect 16809 5414 16823 5466
rect 16847 5414 16861 5466
rect 16861 5414 16873 5466
rect 16873 5414 16903 5466
rect 16927 5414 16937 5466
rect 16937 5414 16983 5466
rect 16687 5412 16743 5414
rect 16767 5412 16823 5414
rect 16847 5412 16903 5414
rect 16927 5412 16983 5414
rect 16687 4378 16743 4380
rect 16767 4378 16823 4380
rect 16847 4378 16903 4380
rect 16927 4378 16983 4380
rect 16687 4326 16733 4378
rect 16733 4326 16743 4378
rect 16767 4326 16797 4378
rect 16797 4326 16809 4378
rect 16809 4326 16823 4378
rect 16847 4326 16861 4378
rect 16861 4326 16873 4378
rect 16873 4326 16903 4378
rect 16927 4326 16937 4378
rect 16937 4326 16983 4378
rect 16687 4324 16743 4326
rect 16767 4324 16823 4326
rect 16847 4324 16903 4326
rect 16927 4324 16983 4326
rect 16302 3984 16358 4040
rect 16687 3290 16743 3292
rect 16767 3290 16823 3292
rect 16847 3290 16903 3292
rect 16927 3290 16983 3292
rect 16687 3238 16733 3290
rect 16733 3238 16743 3290
rect 16767 3238 16797 3290
rect 16797 3238 16809 3290
rect 16809 3238 16823 3290
rect 16847 3238 16861 3290
rect 16861 3238 16873 3290
rect 16873 3238 16903 3290
rect 16927 3238 16937 3290
rect 16937 3238 16983 3290
rect 16687 3236 16743 3238
rect 16767 3236 16823 3238
rect 16847 3236 16903 3238
rect 16927 3236 16983 3238
rect 12754 2202 12810 2204
rect 12834 2202 12890 2204
rect 12914 2202 12970 2204
rect 12994 2202 13050 2204
rect 12754 2150 12800 2202
rect 12800 2150 12810 2202
rect 12834 2150 12864 2202
rect 12864 2150 12876 2202
rect 12876 2150 12890 2202
rect 12914 2150 12928 2202
rect 12928 2150 12940 2202
rect 12940 2150 12970 2202
rect 12994 2150 13004 2202
rect 13004 2150 13050 2202
rect 12754 2148 12810 2150
rect 12834 2148 12890 2150
rect 12914 2148 12970 2150
rect 12994 2148 13050 2150
rect 13818 312 13874 368
rect 16687 2202 16743 2204
rect 16767 2202 16823 2204
rect 16847 2202 16903 2204
rect 16927 2202 16983 2204
rect 16687 2150 16733 2202
rect 16733 2150 16743 2202
rect 16767 2150 16797 2202
rect 16797 2150 16809 2202
rect 16809 2150 16823 2202
rect 16847 2150 16861 2202
rect 16861 2150 16873 2202
rect 16873 2150 16903 2202
rect 16927 2150 16937 2202
rect 16937 2150 16983 2202
rect 16687 2148 16743 2150
rect 16767 2148 16823 2150
rect 16847 2148 16903 2150
rect 16927 2148 16983 2150
rect 16578 1944 16634 2000
rect 16302 1128 16358 1184
<< metal3 >>
rect 14917 17506 14983 17509
rect 17200 17506 18000 17536
rect 14917 17504 18000 17506
rect 14917 17448 14922 17504
rect 14978 17448 18000 17504
rect 14917 17446 18000 17448
rect 14917 17443 14983 17446
rect 17200 17416 18000 17446
rect 0 16690 800 16720
rect 1485 16690 1551 16693
rect 0 16688 1551 16690
rect 0 16632 1490 16688
rect 1546 16632 1551 16688
rect 0 16630 1551 16632
rect 0 16600 800 16630
rect 1485 16627 1551 16630
rect 16481 16690 16547 16693
rect 17200 16690 18000 16720
rect 16481 16688 18000 16690
rect 16481 16632 16486 16688
rect 16542 16632 18000 16688
rect 16481 16630 18000 16632
rect 16481 16627 16547 16630
rect 17200 16600 18000 16630
rect 0 15874 800 15904
rect 933 15874 999 15877
rect 0 15872 999 15874
rect 0 15816 938 15872
rect 994 15816 999 15872
rect 0 15814 999 15816
rect 0 15784 800 15814
rect 933 15811 999 15814
rect 16665 15874 16731 15877
rect 17200 15874 18000 15904
rect 16665 15872 18000 15874
rect 16665 15816 16670 15872
rect 16726 15816 18000 15872
rect 16665 15814 18000 15816
rect 16665 15811 16731 15814
rect 2912 15808 3228 15809
rect 2912 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3228 15808
rect 2912 15743 3228 15744
rect 6845 15808 7161 15809
rect 6845 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7161 15808
rect 6845 15743 7161 15744
rect 10778 15808 11094 15809
rect 10778 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11094 15808
rect 10778 15743 11094 15744
rect 14711 15808 15027 15809
rect 14711 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15027 15808
rect 17200 15784 18000 15814
rect 14711 15743 15027 15744
rect 4878 15264 5194 15265
rect 4878 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5194 15264
rect 4878 15199 5194 15200
rect 8811 15264 9127 15265
rect 8811 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9127 15264
rect 8811 15199 9127 15200
rect 12744 15264 13060 15265
rect 12744 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13060 15264
rect 12744 15199 13060 15200
rect 16677 15264 16993 15265
rect 16677 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16993 15264
rect 16677 15199 16993 15200
rect 2221 15194 2287 15197
rect 1166 15192 2287 15194
rect 1166 15136 2226 15192
rect 2282 15136 2287 15192
rect 1166 15134 2287 15136
rect 0 15058 800 15088
rect 1166 15058 1226 15134
rect 2221 15131 2287 15134
rect 0 14998 1226 15058
rect 15561 15058 15627 15061
rect 17200 15058 18000 15088
rect 15561 15056 18000 15058
rect 15561 15000 15566 15056
rect 15622 15000 18000 15056
rect 15561 14998 18000 15000
rect 0 14968 800 14998
rect 15561 14995 15627 14998
rect 17200 14968 18000 14998
rect 2912 14720 3228 14721
rect 2912 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3228 14720
rect 2912 14655 3228 14656
rect 6845 14720 7161 14721
rect 6845 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7161 14720
rect 6845 14655 7161 14656
rect 10778 14720 11094 14721
rect 10778 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11094 14720
rect 10778 14655 11094 14656
rect 14711 14720 15027 14721
rect 14711 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15027 14720
rect 14711 14655 15027 14656
rect 16481 14378 16547 14381
rect 16481 14376 17188 14378
rect 16481 14320 16486 14376
rect 16542 14320 17188 14376
rect 16481 14318 17188 14320
rect 16481 14315 16547 14318
rect 17128 14276 17188 14318
rect 17128 14272 17418 14276
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 17128 14216 18000 14272
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 4878 14176 5194 14177
rect 4878 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5194 14176
rect 4878 14111 5194 14112
rect 8811 14176 9127 14177
rect 8811 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9127 14176
rect 8811 14111 9127 14112
rect 12744 14176 13060 14177
rect 12744 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13060 14176
rect 12744 14111 13060 14112
rect 16677 14176 16993 14177
rect 16677 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16993 14176
rect 17200 14152 18000 14216
rect 16677 14111 16993 14112
rect 1485 13696 1551 13701
rect 1485 13640 1490 13696
rect 1546 13640 1551 13696
rect 1485 13635 1551 13640
rect 0 13426 800 13456
rect 1488 13426 1548 13635
rect 2912 13632 3228 13633
rect 2912 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3228 13632
rect 2912 13567 3228 13568
rect 6845 13632 7161 13633
rect 6845 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7161 13632
rect 6845 13567 7161 13568
rect 10778 13632 11094 13633
rect 10778 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11094 13632
rect 10778 13567 11094 13568
rect 14711 13632 15027 13633
rect 14711 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15027 13632
rect 14711 13567 15027 13568
rect 0 13366 1548 13426
rect 16481 13426 16547 13429
rect 17200 13426 18000 13456
rect 16481 13424 18000 13426
rect 16481 13368 16486 13424
rect 16542 13368 18000 13424
rect 16481 13366 18000 13368
rect 0 13336 800 13366
rect 16481 13363 16547 13366
rect 17200 13336 18000 13366
rect 4878 13088 5194 13089
rect 4878 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5194 13088
rect 4878 13023 5194 13024
rect 8811 13088 9127 13089
rect 8811 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9127 13088
rect 8811 13023 9127 13024
rect 12744 13088 13060 13089
rect 12744 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13060 13088
rect 12744 13023 13060 13024
rect 16677 13088 16993 13089
rect 16677 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16993 13088
rect 16677 13023 16993 13024
rect 0 12610 800 12640
rect 933 12610 999 12613
rect 0 12608 999 12610
rect 0 12552 938 12608
rect 994 12552 999 12608
rect 0 12550 999 12552
rect 0 12520 800 12550
rect 933 12547 999 12550
rect 16757 12610 16823 12613
rect 17200 12610 18000 12640
rect 16757 12608 18000 12610
rect 16757 12552 16762 12608
rect 16818 12552 18000 12608
rect 16757 12550 18000 12552
rect 16757 12547 16823 12550
rect 2912 12544 3228 12545
rect 2912 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3228 12544
rect 2912 12479 3228 12480
rect 6845 12544 7161 12545
rect 6845 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7161 12544
rect 6845 12479 7161 12480
rect 10778 12544 11094 12545
rect 10778 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11094 12544
rect 10778 12479 11094 12480
rect 14711 12544 15027 12545
rect 14711 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15027 12544
rect 17200 12520 18000 12550
rect 14711 12479 15027 12480
rect 4878 12000 5194 12001
rect 4878 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5194 12000
rect 4878 11935 5194 11936
rect 8811 12000 9127 12001
rect 8811 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9127 12000
rect 8811 11935 9127 11936
rect 12744 12000 13060 12001
rect 12744 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13060 12000
rect 12744 11935 13060 11936
rect 16677 12000 16993 12001
rect 16677 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16993 12000
rect 16677 11935 16993 11936
rect 0 11794 800 11824
rect 933 11794 999 11797
rect 0 11792 999 11794
rect 0 11736 938 11792
rect 994 11736 999 11792
rect 0 11734 999 11736
rect 0 11704 800 11734
rect 933 11731 999 11734
rect 15101 11794 15167 11797
rect 17200 11794 18000 11824
rect 15101 11792 18000 11794
rect 15101 11736 15106 11792
rect 15162 11736 18000 11792
rect 15101 11734 18000 11736
rect 15101 11731 15167 11734
rect 17200 11704 18000 11734
rect 2912 11456 3228 11457
rect 2912 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3228 11456
rect 2912 11391 3228 11392
rect 6845 11456 7161 11457
rect 6845 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7161 11456
rect 6845 11391 7161 11392
rect 10778 11456 11094 11457
rect 10778 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11094 11456
rect 10778 11391 11094 11392
rect 14711 11456 15027 11457
rect 14711 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15027 11456
rect 14711 11391 15027 11392
rect 11278 11052 11284 11116
rect 11348 11114 11354 11116
rect 11513 11114 11579 11117
rect 11348 11112 11579 11114
rect 11348 11056 11518 11112
rect 11574 11056 11579 11112
rect 11348 11054 11579 11056
rect 11348 11052 11354 11054
rect 11513 11051 11579 11054
rect 14181 11116 14247 11117
rect 14181 11112 14228 11116
rect 14292 11114 14298 11116
rect 14549 11114 14615 11117
rect 14181 11056 14186 11112
rect 14181 11052 14228 11056
rect 14292 11054 14338 11114
rect 14549 11112 17188 11114
rect 14549 11056 14554 11112
rect 14610 11056 17188 11112
rect 14549 11054 17188 11056
rect 14292 11052 14298 11054
rect 14181 11051 14247 11052
rect 14549 11051 14615 11054
rect 17128 11012 17188 11054
rect 17128 11008 17418 11012
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 17128 10952 18000 11008
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 4878 10912 5194 10913
rect 4878 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5194 10912
rect 4878 10847 5194 10848
rect 8811 10912 9127 10913
rect 8811 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9127 10912
rect 8811 10847 9127 10848
rect 12744 10912 13060 10913
rect 12744 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13060 10912
rect 12744 10847 13060 10848
rect 16677 10912 16993 10913
rect 16677 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16993 10912
rect 17200 10888 18000 10952
rect 16677 10847 16993 10848
rect 14406 10508 14412 10572
rect 14476 10570 14482 10572
rect 14825 10570 14891 10573
rect 14476 10568 14891 10570
rect 14476 10512 14830 10568
rect 14886 10512 14891 10568
rect 14476 10510 14891 10512
rect 14476 10508 14482 10510
rect 14825 10507 14891 10510
rect 2912 10368 3228 10369
rect 2912 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3228 10368
rect 2912 10303 3228 10304
rect 6845 10368 7161 10369
rect 6845 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7161 10368
rect 6845 10303 7161 10304
rect 10778 10368 11094 10369
rect 10778 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11094 10368
rect 10778 10303 11094 10304
rect 14711 10368 15027 10369
rect 14711 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15027 10368
rect 14711 10303 15027 10304
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 11973 10162 12039 10165
rect 16297 10162 16363 10165
rect 11973 10160 16363 10162
rect 11973 10104 11978 10160
rect 12034 10104 16302 10160
rect 16358 10104 16363 10160
rect 11973 10102 16363 10104
rect 11973 10099 12039 10102
rect 16297 10099 16363 10102
rect 16481 10162 16547 10165
rect 17200 10162 18000 10192
rect 16481 10160 18000 10162
rect 16481 10104 16486 10160
rect 16542 10104 18000 10160
rect 16481 10102 18000 10104
rect 16481 10099 16547 10102
rect 17200 10072 18000 10102
rect 12249 10026 12315 10029
rect 14641 10026 14707 10029
rect 12249 10024 14707 10026
rect 12249 9968 12254 10024
rect 12310 9968 14646 10024
rect 14702 9968 14707 10024
rect 12249 9966 14707 9968
rect 12249 9963 12315 9966
rect 14641 9963 14707 9966
rect 4878 9824 5194 9825
rect 4878 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5194 9824
rect 4878 9759 5194 9760
rect 8811 9824 9127 9825
rect 8811 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9127 9824
rect 8811 9759 9127 9760
rect 12744 9824 13060 9825
rect 12744 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13060 9824
rect 12744 9759 13060 9760
rect 16677 9824 16993 9825
rect 16677 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16993 9824
rect 16677 9759 16993 9760
rect 16205 9756 16271 9757
rect 16205 9752 16252 9756
rect 16316 9754 16322 9756
rect 16205 9696 16210 9752
rect 16205 9692 16252 9696
rect 16316 9694 16362 9754
rect 16316 9692 16322 9694
rect 16205 9691 16271 9692
rect 3325 9618 3391 9621
rect 5441 9618 5507 9621
rect 3325 9616 5507 9618
rect 3325 9560 3330 9616
rect 3386 9560 5446 9616
rect 5502 9560 5507 9616
rect 3325 9558 5507 9560
rect 3325 9555 3391 9558
rect 5441 9555 5507 9558
rect 13169 9618 13235 9621
rect 14089 9618 14155 9621
rect 13169 9616 14155 9618
rect 13169 9560 13174 9616
rect 13230 9560 14094 9616
rect 14150 9560 14155 9616
rect 13169 9558 14155 9560
rect 13169 9555 13235 9558
rect 14089 9555 14155 9558
rect 0 9346 800 9376
rect 16757 9346 16823 9349
rect 17200 9346 18000 9376
rect 0 9286 2698 9346
rect 0 9256 800 9286
rect 2638 9074 2698 9286
rect 16757 9344 18000 9346
rect 16757 9288 16762 9344
rect 16818 9288 18000 9344
rect 16757 9286 18000 9288
rect 16757 9283 16823 9286
rect 2912 9280 3228 9281
rect 2912 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3228 9280
rect 2912 9215 3228 9216
rect 6845 9280 7161 9281
rect 6845 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7161 9280
rect 6845 9215 7161 9216
rect 10778 9280 11094 9281
rect 10778 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11094 9280
rect 10778 9215 11094 9216
rect 14711 9280 15027 9281
rect 14711 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15027 9280
rect 17200 9256 18000 9286
rect 14711 9215 15027 9216
rect 9305 9074 9371 9077
rect 2638 9072 9371 9074
rect 2638 9016 9310 9072
rect 9366 9016 9371 9072
rect 2638 9014 9371 9016
rect 9305 9011 9371 9014
rect 4878 8736 5194 8737
rect 4878 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5194 8736
rect 4878 8671 5194 8672
rect 8811 8736 9127 8737
rect 8811 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9127 8736
rect 8811 8671 9127 8672
rect 12744 8736 13060 8737
rect 12744 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13060 8736
rect 12744 8671 13060 8672
rect 16677 8736 16993 8737
rect 16677 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16993 8736
rect 16677 8671 16993 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 15101 8530 15167 8533
rect 17200 8530 18000 8560
rect 15101 8528 18000 8530
rect 15101 8472 15106 8528
rect 15162 8472 18000 8528
rect 15101 8470 18000 8472
rect 15101 8467 15167 8470
rect 17200 8440 18000 8470
rect 2912 8192 3228 8193
rect 2912 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3228 8192
rect 2912 8127 3228 8128
rect 6845 8192 7161 8193
rect 6845 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7161 8192
rect 6845 8127 7161 8128
rect 10778 8192 11094 8193
rect 10778 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11094 8192
rect 10778 8127 11094 8128
rect 14711 8192 15027 8193
rect 14711 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15027 8192
rect 14711 8127 15027 8128
rect 16530 7926 17188 7986
rect 16530 7853 16590 7926
rect 12893 7850 12959 7853
rect 14181 7850 14247 7853
rect 12893 7848 14247 7850
rect 12893 7792 12898 7848
rect 12954 7792 14186 7848
rect 14242 7792 14247 7848
rect 12893 7790 14247 7792
rect 12893 7787 12959 7790
rect 14181 7787 14247 7790
rect 16481 7848 16590 7853
rect 16481 7792 16486 7848
rect 16542 7792 16590 7848
rect 16481 7790 16590 7792
rect 16481 7787 16547 7790
rect 17128 7748 17188 7926
rect 17128 7744 17418 7748
rect 0 7714 800 7744
rect 933 7714 999 7717
rect 0 7712 999 7714
rect 0 7656 938 7712
rect 994 7656 999 7712
rect 17128 7688 18000 7744
rect 0 7654 999 7656
rect 0 7624 800 7654
rect 933 7651 999 7654
rect 4878 7648 5194 7649
rect 4878 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5194 7648
rect 4878 7583 5194 7584
rect 8811 7648 9127 7649
rect 8811 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9127 7648
rect 8811 7583 9127 7584
rect 12744 7648 13060 7649
rect 12744 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13060 7648
rect 12744 7583 13060 7584
rect 16677 7648 16993 7649
rect 16677 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16993 7648
rect 17200 7624 18000 7688
rect 16677 7583 16993 7584
rect 2912 7104 3228 7105
rect 2912 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3228 7104
rect 2912 7039 3228 7040
rect 6845 7104 7161 7105
rect 6845 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7161 7104
rect 6845 7039 7161 7040
rect 10778 7104 11094 7105
rect 10778 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11094 7104
rect 10778 7039 11094 7040
rect 14711 7104 15027 7105
rect 14711 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15027 7104
rect 14711 7039 15027 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 5625 6898 5691 6901
rect 14825 6898 14891 6901
rect 5625 6896 14891 6898
rect 5625 6840 5630 6896
rect 5686 6840 14830 6896
rect 14886 6840 14891 6896
rect 5625 6838 14891 6840
rect 5625 6835 5691 6838
rect 14825 6835 14891 6838
rect 16573 6898 16639 6901
rect 17200 6898 18000 6928
rect 16573 6896 18000 6898
rect 16573 6840 16578 6896
rect 16634 6840 18000 6896
rect 16573 6838 18000 6840
rect 16573 6835 16639 6838
rect 17200 6808 18000 6838
rect 4878 6560 5194 6561
rect 4878 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5194 6560
rect 4878 6495 5194 6496
rect 8811 6560 9127 6561
rect 8811 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9127 6560
rect 8811 6495 9127 6496
rect 12744 6560 13060 6561
rect 12744 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13060 6560
rect 12744 6495 13060 6496
rect 16677 6560 16993 6561
rect 16677 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16993 6560
rect 16677 6495 16993 6496
rect 13629 6490 13695 6493
rect 15745 6490 15811 6493
rect 13629 6488 15811 6490
rect 13629 6432 13634 6488
rect 13690 6432 15750 6488
rect 15806 6432 15811 6488
rect 13629 6430 15811 6432
rect 13629 6427 13695 6430
rect 15745 6427 15811 6430
rect 6453 6354 6519 6357
rect 8753 6354 8819 6357
rect 6453 6352 8819 6354
rect 6453 6296 6458 6352
rect 6514 6296 8758 6352
rect 8814 6296 8819 6352
rect 6453 6294 8819 6296
rect 6453 6291 6519 6294
rect 8753 6291 8819 6294
rect 15837 6354 15903 6357
rect 15837 6352 15946 6354
rect 15837 6296 15842 6352
rect 15898 6296 15946 6352
rect 15837 6291 15946 6296
rect 15886 6221 15946 6291
rect 3325 6218 3391 6221
rect 8017 6218 8083 6221
rect 3325 6216 8083 6218
rect 3325 6160 3330 6216
rect 3386 6160 8022 6216
rect 8078 6160 8083 6216
rect 3325 6158 8083 6160
rect 3325 6155 3391 6158
rect 8017 6155 8083 6158
rect 14825 6218 14891 6221
rect 14825 6216 15210 6218
rect 14825 6160 14830 6216
rect 14886 6160 15210 6216
rect 14825 6158 15210 6160
rect 14825 6155 14891 6158
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 15150 6082 15210 6158
rect 15837 6216 15946 6221
rect 15837 6160 15842 6216
rect 15898 6160 15946 6216
rect 15837 6158 15946 6160
rect 15837 6155 15903 6158
rect 17200 6082 18000 6112
rect 15150 6022 18000 6082
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 2912 6016 3228 6017
rect 2912 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3228 6016
rect 2912 5951 3228 5952
rect 6845 6016 7161 6017
rect 6845 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7161 6016
rect 6845 5951 7161 5952
rect 10778 6016 11094 6017
rect 10778 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11094 6016
rect 10778 5951 11094 5952
rect 14711 6016 15027 6017
rect 14711 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15027 6016
rect 17200 5992 18000 6022
rect 14711 5951 15027 5952
rect 7833 5810 7899 5813
rect 8661 5810 8727 5813
rect 7833 5808 8727 5810
rect 7833 5752 7838 5808
rect 7894 5752 8666 5808
rect 8722 5752 8727 5808
rect 7833 5750 8727 5752
rect 7833 5747 7899 5750
rect 8661 5747 8727 5750
rect 7833 5674 7899 5677
rect 8937 5674 9003 5677
rect 7833 5672 9003 5674
rect 7833 5616 7838 5672
rect 7894 5616 8942 5672
rect 8998 5616 9003 5672
rect 7833 5614 9003 5616
rect 7833 5611 7899 5614
rect 8937 5611 9003 5614
rect 1485 5538 1551 5541
rect 11237 5540 11303 5541
rect 11237 5538 11284 5540
rect 798 5536 1551 5538
rect 798 5480 1490 5536
rect 1546 5480 1551 5536
rect 798 5478 1551 5480
rect 11192 5536 11284 5538
rect 11192 5480 11242 5536
rect 11192 5478 11284 5480
rect 798 5296 858 5478
rect 1485 5475 1551 5478
rect 11237 5476 11284 5478
rect 11348 5476 11354 5540
rect 11237 5475 11303 5476
rect 4878 5472 5194 5473
rect 4878 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5194 5472
rect 4878 5407 5194 5408
rect 8811 5472 9127 5473
rect 8811 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9127 5472
rect 8811 5407 9127 5408
rect 12744 5472 13060 5473
rect 12744 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13060 5472
rect 12744 5407 13060 5408
rect 16677 5472 16993 5473
rect 16677 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16993 5472
rect 16677 5407 16993 5408
rect 0 5206 858 5296
rect 7373 5266 7439 5269
rect 8937 5266 9003 5269
rect 7373 5264 9003 5266
rect 7373 5208 7378 5264
rect 7434 5208 8942 5264
rect 8998 5208 9003 5264
rect 7373 5206 9003 5208
rect 0 5176 800 5206
rect 7373 5203 7439 5206
rect 8937 5203 9003 5206
rect 13813 5266 13879 5269
rect 17200 5266 18000 5296
rect 13813 5264 18000 5266
rect 13813 5208 13818 5264
rect 13874 5208 18000 5264
rect 13813 5206 18000 5208
rect 13813 5203 13879 5206
rect 17200 5176 18000 5206
rect 2912 4928 3228 4929
rect 2912 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3228 4928
rect 2912 4863 3228 4864
rect 6845 4928 7161 4929
rect 6845 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7161 4928
rect 6845 4863 7161 4864
rect 10778 4928 11094 4929
rect 10778 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11094 4928
rect 10778 4863 11094 4864
rect 14711 4928 15027 4929
rect 14711 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15027 4928
rect 14711 4863 15027 4864
rect 12433 4586 12499 4589
rect 16990 4586 17188 4620
rect 12433 4584 17188 4586
rect 12433 4528 12438 4584
rect 12494 4560 17188 4584
rect 12494 4528 17050 4560
rect 12433 4526 17050 4528
rect 12433 4523 12499 4526
rect 17128 4484 17188 4560
rect 17128 4480 17418 4484
rect 0 4450 800 4480
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 17128 4424 18000 4480
rect 0 4390 999 4392
rect 0 4360 800 4390
rect 933 4387 999 4390
rect 4878 4384 5194 4385
rect 4878 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5194 4384
rect 4878 4319 5194 4320
rect 8811 4384 9127 4385
rect 8811 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9127 4384
rect 8811 4319 9127 4320
rect 12744 4384 13060 4385
rect 12744 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13060 4384
rect 12744 4319 13060 4320
rect 16677 4384 16993 4385
rect 16677 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16993 4384
rect 17200 4360 18000 4424
rect 16677 4319 16993 4320
rect 13905 4042 13971 4045
rect 16297 4044 16363 4045
rect 14406 4042 14412 4044
rect 13905 4040 14412 4042
rect 13905 3984 13910 4040
rect 13966 3984 14412 4040
rect 13905 3982 14412 3984
rect 13905 3979 13971 3982
rect 14406 3980 14412 3982
rect 14476 3980 14482 4044
rect 16246 3980 16252 4044
rect 16316 4042 16363 4044
rect 16316 4040 16408 4042
rect 16358 3984 16408 4040
rect 16316 3982 16408 3984
rect 16316 3980 16363 3982
rect 16297 3979 16363 3980
rect 2912 3840 3228 3841
rect 2912 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3228 3840
rect 2912 3775 3228 3776
rect 6845 3840 7161 3841
rect 6845 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7161 3840
rect 6845 3775 7161 3776
rect 10778 3840 11094 3841
rect 10778 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11094 3840
rect 10778 3775 11094 3776
rect 14711 3840 15027 3841
rect 14711 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15027 3840
rect 14711 3775 15027 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 14365 3634 14431 3637
rect 17200 3634 18000 3664
rect 14365 3632 18000 3634
rect 14365 3576 14370 3632
rect 14426 3576 18000 3632
rect 14365 3574 18000 3576
rect 14365 3571 14431 3574
rect 17200 3544 18000 3574
rect 4878 3296 5194 3297
rect 4878 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5194 3296
rect 4878 3231 5194 3232
rect 8811 3296 9127 3297
rect 8811 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9127 3296
rect 8811 3231 9127 3232
rect 12744 3296 13060 3297
rect 12744 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13060 3296
rect 12744 3231 13060 3232
rect 16677 3296 16993 3297
rect 16677 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16993 3296
rect 16677 3231 16993 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 15653 2818 15719 2821
rect 17200 2818 18000 2848
rect 15653 2816 18000 2818
rect 15653 2760 15658 2816
rect 15714 2760 18000 2816
rect 15653 2758 18000 2760
rect 15653 2755 15719 2758
rect 2912 2752 3228 2753
rect 2912 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3228 2752
rect 2912 2687 3228 2688
rect 6845 2752 7161 2753
rect 6845 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7161 2752
rect 6845 2687 7161 2688
rect 10778 2752 11094 2753
rect 10778 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11094 2752
rect 10778 2687 11094 2688
rect 14711 2752 15027 2753
rect 14711 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15027 2752
rect 17200 2728 18000 2758
rect 14711 2687 15027 2688
rect 11421 2682 11487 2685
rect 14222 2682 14228 2684
rect 11421 2680 14228 2682
rect 11421 2624 11426 2680
rect 11482 2624 14228 2680
rect 11421 2622 14228 2624
rect 11421 2619 11487 2622
rect 14222 2620 14228 2622
rect 14292 2620 14298 2684
rect 9397 2546 9463 2549
rect 11881 2546 11947 2549
rect 9397 2544 11947 2546
rect 9397 2488 9402 2544
rect 9458 2488 11886 2544
rect 11942 2488 11947 2544
rect 9397 2486 11947 2488
rect 9397 2483 9463 2486
rect 11881 2483 11947 2486
rect 4878 2208 5194 2209
rect 4878 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5194 2208
rect 4878 2143 5194 2144
rect 8811 2208 9127 2209
rect 8811 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9127 2208
rect 8811 2143 9127 2144
rect 12744 2208 13060 2209
rect 12744 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13060 2208
rect 12744 2143 13060 2144
rect 16677 2208 16993 2209
rect 16677 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16993 2208
rect 16677 2143 16993 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
rect 16573 2002 16639 2005
rect 17200 2002 18000 2032
rect 16573 2000 18000 2002
rect 16573 1944 16578 2000
rect 16634 1944 18000 2000
rect 16573 1942 18000 1944
rect 16573 1939 16639 1942
rect 17200 1912 18000 1942
rect 16297 1186 16363 1189
rect 17200 1186 18000 1216
rect 16297 1184 18000 1186
rect 16297 1128 16302 1184
rect 16358 1128 18000 1184
rect 16297 1126 18000 1128
rect 16297 1123 16363 1126
rect 17200 1096 18000 1126
rect 13813 370 13879 373
rect 17200 370 18000 400
rect 13813 368 18000 370
rect 13813 312 13818 368
rect 13874 312 18000 368
rect 13813 310 18000 312
rect 13813 307 13879 310
rect 17200 280 18000 310
<< via3 >>
rect 2918 15804 2982 15808
rect 2918 15748 2922 15804
rect 2922 15748 2978 15804
rect 2978 15748 2982 15804
rect 2918 15744 2982 15748
rect 2998 15804 3062 15808
rect 2998 15748 3002 15804
rect 3002 15748 3058 15804
rect 3058 15748 3062 15804
rect 2998 15744 3062 15748
rect 3078 15804 3142 15808
rect 3078 15748 3082 15804
rect 3082 15748 3138 15804
rect 3138 15748 3142 15804
rect 3078 15744 3142 15748
rect 3158 15804 3222 15808
rect 3158 15748 3162 15804
rect 3162 15748 3218 15804
rect 3218 15748 3222 15804
rect 3158 15744 3222 15748
rect 6851 15804 6915 15808
rect 6851 15748 6855 15804
rect 6855 15748 6911 15804
rect 6911 15748 6915 15804
rect 6851 15744 6915 15748
rect 6931 15804 6995 15808
rect 6931 15748 6935 15804
rect 6935 15748 6991 15804
rect 6991 15748 6995 15804
rect 6931 15744 6995 15748
rect 7011 15804 7075 15808
rect 7011 15748 7015 15804
rect 7015 15748 7071 15804
rect 7071 15748 7075 15804
rect 7011 15744 7075 15748
rect 7091 15804 7155 15808
rect 7091 15748 7095 15804
rect 7095 15748 7151 15804
rect 7151 15748 7155 15804
rect 7091 15744 7155 15748
rect 10784 15804 10848 15808
rect 10784 15748 10788 15804
rect 10788 15748 10844 15804
rect 10844 15748 10848 15804
rect 10784 15744 10848 15748
rect 10864 15804 10928 15808
rect 10864 15748 10868 15804
rect 10868 15748 10924 15804
rect 10924 15748 10928 15804
rect 10864 15744 10928 15748
rect 10944 15804 11008 15808
rect 10944 15748 10948 15804
rect 10948 15748 11004 15804
rect 11004 15748 11008 15804
rect 10944 15744 11008 15748
rect 11024 15804 11088 15808
rect 11024 15748 11028 15804
rect 11028 15748 11084 15804
rect 11084 15748 11088 15804
rect 11024 15744 11088 15748
rect 14717 15804 14781 15808
rect 14717 15748 14721 15804
rect 14721 15748 14777 15804
rect 14777 15748 14781 15804
rect 14717 15744 14781 15748
rect 14797 15804 14861 15808
rect 14797 15748 14801 15804
rect 14801 15748 14857 15804
rect 14857 15748 14861 15804
rect 14797 15744 14861 15748
rect 14877 15804 14941 15808
rect 14877 15748 14881 15804
rect 14881 15748 14937 15804
rect 14937 15748 14941 15804
rect 14877 15744 14941 15748
rect 14957 15804 15021 15808
rect 14957 15748 14961 15804
rect 14961 15748 15017 15804
rect 15017 15748 15021 15804
rect 14957 15744 15021 15748
rect 4884 15260 4948 15264
rect 4884 15204 4888 15260
rect 4888 15204 4944 15260
rect 4944 15204 4948 15260
rect 4884 15200 4948 15204
rect 4964 15260 5028 15264
rect 4964 15204 4968 15260
rect 4968 15204 5024 15260
rect 5024 15204 5028 15260
rect 4964 15200 5028 15204
rect 5044 15260 5108 15264
rect 5044 15204 5048 15260
rect 5048 15204 5104 15260
rect 5104 15204 5108 15260
rect 5044 15200 5108 15204
rect 5124 15260 5188 15264
rect 5124 15204 5128 15260
rect 5128 15204 5184 15260
rect 5184 15204 5188 15260
rect 5124 15200 5188 15204
rect 8817 15260 8881 15264
rect 8817 15204 8821 15260
rect 8821 15204 8877 15260
rect 8877 15204 8881 15260
rect 8817 15200 8881 15204
rect 8897 15260 8961 15264
rect 8897 15204 8901 15260
rect 8901 15204 8957 15260
rect 8957 15204 8961 15260
rect 8897 15200 8961 15204
rect 8977 15260 9041 15264
rect 8977 15204 8981 15260
rect 8981 15204 9037 15260
rect 9037 15204 9041 15260
rect 8977 15200 9041 15204
rect 9057 15260 9121 15264
rect 9057 15204 9061 15260
rect 9061 15204 9117 15260
rect 9117 15204 9121 15260
rect 9057 15200 9121 15204
rect 12750 15260 12814 15264
rect 12750 15204 12754 15260
rect 12754 15204 12810 15260
rect 12810 15204 12814 15260
rect 12750 15200 12814 15204
rect 12830 15260 12894 15264
rect 12830 15204 12834 15260
rect 12834 15204 12890 15260
rect 12890 15204 12894 15260
rect 12830 15200 12894 15204
rect 12910 15260 12974 15264
rect 12910 15204 12914 15260
rect 12914 15204 12970 15260
rect 12970 15204 12974 15260
rect 12910 15200 12974 15204
rect 12990 15260 13054 15264
rect 12990 15204 12994 15260
rect 12994 15204 13050 15260
rect 13050 15204 13054 15260
rect 12990 15200 13054 15204
rect 16683 15260 16747 15264
rect 16683 15204 16687 15260
rect 16687 15204 16743 15260
rect 16743 15204 16747 15260
rect 16683 15200 16747 15204
rect 16763 15260 16827 15264
rect 16763 15204 16767 15260
rect 16767 15204 16823 15260
rect 16823 15204 16827 15260
rect 16763 15200 16827 15204
rect 16843 15260 16907 15264
rect 16843 15204 16847 15260
rect 16847 15204 16903 15260
rect 16903 15204 16907 15260
rect 16843 15200 16907 15204
rect 16923 15260 16987 15264
rect 16923 15204 16927 15260
rect 16927 15204 16983 15260
rect 16983 15204 16987 15260
rect 16923 15200 16987 15204
rect 2918 14716 2982 14720
rect 2918 14660 2922 14716
rect 2922 14660 2978 14716
rect 2978 14660 2982 14716
rect 2918 14656 2982 14660
rect 2998 14716 3062 14720
rect 2998 14660 3002 14716
rect 3002 14660 3058 14716
rect 3058 14660 3062 14716
rect 2998 14656 3062 14660
rect 3078 14716 3142 14720
rect 3078 14660 3082 14716
rect 3082 14660 3138 14716
rect 3138 14660 3142 14716
rect 3078 14656 3142 14660
rect 3158 14716 3222 14720
rect 3158 14660 3162 14716
rect 3162 14660 3218 14716
rect 3218 14660 3222 14716
rect 3158 14656 3222 14660
rect 6851 14716 6915 14720
rect 6851 14660 6855 14716
rect 6855 14660 6911 14716
rect 6911 14660 6915 14716
rect 6851 14656 6915 14660
rect 6931 14716 6995 14720
rect 6931 14660 6935 14716
rect 6935 14660 6991 14716
rect 6991 14660 6995 14716
rect 6931 14656 6995 14660
rect 7011 14716 7075 14720
rect 7011 14660 7015 14716
rect 7015 14660 7071 14716
rect 7071 14660 7075 14716
rect 7011 14656 7075 14660
rect 7091 14716 7155 14720
rect 7091 14660 7095 14716
rect 7095 14660 7151 14716
rect 7151 14660 7155 14716
rect 7091 14656 7155 14660
rect 10784 14716 10848 14720
rect 10784 14660 10788 14716
rect 10788 14660 10844 14716
rect 10844 14660 10848 14716
rect 10784 14656 10848 14660
rect 10864 14716 10928 14720
rect 10864 14660 10868 14716
rect 10868 14660 10924 14716
rect 10924 14660 10928 14716
rect 10864 14656 10928 14660
rect 10944 14716 11008 14720
rect 10944 14660 10948 14716
rect 10948 14660 11004 14716
rect 11004 14660 11008 14716
rect 10944 14656 11008 14660
rect 11024 14716 11088 14720
rect 11024 14660 11028 14716
rect 11028 14660 11084 14716
rect 11084 14660 11088 14716
rect 11024 14656 11088 14660
rect 14717 14716 14781 14720
rect 14717 14660 14721 14716
rect 14721 14660 14777 14716
rect 14777 14660 14781 14716
rect 14717 14656 14781 14660
rect 14797 14716 14861 14720
rect 14797 14660 14801 14716
rect 14801 14660 14857 14716
rect 14857 14660 14861 14716
rect 14797 14656 14861 14660
rect 14877 14716 14941 14720
rect 14877 14660 14881 14716
rect 14881 14660 14937 14716
rect 14937 14660 14941 14716
rect 14877 14656 14941 14660
rect 14957 14716 15021 14720
rect 14957 14660 14961 14716
rect 14961 14660 15017 14716
rect 15017 14660 15021 14716
rect 14957 14656 15021 14660
rect 4884 14172 4948 14176
rect 4884 14116 4888 14172
rect 4888 14116 4944 14172
rect 4944 14116 4948 14172
rect 4884 14112 4948 14116
rect 4964 14172 5028 14176
rect 4964 14116 4968 14172
rect 4968 14116 5024 14172
rect 5024 14116 5028 14172
rect 4964 14112 5028 14116
rect 5044 14172 5108 14176
rect 5044 14116 5048 14172
rect 5048 14116 5104 14172
rect 5104 14116 5108 14172
rect 5044 14112 5108 14116
rect 5124 14172 5188 14176
rect 5124 14116 5128 14172
rect 5128 14116 5184 14172
rect 5184 14116 5188 14172
rect 5124 14112 5188 14116
rect 8817 14172 8881 14176
rect 8817 14116 8821 14172
rect 8821 14116 8877 14172
rect 8877 14116 8881 14172
rect 8817 14112 8881 14116
rect 8897 14172 8961 14176
rect 8897 14116 8901 14172
rect 8901 14116 8957 14172
rect 8957 14116 8961 14172
rect 8897 14112 8961 14116
rect 8977 14172 9041 14176
rect 8977 14116 8981 14172
rect 8981 14116 9037 14172
rect 9037 14116 9041 14172
rect 8977 14112 9041 14116
rect 9057 14172 9121 14176
rect 9057 14116 9061 14172
rect 9061 14116 9117 14172
rect 9117 14116 9121 14172
rect 9057 14112 9121 14116
rect 12750 14172 12814 14176
rect 12750 14116 12754 14172
rect 12754 14116 12810 14172
rect 12810 14116 12814 14172
rect 12750 14112 12814 14116
rect 12830 14172 12894 14176
rect 12830 14116 12834 14172
rect 12834 14116 12890 14172
rect 12890 14116 12894 14172
rect 12830 14112 12894 14116
rect 12910 14172 12974 14176
rect 12910 14116 12914 14172
rect 12914 14116 12970 14172
rect 12970 14116 12974 14172
rect 12910 14112 12974 14116
rect 12990 14172 13054 14176
rect 12990 14116 12994 14172
rect 12994 14116 13050 14172
rect 13050 14116 13054 14172
rect 12990 14112 13054 14116
rect 16683 14172 16747 14176
rect 16683 14116 16687 14172
rect 16687 14116 16743 14172
rect 16743 14116 16747 14172
rect 16683 14112 16747 14116
rect 16763 14172 16827 14176
rect 16763 14116 16767 14172
rect 16767 14116 16823 14172
rect 16823 14116 16827 14172
rect 16763 14112 16827 14116
rect 16843 14172 16907 14176
rect 16843 14116 16847 14172
rect 16847 14116 16903 14172
rect 16903 14116 16907 14172
rect 16843 14112 16907 14116
rect 16923 14172 16987 14176
rect 16923 14116 16927 14172
rect 16927 14116 16983 14172
rect 16983 14116 16987 14172
rect 16923 14112 16987 14116
rect 2918 13628 2982 13632
rect 2918 13572 2922 13628
rect 2922 13572 2978 13628
rect 2978 13572 2982 13628
rect 2918 13568 2982 13572
rect 2998 13628 3062 13632
rect 2998 13572 3002 13628
rect 3002 13572 3058 13628
rect 3058 13572 3062 13628
rect 2998 13568 3062 13572
rect 3078 13628 3142 13632
rect 3078 13572 3082 13628
rect 3082 13572 3138 13628
rect 3138 13572 3142 13628
rect 3078 13568 3142 13572
rect 3158 13628 3222 13632
rect 3158 13572 3162 13628
rect 3162 13572 3218 13628
rect 3218 13572 3222 13628
rect 3158 13568 3222 13572
rect 6851 13628 6915 13632
rect 6851 13572 6855 13628
rect 6855 13572 6911 13628
rect 6911 13572 6915 13628
rect 6851 13568 6915 13572
rect 6931 13628 6995 13632
rect 6931 13572 6935 13628
rect 6935 13572 6991 13628
rect 6991 13572 6995 13628
rect 6931 13568 6995 13572
rect 7011 13628 7075 13632
rect 7011 13572 7015 13628
rect 7015 13572 7071 13628
rect 7071 13572 7075 13628
rect 7011 13568 7075 13572
rect 7091 13628 7155 13632
rect 7091 13572 7095 13628
rect 7095 13572 7151 13628
rect 7151 13572 7155 13628
rect 7091 13568 7155 13572
rect 10784 13628 10848 13632
rect 10784 13572 10788 13628
rect 10788 13572 10844 13628
rect 10844 13572 10848 13628
rect 10784 13568 10848 13572
rect 10864 13628 10928 13632
rect 10864 13572 10868 13628
rect 10868 13572 10924 13628
rect 10924 13572 10928 13628
rect 10864 13568 10928 13572
rect 10944 13628 11008 13632
rect 10944 13572 10948 13628
rect 10948 13572 11004 13628
rect 11004 13572 11008 13628
rect 10944 13568 11008 13572
rect 11024 13628 11088 13632
rect 11024 13572 11028 13628
rect 11028 13572 11084 13628
rect 11084 13572 11088 13628
rect 11024 13568 11088 13572
rect 14717 13628 14781 13632
rect 14717 13572 14721 13628
rect 14721 13572 14777 13628
rect 14777 13572 14781 13628
rect 14717 13568 14781 13572
rect 14797 13628 14861 13632
rect 14797 13572 14801 13628
rect 14801 13572 14857 13628
rect 14857 13572 14861 13628
rect 14797 13568 14861 13572
rect 14877 13628 14941 13632
rect 14877 13572 14881 13628
rect 14881 13572 14937 13628
rect 14937 13572 14941 13628
rect 14877 13568 14941 13572
rect 14957 13628 15021 13632
rect 14957 13572 14961 13628
rect 14961 13572 15017 13628
rect 15017 13572 15021 13628
rect 14957 13568 15021 13572
rect 4884 13084 4948 13088
rect 4884 13028 4888 13084
rect 4888 13028 4944 13084
rect 4944 13028 4948 13084
rect 4884 13024 4948 13028
rect 4964 13084 5028 13088
rect 4964 13028 4968 13084
rect 4968 13028 5024 13084
rect 5024 13028 5028 13084
rect 4964 13024 5028 13028
rect 5044 13084 5108 13088
rect 5044 13028 5048 13084
rect 5048 13028 5104 13084
rect 5104 13028 5108 13084
rect 5044 13024 5108 13028
rect 5124 13084 5188 13088
rect 5124 13028 5128 13084
rect 5128 13028 5184 13084
rect 5184 13028 5188 13084
rect 5124 13024 5188 13028
rect 8817 13084 8881 13088
rect 8817 13028 8821 13084
rect 8821 13028 8877 13084
rect 8877 13028 8881 13084
rect 8817 13024 8881 13028
rect 8897 13084 8961 13088
rect 8897 13028 8901 13084
rect 8901 13028 8957 13084
rect 8957 13028 8961 13084
rect 8897 13024 8961 13028
rect 8977 13084 9041 13088
rect 8977 13028 8981 13084
rect 8981 13028 9037 13084
rect 9037 13028 9041 13084
rect 8977 13024 9041 13028
rect 9057 13084 9121 13088
rect 9057 13028 9061 13084
rect 9061 13028 9117 13084
rect 9117 13028 9121 13084
rect 9057 13024 9121 13028
rect 12750 13084 12814 13088
rect 12750 13028 12754 13084
rect 12754 13028 12810 13084
rect 12810 13028 12814 13084
rect 12750 13024 12814 13028
rect 12830 13084 12894 13088
rect 12830 13028 12834 13084
rect 12834 13028 12890 13084
rect 12890 13028 12894 13084
rect 12830 13024 12894 13028
rect 12910 13084 12974 13088
rect 12910 13028 12914 13084
rect 12914 13028 12970 13084
rect 12970 13028 12974 13084
rect 12910 13024 12974 13028
rect 12990 13084 13054 13088
rect 12990 13028 12994 13084
rect 12994 13028 13050 13084
rect 13050 13028 13054 13084
rect 12990 13024 13054 13028
rect 16683 13084 16747 13088
rect 16683 13028 16687 13084
rect 16687 13028 16743 13084
rect 16743 13028 16747 13084
rect 16683 13024 16747 13028
rect 16763 13084 16827 13088
rect 16763 13028 16767 13084
rect 16767 13028 16823 13084
rect 16823 13028 16827 13084
rect 16763 13024 16827 13028
rect 16843 13084 16907 13088
rect 16843 13028 16847 13084
rect 16847 13028 16903 13084
rect 16903 13028 16907 13084
rect 16843 13024 16907 13028
rect 16923 13084 16987 13088
rect 16923 13028 16927 13084
rect 16927 13028 16983 13084
rect 16983 13028 16987 13084
rect 16923 13024 16987 13028
rect 2918 12540 2982 12544
rect 2918 12484 2922 12540
rect 2922 12484 2978 12540
rect 2978 12484 2982 12540
rect 2918 12480 2982 12484
rect 2998 12540 3062 12544
rect 2998 12484 3002 12540
rect 3002 12484 3058 12540
rect 3058 12484 3062 12540
rect 2998 12480 3062 12484
rect 3078 12540 3142 12544
rect 3078 12484 3082 12540
rect 3082 12484 3138 12540
rect 3138 12484 3142 12540
rect 3078 12480 3142 12484
rect 3158 12540 3222 12544
rect 3158 12484 3162 12540
rect 3162 12484 3218 12540
rect 3218 12484 3222 12540
rect 3158 12480 3222 12484
rect 6851 12540 6915 12544
rect 6851 12484 6855 12540
rect 6855 12484 6911 12540
rect 6911 12484 6915 12540
rect 6851 12480 6915 12484
rect 6931 12540 6995 12544
rect 6931 12484 6935 12540
rect 6935 12484 6991 12540
rect 6991 12484 6995 12540
rect 6931 12480 6995 12484
rect 7011 12540 7075 12544
rect 7011 12484 7015 12540
rect 7015 12484 7071 12540
rect 7071 12484 7075 12540
rect 7011 12480 7075 12484
rect 7091 12540 7155 12544
rect 7091 12484 7095 12540
rect 7095 12484 7151 12540
rect 7151 12484 7155 12540
rect 7091 12480 7155 12484
rect 10784 12540 10848 12544
rect 10784 12484 10788 12540
rect 10788 12484 10844 12540
rect 10844 12484 10848 12540
rect 10784 12480 10848 12484
rect 10864 12540 10928 12544
rect 10864 12484 10868 12540
rect 10868 12484 10924 12540
rect 10924 12484 10928 12540
rect 10864 12480 10928 12484
rect 10944 12540 11008 12544
rect 10944 12484 10948 12540
rect 10948 12484 11004 12540
rect 11004 12484 11008 12540
rect 10944 12480 11008 12484
rect 11024 12540 11088 12544
rect 11024 12484 11028 12540
rect 11028 12484 11084 12540
rect 11084 12484 11088 12540
rect 11024 12480 11088 12484
rect 14717 12540 14781 12544
rect 14717 12484 14721 12540
rect 14721 12484 14777 12540
rect 14777 12484 14781 12540
rect 14717 12480 14781 12484
rect 14797 12540 14861 12544
rect 14797 12484 14801 12540
rect 14801 12484 14857 12540
rect 14857 12484 14861 12540
rect 14797 12480 14861 12484
rect 14877 12540 14941 12544
rect 14877 12484 14881 12540
rect 14881 12484 14937 12540
rect 14937 12484 14941 12540
rect 14877 12480 14941 12484
rect 14957 12540 15021 12544
rect 14957 12484 14961 12540
rect 14961 12484 15017 12540
rect 15017 12484 15021 12540
rect 14957 12480 15021 12484
rect 4884 11996 4948 12000
rect 4884 11940 4888 11996
rect 4888 11940 4944 11996
rect 4944 11940 4948 11996
rect 4884 11936 4948 11940
rect 4964 11996 5028 12000
rect 4964 11940 4968 11996
rect 4968 11940 5024 11996
rect 5024 11940 5028 11996
rect 4964 11936 5028 11940
rect 5044 11996 5108 12000
rect 5044 11940 5048 11996
rect 5048 11940 5104 11996
rect 5104 11940 5108 11996
rect 5044 11936 5108 11940
rect 5124 11996 5188 12000
rect 5124 11940 5128 11996
rect 5128 11940 5184 11996
rect 5184 11940 5188 11996
rect 5124 11936 5188 11940
rect 8817 11996 8881 12000
rect 8817 11940 8821 11996
rect 8821 11940 8877 11996
rect 8877 11940 8881 11996
rect 8817 11936 8881 11940
rect 8897 11996 8961 12000
rect 8897 11940 8901 11996
rect 8901 11940 8957 11996
rect 8957 11940 8961 11996
rect 8897 11936 8961 11940
rect 8977 11996 9041 12000
rect 8977 11940 8981 11996
rect 8981 11940 9037 11996
rect 9037 11940 9041 11996
rect 8977 11936 9041 11940
rect 9057 11996 9121 12000
rect 9057 11940 9061 11996
rect 9061 11940 9117 11996
rect 9117 11940 9121 11996
rect 9057 11936 9121 11940
rect 12750 11996 12814 12000
rect 12750 11940 12754 11996
rect 12754 11940 12810 11996
rect 12810 11940 12814 11996
rect 12750 11936 12814 11940
rect 12830 11996 12894 12000
rect 12830 11940 12834 11996
rect 12834 11940 12890 11996
rect 12890 11940 12894 11996
rect 12830 11936 12894 11940
rect 12910 11996 12974 12000
rect 12910 11940 12914 11996
rect 12914 11940 12970 11996
rect 12970 11940 12974 11996
rect 12910 11936 12974 11940
rect 12990 11996 13054 12000
rect 12990 11940 12994 11996
rect 12994 11940 13050 11996
rect 13050 11940 13054 11996
rect 12990 11936 13054 11940
rect 16683 11996 16747 12000
rect 16683 11940 16687 11996
rect 16687 11940 16743 11996
rect 16743 11940 16747 11996
rect 16683 11936 16747 11940
rect 16763 11996 16827 12000
rect 16763 11940 16767 11996
rect 16767 11940 16823 11996
rect 16823 11940 16827 11996
rect 16763 11936 16827 11940
rect 16843 11996 16907 12000
rect 16843 11940 16847 11996
rect 16847 11940 16903 11996
rect 16903 11940 16907 11996
rect 16843 11936 16907 11940
rect 16923 11996 16987 12000
rect 16923 11940 16927 11996
rect 16927 11940 16983 11996
rect 16983 11940 16987 11996
rect 16923 11936 16987 11940
rect 2918 11452 2982 11456
rect 2918 11396 2922 11452
rect 2922 11396 2978 11452
rect 2978 11396 2982 11452
rect 2918 11392 2982 11396
rect 2998 11452 3062 11456
rect 2998 11396 3002 11452
rect 3002 11396 3058 11452
rect 3058 11396 3062 11452
rect 2998 11392 3062 11396
rect 3078 11452 3142 11456
rect 3078 11396 3082 11452
rect 3082 11396 3138 11452
rect 3138 11396 3142 11452
rect 3078 11392 3142 11396
rect 3158 11452 3222 11456
rect 3158 11396 3162 11452
rect 3162 11396 3218 11452
rect 3218 11396 3222 11452
rect 3158 11392 3222 11396
rect 6851 11452 6915 11456
rect 6851 11396 6855 11452
rect 6855 11396 6911 11452
rect 6911 11396 6915 11452
rect 6851 11392 6915 11396
rect 6931 11452 6995 11456
rect 6931 11396 6935 11452
rect 6935 11396 6991 11452
rect 6991 11396 6995 11452
rect 6931 11392 6995 11396
rect 7011 11452 7075 11456
rect 7011 11396 7015 11452
rect 7015 11396 7071 11452
rect 7071 11396 7075 11452
rect 7011 11392 7075 11396
rect 7091 11452 7155 11456
rect 7091 11396 7095 11452
rect 7095 11396 7151 11452
rect 7151 11396 7155 11452
rect 7091 11392 7155 11396
rect 10784 11452 10848 11456
rect 10784 11396 10788 11452
rect 10788 11396 10844 11452
rect 10844 11396 10848 11452
rect 10784 11392 10848 11396
rect 10864 11452 10928 11456
rect 10864 11396 10868 11452
rect 10868 11396 10924 11452
rect 10924 11396 10928 11452
rect 10864 11392 10928 11396
rect 10944 11452 11008 11456
rect 10944 11396 10948 11452
rect 10948 11396 11004 11452
rect 11004 11396 11008 11452
rect 10944 11392 11008 11396
rect 11024 11452 11088 11456
rect 11024 11396 11028 11452
rect 11028 11396 11084 11452
rect 11084 11396 11088 11452
rect 11024 11392 11088 11396
rect 14717 11452 14781 11456
rect 14717 11396 14721 11452
rect 14721 11396 14777 11452
rect 14777 11396 14781 11452
rect 14717 11392 14781 11396
rect 14797 11452 14861 11456
rect 14797 11396 14801 11452
rect 14801 11396 14857 11452
rect 14857 11396 14861 11452
rect 14797 11392 14861 11396
rect 14877 11452 14941 11456
rect 14877 11396 14881 11452
rect 14881 11396 14937 11452
rect 14937 11396 14941 11452
rect 14877 11392 14941 11396
rect 14957 11452 15021 11456
rect 14957 11396 14961 11452
rect 14961 11396 15017 11452
rect 15017 11396 15021 11452
rect 14957 11392 15021 11396
rect 11284 11052 11348 11116
rect 14228 11112 14292 11116
rect 14228 11056 14242 11112
rect 14242 11056 14292 11112
rect 14228 11052 14292 11056
rect 4884 10908 4948 10912
rect 4884 10852 4888 10908
rect 4888 10852 4944 10908
rect 4944 10852 4948 10908
rect 4884 10848 4948 10852
rect 4964 10908 5028 10912
rect 4964 10852 4968 10908
rect 4968 10852 5024 10908
rect 5024 10852 5028 10908
rect 4964 10848 5028 10852
rect 5044 10908 5108 10912
rect 5044 10852 5048 10908
rect 5048 10852 5104 10908
rect 5104 10852 5108 10908
rect 5044 10848 5108 10852
rect 5124 10908 5188 10912
rect 5124 10852 5128 10908
rect 5128 10852 5184 10908
rect 5184 10852 5188 10908
rect 5124 10848 5188 10852
rect 8817 10908 8881 10912
rect 8817 10852 8821 10908
rect 8821 10852 8877 10908
rect 8877 10852 8881 10908
rect 8817 10848 8881 10852
rect 8897 10908 8961 10912
rect 8897 10852 8901 10908
rect 8901 10852 8957 10908
rect 8957 10852 8961 10908
rect 8897 10848 8961 10852
rect 8977 10908 9041 10912
rect 8977 10852 8981 10908
rect 8981 10852 9037 10908
rect 9037 10852 9041 10908
rect 8977 10848 9041 10852
rect 9057 10908 9121 10912
rect 9057 10852 9061 10908
rect 9061 10852 9117 10908
rect 9117 10852 9121 10908
rect 9057 10848 9121 10852
rect 12750 10908 12814 10912
rect 12750 10852 12754 10908
rect 12754 10852 12810 10908
rect 12810 10852 12814 10908
rect 12750 10848 12814 10852
rect 12830 10908 12894 10912
rect 12830 10852 12834 10908
rect 12834 10852 12890 10908
rect 12890 10852 12894 10908
rect 12830 10848 12894 10852
rect 12910 10908 12974 10912
rect 12910 10852 12914 10908
rect 12914 10852 12970 10908
rect 12970 10852 12974 10908
rect 12910 10848 12974 10852
rect 12990 10908 13054 10912
rect 12990 10852 12994 10908
rect 12994 10852 13050 10908
rect 13050 10852 13054 10908
rect 12990 10848 13054 10852
rect 16683 10908 16747 10912
rect 16683 10852 16687 10908
rect 16687 10852 16743 10908
rect 16743 10852 16747 10908
rect 16683 10848 16747 10852
rect 16763 10908 16827 10912
rect 16763 10852 16767 10908
rect 16767 10852 16823 10908
rect 16823 10852 16827 10908
rect 16763 10848 16827 10852
rect 16843 10908 16907 10912
rect 16843 10852 16847 10908
rect 16847 10852 16903 10908
rect 16903 10852 16907 10908
rect 16843 10848 16907 10852
rect 16923 10908 16987 10912
rect 16923 10852 16927 10908
rect 16927 10852 16983 10908
rect 16983 10852 16987 10908
rect 16923 10848 16987 10852
rect 14412 10508 14476 10572
rect 2918 10364 2982 10368
rect 2918 10308 2922 10364
rect 2922 10308 2978 10364
rect 2978 10308 2982 10364
rect 2918 10304 2982 10308
rect 2998 10364 3062 10368
rect 2998 10308 3002 10364
rect 3002 10308 3058 10364
rect 3058 10308 3062 10364
rect 2998 10304 3062 10308
rect 3078 10364 3142 10368
rect 3078 10308 3082 10364
rect 3082 10308 3138 10364
rect 3138 10308 3142 10364
rect 3078 10304 3142 10308
rect 3158 10364 3222 10368
rect 3158 10308 3162 10364
rect 3162 10308 3218 10364
rect 3218 10308 3222 10364
rect 3158 10304 3222 10308
rect 6851 10364 6915 10368
rect 6851 10308 6855 10364
rect 6855 10308 6911 10364
rect 6911 10308 6915 10364
rect 6851 10304 6915 10308
rect 6931 10364 6995 10368
rect 6931 10308 6935 10364
rect 6935 10308 6991 10364
rect 6991 10308 6995 10364
rect 6931 10304 6995 10308
rect 7011 10364 7075 10368
rect 7011 10308 7015 10364
rect 7015 10308 7071 10364
rect 7071 10308 7075 10364
rect 7011 10304 7075 10308
rect 7091 10364 7155 10368
rect 7091 10308 7095 10364
rect 7095 10308 7151 10364
rect 7151 10308 7155 10364
rect 7091 10304 7155 10308
rect 10784 10364 10848 10368
rect 10784 10308 10788 10364
rect 10788 10308 10844 10364
rect 10844 10308 10848 10364
rect 10784 10304 10848 10308
rect 10864 10364 10928 10368
rect 10864 10308 10868 10364
rect 10868 10308 10924 10364
rect 10924 10308 10928 10364
rect 10864 10304 10928 10308
rect 10944 10364 11008 10368
rect 10944 10308 10948 10364
rect 10948 10308 11004 10364
rect 11004 10308 11008 10364
rect 10944 10304 11008 10308
rect 11024 10364 11088 10368
rect 11024 10308 11028 10364
rect 11028 10308 11084 10364
rect 11084 10308 11088 10364
rect 11024 10304 11088 10308
rect 14717 10364 14781 10368
rect 14717 10308 14721 10364
rect 14721 10308 14777 10364
rect 14777 10308 14781 10364
rect 14717 10304 14781 10308
rect 14797 10364 14861 10368
rect 14797 10308 14801 10364
rect 14801 10308 14857 10364
rect 14857 10308 14861 10364
rect 14797 10304 14861 10308
rect 14877 10364 14941 10368
rect 14877 10308 14881 10364
rect 14881 10308 14937 10364
rect 14937 10308 14941 10364
rect 14877 10304 14941 10308
rect 14957 10364 15021 10368
rect 14957 10308 14961 10364
rect 14961 10308 15017 10364
rect 15017 10308 15021 10364
rect 14957 10304 15021 10308
rect 4884 9820 4948 9824
rect 4884 9764 4888 9820
rect 4888 9764 4944 9820
rect 4944 9764 4948 9820
rect 4884 9760 4948 9764
rect 4964 9820 5028 9824
rect 4964 9764 4968 9820
rect 4968 9764 5024 9820
rect 5024 9764 5028 9820
rect 4964 9760 5028 9764
rect 5044 9820 5108 9824
rect 5044 9764 5048 9820
rect 5048 9764 5104 9820
rect 5104 9764 5108 9820
rect 5044 9760 5108 9764
rect 5124 9820 5188 9824
rect 5124 9764 5128 9820
rect 5128 9764 5184 9820
rect 5184 9764 5188 9820
rect 5124 9760 5188 9764
rect 8817 9820 8881 9824
rect 8817 9764 8821 9820
rect 8821 9764 8877 9820
rect 8877 9764 8881 9820
rect 8817 9760 8881 9764
rect 8897 9820 8961 9824
rect 8897 9764 8901 9820
rect 8901 9764 8957 9820
rect 8957 9764 8961 9820
rect 8897 9760 8961 9764
rect 8977 9820 9041 9824
rect 8977 9764 8981 9820
rect 8981 9764 9037 9820
rect 9037 9764 9041 9820
rect 8977 9760 9041 9764
rect 9057 9820 9121 9824
rect 9057 9764 9061 9820
rect 9061 9764 9117 9820
rect 9117 9764 9121 9820
rect 9057 9760 9121 9764
rect 12750 9820 12814 9824
rect 12750 9764 12754 9820
rect 12754 9764 12810 9820
rect 12810 9764 12814 9820
rect 12750 9760 12814 9764
rect 12830 9820 12894 9824
rect 12830 9764 12834 9820
rect 12834 9764 12890 9820
rect 12890 9764 12894 9820
rect 12830 9760 12894 9764
rect 12910 9820 12974 9824
rect 12910 9764 12914 9820
rect 12914 9764 12970 9820
rect 12970 9764 12974 9820
rect 12910 9760 12974 9764
rect 12990 9820 13054 9824
rect 12990 9764 12994 9820
rect 12994 9764 13050 9820
rect 13050 9764 13054 9820
rect 12990 9760 13054 9764
rect 16683 9820 16747 9824
rect 16683 9764 16687 9820
rect 16687 9764 16743 9820
rect 16743 9764 16747 9820
rect 16683 9760 16747 9764
rect 16763 9820 16827 9824
rect 16763 9764 16767 9820
rect 16767 9764 16823 9820
rect 16823 9764 16827 9820
rect 16763 9760 16827 9764
rect 16843 9820 16907 9824
rect 16843 9764 16847 9820
rect 16847 9764 16903 9820
rect 16903 9764 16907 9820
rect 16843 9760 16907 9764
rect 16923 9820 16987 9824
rect 16923 9764 16927 9820
rect 16927 9764 16983 9820
rect 16983 9764 16987 9820
rect 16923 9760 16987 9764
rect 16252 9752 16316 9756
rect 16252 9696 16266 9752
rect 16266 9696 16316 9752
rect 16252 9692 16316 9696
rect 2918 9276 2982 9280
rect 2918 9220 2922 9276
rect 2922 9220 2978 9276
rect 2978 9220 2982 9276
rect 2918 9216 2982 9220
rect 2998 9276 3062 9280
rect 2998 9220 3002 9276
rect 3002 9220 3058 9276
rect 3058 9220 3062 9276
rect 2998 9216 3062 9220
rect 3078 9276 3142 9280
rect 3078 9220 3082 9276
rect 3082 9220 3138 9276
rect 3138 9220 3142 9276
rect 3078 9216 3142 9220
rect 3158 9276 3222 9280
rect 3158 9220 3162 9276
rect 3162 9220 3218 9276
rect 3218 9220 3222 9276
rect 3158 9216 3222 9220
rect 6851 9276 6915 9280
rect 6851 9220 6855 9276
rect 6855 9220 6911 9276
rect 6911 9220 6915 9276
rect 6851 9216 6915 9220
rect 6931 9276 6995 9280
rect 6931 9220 6935 9276
rect 6935 9220 6991 9276
rect 6991 9220 6995 9276
rect 6931 9216 6995 9220
rect 7011 9276 7075 9280
rect 7011 9220 7015 9276
rect 7015 9220 7071 9276
rect 7071 9220 7075 9276
rect 7011 9216 7075 9220
rect 7091 9276 7155 9280
rect 7091 9220 7095 9276
rect 7095 9220 7151 9276
rect 7151 9220 7155 9276
rect 7091 9216 7155 9220
rect 10784 9276 10848 9280
rect 10784 9220 10788 9276
rect 10788 9220 10844 9276
rect 10844 9220 10848 9276
rect 10784 9216 10848 9220
rect 10864 9276 10928 9280
rect 10864 9220 10868 9276
rect 10868 9220 10924 9276
rect 10924 9220 10928 9276
rect 10864 9216 10928 9220
rect 10944 9276 11008 9280
rect 10944 9220 10948 9276
rect 10948 9220 11004 9276
rect 11004 9220 11008 9276
rect 10944 9216 11008 9220
rect 11024 9276 11088 9280
rect 11024 9220 11028 9276
rect 11028 9220 11084 9276
rect 11084 9220 11088 9276
rect 11024 9216 11088 9220
rect 14717 9276 14781 9280
rect 14717 9220 14721 9276
rect 14721 9220 14777 9276
rect 14777 9220 14781 9276
rect 14717 9216 14781 9220
rect 14797 9276 14861 9280
rect 14797 9220 14801 9276
rect 14801 9220 14857 9276
rect 14857 9220 14861 9276
rect 14797 9216 14861 9220
rect 14877 9276 14941 9280
rect 14877 9220 14881 9276
rect 14881 9220 14937 9276
rect 14937 9220 14941 9276
rect 14877 9216 14941 9220
rect 14957 9276 15021 9280
rect 14957 9220 14961 9276
rect 14961 9220 15017 9276
rect 15017 9220 15021 9276
rect 14957 9216 15021 9220
rect 4884 8732 4948 8736
rect 4884 8676 4888 8732
rect 4888 8676 4944 8732
rect 4944 8676 4948 8732
rect 4884 8672 4948 8676
rect 4964 8732 5028 8736
rect 4964 8676 4968 8732
rect 4968 8676 5024 8732
rect 5024 8676 5028 8732
rect 4964 8672 5028 8676
rect 5044 8732 5108 8736
rect 5044 8676 5048 8732
rect 5048 8676 5104 8732
rect 5104 8676 5108 8732
rect 5044 8672 5108 8676
rect 5124 8732 5188 8736
rect 5124 8676 5128 8732
rect 5128 8676 5184 8732
rect 5184 8676 5188 8732
rect 5124 8672 5188 8676
rect 8817 8732 8881 8736
rect 8817 8676 8821 8732
rect 8821 8676 8877 8732
rect 8877 8676 8881 8732
rect 8817 8672 8881 8676
rect 8897 8732 8961 8736
rect 8897 8676 8901 8732
rect 8901 8676 8957 8732
rect 8957 8676 8961 8732
rect 8897 8672 8961 8676
rect 8977 8732 9041 8736
rect 8977 8676 8981 8732
rect 8981 8676 9037 8732
rect 9037 8676 9041 8732
rect 8977 8672 9041 8676
rect 9057 8732 9121 8736
rect 9057 8676 9061 8732
rect 9061 8676 9117 8732
rect 9117 8676 9121 8732
rect 9057 8672 9121 8676
rect 12750 8732 12814 8736
rect 12750 8676 12754 8732
rect 12754 8676 12810 8732
rect 12810 8676 12814 8732
rect 12750 8672 12814 8676
rect 12830 8732 12894 8736
rect 12830 8676 12834 8732
rect 12834 8676 12890 8732
rect 12890 8676 12894 8732
rect 12830 8672 12894 8676
rect 12910 8732 12974 8736
rect 12910 8676 12914 8732
rect 12914 8676 12970 8732
rect 12970 8676 12974 8732
rect 12910 8672 12974 8676
rect 12990 8732 13054 8736
rect 12990 8676 12994 8732
rect 12994 8676 13050 8732
rect 13050 8676 13054 8732
rect 12990 8672 13054 8676
rect 16683 8732 16747 8736
rect 16683 8676 16687 8732
rect 16687 8676 16743 8732
rect 16743 8676 16747 8732
rect 16683 8672 16747 8676
rect 16763 8732 16827 8736
rect 16763 8676 16767 8732
rect 16767 8676 16823 8732
rect 16823 8676 16827 8732
rect 16763 8672 16827 8676
rect 16843 8732 16907 8736
rect 16843 8676 16847 8732
rect 16847 8676 16903 8732
rect 16903 8676 16907 8732
rect 16843 8672 16907 8676
rect 16923 8732 16987 8736
rect 16923 8676 16927 8732
rect 16927 8676 16983 8732
rect 16983 8676 16987 8732
rect 16923 8672 16987 8676
rect 2918 8188 2982 8192
rect 2918 8132 2922 8188
rect 2922 8132 2978 8188
rect 2978 8132 2982 8188
rect 2918 8128 2982 8132
rect 2998 8188 3062 8192
rect 2998 8132 3002 8188
rect 3002 8132 3058 8188
rect 3058 8132 3062 8188
rect 2998 8128 3062 8132
rect 3078 8188 3142 8192
rect 3078 8132 3082 8188
rect 3082 8132 3138 8188
rect 3138 8132 3142 8188
rect 3078 8128 3142 8132
rect 3158 8188 3222 8192
rect 3158 8132 3162 8188
rect 3162 8132 3218 8188
rect 3218 8132 3222 8188
rect 3158 8128 3222 8132
rect 6851 8188 6915 8192
rect 6851 8132 6855 8188
rect 6855 8132 6911 8188
rect 6911 8132 6915 8188
rect 6851 8128 6915 8132
rect 6931 8188 6995 8192
rect 6931 8132 6935 8188
rect 6935 8132 6991 8188
rect 6991 8132 6995 8188
rect 6931 8128 6995 8132
rect 7011 8188 7075 8192
rect 7011 8132 7015 8188
rect 7015 8132 7071 8188
rect 7071 8132 7075 8188
rect 7011 8128 7075 8132
rect 7091 8188 7155 8192
rect 7091 8132 7095 8188
rect 7095 8132 7151 8188
rect 7151 8132 7155 8188
rect 7091 8128 7155 8132
rect 10784 8188 10848 8192
rect 10784 8132 10788 8188
rect 10788 8132 10844 8188
rect 10844 8132 10848 8188
rect 10784 8128 10848 8132
rect 10864 8188 10928 8192
rect 10864 8132 10868 8188
rect 10868 8132 10924 8188
rect 10924 8132 10928 8188
rect 10864 8128 10928 8132
rect 10944 8188 11008 8192
rect 10944 8132 10948 8188
rect 10948 8132 11004 8188
rect 11004 8132 11008 8188
rect 10944 8128 11008 8132
rect 11024 8188 11088 8192
rect 11024 8132 11028 8188
rect 11028 8132 11084 8188
rect 11084 8132 11088 8188
rect 11024 8128 11088 8132
rect 14717 8188 14781 8192
rect 14717 8132 14721 8188
rect 14721 8132 14777 8188
rect 14777 8132 14781 8188
rect 14717 8128 14781 8132
rect 14797 8188 14861 8192
rect 14797 8132 14801 8188
rect 14801 8132 14857 8188
rect 14857 8132 14861 8188
rect 14797 8128 14861 8132
rect 14877 8188 14941 8192
rect 14877 8132 14881 8188
rect 14881 8132 14937 8188
rect 14937 8132 14941 8188
rect 14877 8128 14941 8132
rect 14957 8188 15021 8192
rect 14957 8132 14961 8188
rect 14961 8132 15017 8188
rect 15017 8132 15021 8188
rect 14957 8128 15021 8132
rect 4884 7644 4948 7648
rect 4884 7588 4888 7644
rect 4888 7588 4944 7644
rect 4944 7588 4948 7644
rect 4884 7584 4948 7588
rect 4964 7644 5028 7648
rect 4964 7588 4968 7644
rect 4968 7588 5024 7644
rect 5024 7588 5028 7644
rect 4964 7584 5028 7588
rect 5044 7644 5108 7648
rect 5044 7588 5048 7644
rect 5048 7588 5104 7644
rect 5104 7588 5108 7644
rect 5044 7584 5108 7588
rect 5124 7644 5188 7648
rect 5124 7588 5128 7644
rect 5128 7588 5184 7644
rect 5184 7588 5188 7644
rect 5124 7584 5188 7588
rect 8817 7644 8881 7648
rect 8817 7588 8821 7644
rect 8821 7588 8877 7644
rect 8877 7588 8881 7644
rect 8817 7584 8881 7588
rect 8897 7644 8961 7648
rect 8897 7588 8901 7644
rect 8901 7588 8957 7644
rect 8957 7588 8961 7644
rect 8897 7584 8961 7588
rect 8977 7644 9041 7648
rect 8977 7588 8981 7644
rect 8981 7588 9037 7644
rect 9037 7588 9041 7644
rect 8977 7584 9041 7588
rect 9057 7644 9121 7648
rect 9057 7588 9061 7644
rect 9061 7588 9117 7644
rect 9117 7588 9121 7644
rect 9057 7584 9121 7588
rect 12750 7644 12814 7648
rect 12750 7588 12754 7644
rect 12754 7588 12810 7644
rect 12810 7588 12814 7644
rect 12750 7584 12814 7588
rect 12830 7644 12894 7648
rect 12830 7588 12834 7644
rect 12834 7588 12890 7644
rect 12890 7588 12894 7644
rect 12830 7584 12894 7588
rect 12910 7644 12974 7648
rect 12910 7588 12914 7644
rect 12914 7588 12970 7644
rect 12970 7588 12974 7644
rect 12910 7584 12974 7588
rect 12990 7644 13054 7648
rect 12990 7588 12994 7644
rect 12994 7588 13050 7644
rect 13050 7588 13054 7644
rect 12990 7584 13054 7588
rect 16683 7644 16747 7648
rect 16683 7588 16687 7644
rect 16687 7588 16743 7644
rect 16743 7588 16747 7644
rect 16683 7584 16747 7588
rect 16763 7644 16827 7648
rect 16763 7588 16767 7644
rect 16767 7588 16823 7644
rect 16823 7588 16827 7644
rect 16763 7584 16827 7588
rect 16843 7644 16907 7648
rect 16843 7588 16847 7644
rect 16847 7588 16903 7644
rect 16903 7588 16907 7644
rect 16843 7584 16907 7588
rect 16923 7644 16987 7648
rect 16923 7588 16927 7644
rect 16927 7588 16983 7644
rect 16983 7588 16987 7644
rect 16923 7584 16987 7588
rect 2918 7100 2982 7104
rect 2918 7044 2922 7100
rect 2922 7044 2978 7100
rect 2978 7044 2982 7100
rect 2918 7040 2982 7044
rect 2998 7100 3062 7104
rect 2998 7044 3002 7100
rect 3002 7044 3058 7100
rect 3058 7044 3062 7100
rect 2998 7040 3062 7044
rect 3078 7100 3142 7104
rect 3078 7044 3082 7100
rect 3082 7044 3138 7100
rect 3138 7044 3142 7100
rect 3078 7040 3142 7044
rect 3158 7100 3222 7104
rect 3158 7044 3162 7100
rect 3162 7044 3218 7100
rect 3218 7044 3222 7100
rect 3158 7040 3222 7044
rect 6851 7100 6915 7104
rect 6851 7044 6855 7100
rect 6855 7044 6911 7100
rect 6911 7044 6915 7100
rect 6851 7040 6915 7044
rect 6931 7100 6995 7104
rect 6931 7044 6935 7100
rect 6935 7044 6991 7100
rect 6991 7044 6995 7100
rect 6931 7040 6995 7044
rect 7011 7100 7075 7104
rect 7011 7044 7015 7100
rect 7015 7044 7071 7100
rect 7071 7044 7075 7100
rect 7011 7040 7075 7044
rect 7091 7100 7155 7104
rect 7091 7044 7095 7100
rect 7095 7044 7151 7100
rect 7151 7044 7155 7100
rect 7091 7040 7155 7044
rect 10784 7100 10848 7104
rect 10784 7044 10788 7100
rect 10788 7044 10844 7100
rect 10844 7044 10848 7100
rect 10784 7040 10848 7044
rect 10864 7100 10928 7104
rect 10864 7044 10868 7100
rect 10868 7044 10924 7100
rect 10924 7044 10928 7100
rect 10864 7040 10928 7044
rect 10944 7100 11008 7104
rect 10944 7044 10948 7100
rect 10948 7044 11004 7100
rect 11004 7044 11008 7100
rect 10944 7040 11008 7044
rect 11024 7100 11088 7104
rect 11024 7044 11028 7100
rect 11028 7044 11084 7100
rect 11084 7044 11088 7100
rect 11024 7040 11088 7044
rect 14717 7100 14781 7104
rect 14717 7044 14721 7100
rect 14721 7044 14777 7100
rect 14777 7044 14781 7100
rect 14717 7040 14781 7044
rect 14797 7100 14861 7104
rect 14797 7044 14801 7100
rect 14801 7044 14857 7100
rect 14857 7044 14861 7100
rect 14797 7040 14861 7044
rect 14877 7100 14941 7104
rect 14877 7044 14881 7100
rect 14881 7044 14937 7100
rect 14937 7044 14941 7100
rect 14877 7040 14941 7044
rect 14957 7100 15021 7104
rect 14957 7044 14961 7100
rect 14961 7044 15017 7100
rect 15017 7044 15021 7100
rect 14957 7040 15021 7044
rect 4884 6556 4948 6560
rect 4884 6500 4888 6556
rect 4888 6500 4944 6556
rect 4944 6500 4948 6556
rect 4884 6496 4948 6500
rect 4964 6556 5028 6560
rect 4964 6500 4968 6556
rect 4968 6500 5024 6556
rect 5024 6500 5028 6556
rect 4964 6496 5028 6500
rect 5044 6556 5108 6560
rect 5044 6500 5048 6556
rect 5048 6500 5104 6556
rect 5104 6500 5108 6556
rect 5044 6496 5108 6500
rect 5124 6556 5188 6560
rect 5124 6500 5128 6556
rect 5128 6500 5184 6556
rect 5184 6500 5188 6556
rect 5124 6496 5188 6500
rect 8817 6556 8881 6560
rect 8817 6500 8821 6556
rect 8821 6500 8877 6556
rect 8877 6500 8881 6556
rect 8817 6496 8881 6500
rect 8897 6556 8961 6560
rect 8897 6500 8901 6556
rect 8901 6500 8957 6556
rect 8957 6500 8961 6556
rect 8897 6496 8961 6500
rect 8977 6556 9041 6560
rect 8977 6500 8981 6556
rect 8981 6500 9037 6556
rect 9037 6500 9041 6556
rect 8977 6496 9041 6500
rect 9057 6556 9121 6560
rect 9057 6500 9061 6556
rect 9061 6500 9117 6556
rect 9117 6500 9121 6556
rect 9057 6496 9121 6500
rect 12750 6556 12814 6560
rect 12750 6500 12754 6556
rect 12754 6500 12810 6556
rect 12810 6500 12814 6556
rect 12750 6496 12814 6500
rect 12830 6556 12894 6560
rect 12830 6500 12834 6556
rect 12834 6500 12890 6556
rect 12890 6500 12894 6556
rect 12830 6496 12894 6500
rect 12910 6556 12974 6560
rect 12910 6500 12914 6556
rect 12914 6500 12970 6556
rect 12970 6500 12974 6556
rect 12910 6496 12974 6500
rect 12990 6556 13054 6560
rect 12990 6500 12994 6556
rect 12994 6500 13050 6556
rect 13050 6500 13054 6556
rect 12990 6496 13054 6500
rect 16683 6556 16747 6560
rect 16683 6500 16687 6556
rect 16687 6500 16743 6556
rect 16743 6500 16747 6556
rect 16683 6496 16747 6500
rect 16763 6556 16827 6560
rect 16763 6500 16767 6556
rect 16767 6500 16823 6556
rect 16823 6500 16827 6556
rect 16763 6496 16827 6500
rect 16843 6556 16907 6560
rect 16843 6500 16847 6556
rect 16847 6500 16903 6556
rect 16903 6500 16907 6556
rect 16843 6496 16907 6500
rect 16923 6556 16987 6560
rect 16923 6500 16927 6556
rect 16927 6500 16983 6556
rect 16983 6500 16987 6556
rect 16923 6496 16987 6500
rect 2918 6012 2982 6016
rect 2918 5956 2922 6012
rect 2922 5956 2978 6012
rect 2978 5956 2982 6012
rect 2918 5952 2982 5956
rect 2998 6012 3062 6016
rect 2998 5956 3002 6012
rect 3002 5956 3058 6012
rect 3058 5956 3062 6012
rect 2998 5952 3062 5956
rect 3078 6012 3142 6016
rect 3078 5956 3082 6012
rect 3082 5956 3138 6012
rect 3138 5956 3142 6012
rect 3078 5952 3142 5956
rect 3158 6012 3222 6016
rect 3158 5956 3162 6012
rect 3162 5956 3218 6012
rect 3218 5956 3222 6012
rect 3158 5952 3222 5956
rect 6851 6012 6915 6016
rect 6851 5956 6855 6012
rect 6855 5956 6911 6012
rect 6911 5956 6915 6012
rect 6851 5952 6915 5956
rect 6931 6012 6995 6016
rect 6931 5956 6935 6012
rect 6935 5956 6991 6012
rect 6991 5956 6995 6012
rect 6931 5952 6995 5956
rect 7011 6012 7075 6016
rect 7011 5956 7015 6012
rect 7015 5956 7071 6012
rect 7071 5956 7075 6012
rect 7011 5952 7075 5956
rect 7091 6012 7155 6016
rect 7091 5956 7095 6012
rect 7095 5956 7151 6012
rect 7151 5956 7155 6012
rect 7091 5952 7155 5956
rect 10784 6012 10848 6016
rect 10784 5956 10788 6012
rect 10788 5956 10844 6012
rect 10844 5956 10848 6012
rect 10784 5952 10848 5956
rect 10864 6012 10928 6016
rect 10864 5956 10868 6012
rect 10868 5956 10924 6012
rect 10924 5956 10928 6012
rect 10864 5952 10928 5956
rect 10944 6012 11008 6016
rect 10944 5956 10948 6012
rect 10948 5956 11004 6012
rect 11004 5956 11008 6012
rect 10944 5952 11008 5956
rect 11024 6012 11088 6016
rect 11024 5956 11028 6012
rect 11028 5956 11084 6012
rect 11084 5956 11088 6012
rect 11024 5952 11088 5956
rect 14717 6012 14781 6016
rect 14717 5956 14721 6012
rect 14721 5956 14777 6012
rect 14777 5956 14781 6012
rect 14717 5952 14781 5956
rect 14797 6012 14861 6016
rect 14797 5956 14801 6012
rect 14801 5956 14857 6012
rect 14857 5956 14861 6012
rect 14797 5952 14861 5956
rect 14877 6012 14941 6016
rect 14877 5956 14881 6012
rect 14881 5956 14937 6012
rect 14937 5956 14941 6012
rect 14877 5952 14941 5956
rect 14957 6012 15021 6016
rect 14957 5956 14961 6012
rect 14961 5956 15017 6012
rect 15017 5956 15021 6012
rect 14957 5952 15021 5956
rect 11284 5536 11348 5540
rect 11284 5480 11298 5536
rect 11298 5480 11348 5536
rect 11284 5476 11348 5480
rect 4884 5468 4948 5472
rect 4884 5412 4888 5468
rect 4888 5412 4944 5468
rect 4944 5412 4948 5468
rect 4884 5408 4948 5412
rect 4964 5468 5028 5472
rect 4964 5412 4968 5468
rect 4968 5412 5024 5468
rect 5024 5412 5028 5468
rect 4964 5408 5028 5412
rect 5044 5468 5108 5472
rect 5044 5412 5048 5468
rect 5048 5412 5104 5468
rect 5104 5412 5108 5468
rect 5044 5408 5108 5412
rect 5124 5468 5188 5472
rect 5124 5412 5128 5468
rect 5128 5412 5184 5468
rect 5184 5412 5188 5468
rect 5124 5408 5188 5412
rect 8817 5468 8881 5472
rect 8817 5412 8821 5468
rect 8821 5412 8877 5468
rect 8877 5412 8881 5468
rect 8817 5408 8881 5412
rect 8897 5468 8961 5472
rect 8897 5412 8901 5468
rect 8901 5412 8957 5468
rect 8957 5412 8961 5468
rect 8897 5408 8961 5412
rect 8977 5468 9041 5472
rect 8977 5412 8981 5468
rect 8981 5412 9037 5468
rect 9037 5412 9041 5468
rect 8977 5408 9041 5412
rect 9057 5468 9121 5472
rect 9057 5412 9061 5468
rect 9061 5412 9117 5468
rect 9117 5412 9121 5468
rect 9057 5408 9121 5412
rect 12750 5468 12814 5472
rect 12750 5412 12754 5468
rect 12754 5412 12810 5468
rect 12810 5412 12814 5468
rect 12750 5408 12814 5412
rect 12830 5468 12894 5472
rect 12830 5412 12834 5468
rect 12834 5412 12890 5468
rect 12890 5412 12894 5468
rect 12830 5408 12894 5412
rect 12910 5468 12974 5472
rect 12910 5412 12914 5468
rect 12914 5412 12970 5468
rect 12970 5412 12974 5468
rect 12910 5408 12974 5412
rect 12990 5468 13054 5472
rect 12990 5412 12994 5468
rect 12994 5412 13050 5468
rect 13050 5412 13054 5468
rect 12990 5408 13054 5412
rect 16683 5468 16747 5472
rect 16683 5412 16687 5468
rect 16687 5412 16743 5468
rect 16743 5412 16747 5468
rect 16683 5408 16747 5412
rect 16763 5468 16827 5472
rect 16763 5412 16767 5468
rect 16767 5412 16823 5468
rect 16823 5412 16827 5468
rect 16763 5408 16827 5412
rect 16843 5468 16907 5472
rect 16843 5412 16847 5468
rect 16847 5412 16903 5468
rect 16903 5412 16907 5468
rect 16843 5408 16907 5412
rect 16923 5468 16987 5472
rect 16923 5412 16927 5468
rect 16927 5412 16983 5468
rect 16983 5412 16987 5468
rect 16923 5408 16987 5412
rect 2918 4924 2982 4928
rect 2918 4868 2922 4924
rect 2922 4868 2978 4924
rect 2978 4868 2982 4924
rect 2918 4864 2982 4868
rect 2998 4924 3062 4928
rect 2998 4868 3002 4924
rect 3002 4868 3058 4924
rect 3058 4868 3062 4924
rect 2998 4864 3062 4868
rect 3078 4924 3142 4928
rect 3078 4868 3082 4924
rect 3082 4868 3138 4924
rect 3138 4868 3142 4924
rect 3078 4864 3142 4868
rect 3158 4924 3222 4928
rect 3158 4868 3162 4924
rect 3162 4868 3218 4924
rect 3218 4868 3222 4924
rect 3158 4864 3222 4868
rect 6851 4924 6915 4928
rect 6851 4868 6855 4924
rect 6855 4868 6911 4924
rect 6911 4868 6915 4924
rect 6851 4864 6915 4868
rect 6931 4924 6995 4928
rect 6931 4868 6935 4924
rect 6935 4868 6991 4924
rect 6991 4868 6995 4924
rect 6931 4864 6995 4868
rect 7011 4924 7075 4928
rect 7011 4868 7015 4924
rect 7015 4868 7071 4924
rect 7071 4868 7075 4924
rect 7011 4864 7075 4868
rect 7091 4924 7155 4928
rect 7091 4868 7095 4924
rect 7095 4868 7151 4924
rect 7151 4868 7155 4924
rect 7091 4864 7155 4868
rect 10784 4924 10848 4928
rect 10784 4868 10788 4924
rect 10788 4868 10844 4924
rect 10844 4868 10848 4924
rect 10784 4864 10848 4868
rect 10864 4924 10928 4928
rect 10864 4868 10868 4924
rect 10868 4868 10924 4924
rect 10924 4868 10928 4924
rect 10864 4864 10928 4868
rect 10944 4924 11008 4928
rect 10944 4868 10948 4924
rect 10948 4868 11004 4924
rect 11004 4868 11008 4924
rect 10944 4864 11008 4868
rect 11024 4924 11088 4928
rect 11024 4868 11028 4924
rect 11028 4868 11084 4924
rect 11084 4868 11088 4924
rect 11024 4864 11088 4868
rect 14717 4924 14781 4928
rect 14717 4868 14721 4924
rect 14721 4868 14777 4924
rect 14777 4868 14781 4924
rect 14717 4864 14781 4868
rect 14797 4924 14861 4928
rect 14797 4868 14801 4924
rect 14801 4868 14857 4924
rect 14857 4868 14861 4924
rect 14797 4864 14861 4868
rect 14877 4924 14941 4928
rect 14877 4868 14881 4924
rect 14881 4868 14937 4924
rect 14937 4868 14941 4924
rect 14877 4864 14941 4868
rect 14957 4924 15021 4928
rect 14957 4868 14961 4924
rect 14961 4868 15017 4924
rect 15017 4868 15021 4924
rect 14957 4864 15021 4868
rect 4884 4380 4948 4384
rect 4884 4324 4888 4380
rect 4888 4324 4944 4380
rect 4944 4324 4948 4380
rect 4884 4320 4948 4324
rect 4964 4380 5028 4384
rect 4964 4324 4968 4380
rect 4968 4324 5024 4380
rect 5024 4324 5028 4380
rect 4964 4320 5028 4324
rect 5044 4380 5108 4384
rect 5044 4324 5048 4380
rect 5048 4324 5104 4380
rect 5104 4324 5108 4380
rect 5044 4320 5108 4324
rect 5124 4380 5188 4384
rect 5124 4324 5128 4380
rect 5128 4324 5184 4380
rect 5184 4324 5188 4380
rect 5124 4320 5188 4324
rect 8817 4380 8881 4384
rect 8817 4324 8821 4380
rect 8821 4324 8877 4380
rect 8877 4324 8881 4380
rect 8817 4320 8881 4324
rect 8897 4380 8961 4384
rect 8897 4324 8901 4380
rect 8901 4324 8957 4380
rect 8957 4324 8961 4380
rect 8897 4320 8961 4324
rect 8977 4380 9041 4384
rect 8977 4324 8981 4380
rect 8981 4324 9037 4380
rect 9037 4324 9041 4380
rect 8977 4320 9041 4324
rect 9057 4380 9121 4384
rect 9057 4324 9061 4380
rect 9061 4324 9117 4380
rect 9117 4324 9121 4380
rect 9057 4320 9121 4324
rect 12750 4380 12814 4384
rect 12750 4324 12754 4380
rect 12754 4324 12810 4380
rect 12810 4324 12814 4380
rect 12750 4320 12814 4324
rect 12830 4380 12894 4384
rect 12830 4324 12834 4380
rect 12834 4324 12890 4380
rect 12890 4324 12894 4380
rect 12830 4320 12894 4324
rect 12910 4380 12974 4384
rect 12910 4324 12914 4380
rect 12914 4324 12970 4380
rect 12970 4324 12974 4380
rect 12910 4320 12974 4324
rect 12990 4380 13054 4384
rect 12990 4324 12994 4380
rect 12994 4324 13050 4380
rect 13050 4324 13054 4380
rect 12990 4320 13054 4324
rect 16683 4380 16747 4384
rect 16683 4324 16687 4380
rect 16687 4324 16743 4380
rect 16743 4324 16747 4380
rect 16683 4320 16747 4324
rect 16763 4380 16827 4384
rect 16763 4324 16767 4380
rect 16767 4324 16823 4380
rect 16823 4324 16827 4380
rect 16763 4320 16827 4324
rect 16843 4380 16907 4384
rect 16843 4324 16847 4380
rect 16847 4324 16903 4380
rect 16903 4324 16907 4380
rect 16843 4320 16907 4324
rect 16923 4380 16987 4384
rect 16923 4324 16927 4380
rect 16927 4324 16983 4380
rect 16983 4324 16987 4380
rect 16923 4320 16987 4324
rect 14412 3980 14476 4044
rect 16252 4040 16316 4044
rect 16252 3984 16302 4040
rect 16302 3984 16316 4040
rect 16252 3980 16316 3984
rect 2918 3836 2982 3840
rect 2918 3780 2922 3836
rect 2922 3780 2978 3836
rect 2978 3780 2982 3836
rect 2918 3776 2982 3780
rect 2998 3836 3062 3840
rect 2998 3780 3002 3836
rect 3002 3780 3058 3836
rect 3058 3780 3062 3836
rect 2998 3776 3062 3780
rect 3078 3836 3142 3840
rect 3078 3780 3082 3836
rect 3082 3780 3138 3836
rect 3138 3780 3142 3836
rect 3078 3776 3142 3780
rect 3158 3836 3222 3840
rect 3158 3780 3162 3836
rect 3162 3780 3218 3836
rect 3218 3780 3222 3836
rect 3158 3776 3222 3780
rect 6851 3836 6915 3840
rect 6851 3780 6855 3836
rect 6855 3780 6911 3836
rect 6911 3780 6915 3836
rect 6851 3776 6915 3780
rect 6931 3836 6995 3840
rect 6931 3780 6935 3836
rect 6935 3780 6991 3836
rect 6991 3780 6995 3836
rect 6931 3776 6995 3780
rect 7011 3836 7075 3840
rect 7011 3780 7015 3836
rect 7015 3780 7071 3836
rect 7071 3780 7075 3836
rect 7011 3776 7075 3780
rect 7091 3836 7155 3840
rect 7091 3780 7095 3836
rect 7095 3780 7151 3836
rect 7151 3780 7155 3836
rect 7091 3776 7155 3780
rect 10784 3836 10848 3840
rect 10784 3780 10788 3836
rect 10788 3780 10844 3836
rect 10844 3780 10848 3836
rect 10784 3776 10848 3780
rect 10864 3836 10928 3840
rect 10864 3780 10868 3836
rect 10868 3780 10924 3836
rect 10924 3780 10928 3836
rect 10864 3776 10928 3780
rect 10944 3836 11008 3840
rect 10944 3780 10948 3836
rect 10948 3780 11004 3836
rect 11004 3780 11008 3836
rect 10944 3776 11008 3780
rect 11024 3836 11088 3840
rect 11024 3780 11028 3836
rect 11028 3780 11084 3836
rect 11084 3780 11088 3836
rect 11024 3776 11088 3780
rect 14717 3836 14781 3840
rect 14717 3780 14721 3836
rect 14721 3780 14777 3836
rect 14777 3780 14781 3836
rect 14717 3776 14781 3780
rect 14797 3836 14861 3840
rect 14797 3780 14801 3836
rect 14801 3780 14857 3836
rect 14857 3780 14861 3836
rect 14797 3776 14861 3780
rect 14877 3836 14941 3840
rect 14877 3780 14881 3836
rect 14881 3780 14937 3836
rect 14937 3780 14941 3836
rect 14877 3776 14941 3780
rect 14957 3836 15021 3840
rect 14957 3780 14961 3836
rect 14961 3780 15017 3836
rect 15017 3780 15021 3836
rect 14957 3776 15021 3780
rect 4884 3292 4948 3296
rect 4884 3236 4888 3292
rect 4888 3236 4944 3292
rect 4944 3236 4948 3292
rect 4884 3232 4948 3236
rect 4964 3292 5028 3296
rect 4964 3236 4968 3292
rect 4968 3236 5024 3292
rect 5024 3236 5028 3292
rect 4964 3232 5028 3236
rect 5044 3292 5108 3296
rect 5044 3236 5048 3292
rect 5048 3236 5104 3292
rect 5104 3236 5108 3292
rect 5044 3232 5108 3236
rect 5124 3292 5188 3296
rect 5124 3236 5128 3292
rect 5128 3236 5184 3292
rect 5184 3236 5188 3292
rect 5124 3232 5188 3236
rect 8817 3292 8881 3296
rect 8817 3236 8821 3292
rect 8821 3236 8877 3292
rect 8877 3236 8881 3292
rect 8817 3232 8881 3236
rect 8897 3292 8961 3296
rect 8897 3236 8901 3292
rect 8901 3236 8957 3292
rect 8957 3236 8961 3292
rect 8897 3232 8961 3236
rect 8977 3292 9041 3296
rect 8977 3236 8981 3292
rect 8981 3236 9037 3292
rect 9037 3236 9041 3292
rect 8977 3232 9041 3236
rect 9057 3292 9121 3296
rect 9057 3236 9061 3292
rect 9061 3236 9117 3292
rect 9117 3236 9121 3292
rect 9057 3232 9121 3236
rect 12750 3292 12814 3296
rect 12750 3236 12754 3292
rect 12754 3236 12810 3292
rect 12810 3236 12814 3292
rect 12750 3232 12814 3236
rect 12830 3292 12894 3296
rect 12830 3236 12834 3292
rect 12834 3236 12890 3292
rect 12890 3236 12894 3292
rect 12830 3232 12894 3236
rect 12910 3292 12974 3296
rect 12910 3236 12914 3292
rect 12914 3236 12970 3292
rect 12970 3236 12974 3292
rect 12910 3232 12974 3236
rect 12990 3292 13054 3296
rect 12990 3236 12994 3292
rect 12994 3236 13050 3292
rect 13050 3236 13054 3292
rect 12990 3232 13054 3236
rect 16683 3292 16747 3296
rect 16683 3236 16687 3292
rect 16687 3236 16743 3292
rect 16743 3236 16747 3292
rect 16683 3232 16747 3236
rect 16763 3292 16827 3296
rect 16763 3236 16767 3292
rect 16767 3236 16823 3292
rect 16823 3236 16827 3292
rect 16763 3232 16827 3236
rect 16843 3292 16907 3296
rect 16843 3236 16847 3292
rect 16847 3236 16903 3292
rect 16903 3236 16907 3292
rect 16843 3232 16907 3236
rect 16923 3292 16987 3296
rect 16923 3236 16927 3292
rect 16927 3236 16983 3292
rect 16983 3236 16987 3292
rect 16923 3232 16987 3236
rect 2918 2748 2982 2752
rect 2918 2692 2922 2748
rect 2922 2692 2978 2748
rect 2978 2692 2982 2748
rect 2918 2688 2982 2692
rect 2998 2748 3062 2752
rect 2998 2692 3002 2748
rect 3002 2692 3058 2748
rect 3058 2692 3062 2748
rect 2998 2688 3062 2692
rect 3078 2748 3142 2752
rect 3078 2692 3082 2748
rect 3082 2692 3138 2748
rect 3138 2692 3142 2748
rect 3078 2688 3142 2692
rect 3158 2748 3222 2752
rect 3158 2692 3162 2748
rect 3162 2692 3218 2748
rect 3218 2692 3222 2748
rect 3158 2688 3222 2692
rect 6851 2748 6915 2752
rect 6851 2692 6855 2748
rect 6855 2692 6911 2748
rect 6911 2692 6915 2748
rect 6851 2688 6915 2692
rect 6931 2748 6995 2752
rect 6931 2692 6935 2748
rect 6935 2692 6991 2748
rect 6991 2692 6995 2748
rect 6931 2688 6995 2692
rect 7011 2748 7075 2752
rect 7011 2692 7015 2748
rect 7015 2692 7071 2748
rect 7071 2692 7075 2748
rect 7011 2688 7075 2692
rect 7091 2748 7155 2752
rect 7091 2692 7095 2748
rect 7095 2692 7151 2748
rect 7151 2692 7155 2748
rect 7091 2688 7155 2692
rect 10784 2748 10848 2752
rect 10784 2692 10788 2748
rect 10788 2692 10844 2748
rect 10844 2692 10848 2748
rect 10784 2688 10848 2692
rect 10864 2748 10928 2752
rect 10864 2692 10868 2748
rect 10868 2692 10924 2748
rect 10924 2692 10928 2748
rect 10864 2688 10928 2692
rect 10944 2748 11008 2752
rect 10944 2692 10948 2748
rect 10948 2692 11004 2748
rect 11004 2692 11008 2748
rect 10944 2688 11008 2692
rect 11024 2748 11088 2752
rect 11024 2692 11028 2748
rect 11028 2692 11084 2748
rect 11084 2692 11088 2748
rect 11024 2688 11088 2692
rect 14717 2748 14781 2752
rect 14717 2692 14721 2748
rect 14721 2692 14777 2748
rect 14777 2692 14781 2748
rect 14717 2688 14781 2692
rect 14797 2748 14861 2752
rect 14797 2692 14801 2748
rect 14801 2692 14857 2748
rect 14857 2692 14861 2748
rect 14797 2688 14861 2692
rect 14877 2748 14941 2752
rect 14877 2692 14881 2748
rect 14881 2692 14937 2748
rect 14937 2692 14941 2748
rect 14877 2688 14941 2692
rect 14957 2748 15021 2752
rect 14957 2692 14961 2748
rect 14961 2692 15017 2748
rect 15017 2692 15021 2748
rect 14957 2688 15021 2692
rect 14228 2620 14292 2684
rect 4884 2204 4948 2208
rect 4884 2148 4888 2204
rect 4888 2148 4944 2204
rect 4944 2148 4948 2204
rect 4884 2144 4948 2148
rect 4964 2204 5028 2208
rect 4964 2148 4968 2204
rect 4968 2148 5024 2204
rect 5024 2148 5028 2204
rect 4964 2144 5028 2148
rect 5044 2204 5108 2208
rect 5044 2148 5048 2204
rect 5048 2148 5104 2204
rect 5104 2148 5108 2204
rect 5044 2144 5108 2148
rect 5124 2204 5188 2208
rect 5124 2148 5128 2204
rect 5128 2148 5184 2204
rect 5184 2148 5188 2204
rect 5124 2144 5188 2148
rect 8817 2204 8881 2208
rect 8817 2148 8821 2204
rect 8821 2148 8877 2204
rect 8877 2148 8881 2204
rect 8817 2144 8881 2148
rect 8897 2204 8961 2208
rect 8897 2148 8901 2204
rect 8901 2148 8957 2204
rect 8957 2148 8961 2204
rect 8897 2144 8961 2148
rect 8977 2204 9041 2208
rect 8977 2148 8981 2204
rect 8981 2148 9037 2204
rect 9037 2148 9041 2204
rect 8977 2144 9041 2148
rect 9057 2204 9121 2208
rect 9057 2148 9061 2204
rect 9061 2148 9117 2204
rect 9117 2148 9121 2204
rect 9057 2144 9121 2148
rect 12750 2204 12814 2208
rect 12750 2148 12754 2204
rect 12754 2148 12810 2204
rect 12810 2148 12814 2204
rect 12750 2144 12814 2148
rect 12830 2204 12894 2208
rect 12830 2148 12834 2204
rect 12834 2148 12890 2204
rect 12890 2148 12894 2204
rect 12830 2144 12894 2148
rect 12910 2204 12974 2208
rect 12910 2148 12914 2204
rect 12914 2148 12970 2204
rect 12970 2148 12974 2204
rect 12910 2144 12974 2148
rect 12990 2204 13054 2208
rect 12990 2148 12994 2204
rect 12994 2148 13050 2204
rect 13050 2148 13054 2204
rect 12990 2144 13054 2148
rect 16683 2204 16747 2208
rect 16683 2148 16687 2204
rect 16687 2148 16743 2204
rect 16743 2148 16747 2204
rect 16683 2144 16747 2148
rect 16763 2204 16827 2208
rect 16763 2148 16767 2204
rect 16767 2148 16823 2204
rect 16823 2148 16827 2204
rect 16763 2144 16827 2148
rect 16843 2204 16907 2208
rect 16843 2148 16847 2204
rect 16847 2148 16903 2204
rect 16903 2148 16907 2204
rect 16843 2144 16907 2148
rect 16923 2204 16987 2208
rect 16923 2148 16927 2204
rect 16927 2148 16983 2204
rect 16983 2148 16987 2204
rect 16923 2144 16987 2148
<< metal4 >>
rect 2910 15808 3230 15824
rect 2910 15744 2918 15808
rect 2982 15744 2998 15808
rect 3062 15744 3078 15808
rect 3142 15744 3158 15808
rect 3222 15744 3230 15808
rect 2910 14720 3230 15744
rect 2910 14656 2918 14720
rect 2982 14656 2998 14720
rect 3062 14656 3078 14720
rect 3142 14656 3158 14720
rect 3222 14656 3230 14720
rect 2910 13632 3230 14656
rect 2910 13568 2918 13632
rect 2982 13568 2998 13632
rect 3062 13568 3078 13632
rect 3142 13568 3158 13632
rect 3222 13568 3230 13632
rect 2910 12544 3230 13568
rect 2910 12480 2918 12544
rect 2982 12480 2998 12544
rect 3062 12480 3078 12544
rect 3142 12480 3158 12544
rect 3222 12480 3230 12544
rect 2910 11456 3230 12480
rect 2910 11392 2918 11456
rect 2982 11392 2998 11456
rect 3062 11392 3078 11456
rect 3142 11392 3158 11456
rect 3222 11392 3230 11456
rect 2910 10368 3230 11392
rect 2910 10304 2918 10368
rect 2982 10304 2998 10368
rect 3062 10304 3078 10368
rect 3142 10304 3158 10368
rect 3222 10304 3230 10368
rect 2910 9280 3230 10304
rect 2910 9216 2918 9280
rect 2982 9216 2998 9280
rect 3062 9216 3078 9280
rect 3142 9216 3158 9280
rect 3222 9216 3230 9280
rect 2910 8192 3230 9216
rect 2910 8128 2918 8192
rect 2982 8128 2998 8192
rect 3062 8128 3078 8192
rect 3142 8128 3158 8192
rect 3222 8128 3230 8192
rect 2910 7104 3230 8128
rect 2910 7040 2918 7104
rect 2982 7040 2998 7104
rect 3062 7040 3078 7104
rect 3142 7040 3158 7104
rect 3222 7040 3230 7104
rect 2910 6016 3230 7040
rect 2910 5952 2918 6016
rect 2982 5952 2998 6016
rect 3062 5952 3078 6016
rect 3142 5952 3158 6016
rect 3222 5952 3230 6016
rect 2910 4928 3230 5952
rect 2910 4864 2918 4928
rect 2982 4864 2998 4928
rect 3062 4864 3078 4928
rect 3142 4864 3158 4928
rect 3222 4864 3230 4928
rect 2910 3840 3230 4864
rect 2910 3776 2918 3840
rect 2982 3776 2998 3840
rect 3062 3776 3078 3840
rect 3142 3776 3158 3840
rect 3222 3776 3230 3840
rect 2910 2752 3230 3776
rect 2910 2688 2918 2752
rect 2982 2688 2998 2752
rect 3062 2688 3078 2752
rect 3142 2688 3158 2752
rect 3222 2688 3230 2752
rect 2910 2128 3230 2688
rect 4876 15264 5196 15824
rect 4876 15200 4884 15264
rect 4948 15200 4964 15264
rect 5028 15200 5044 15264
rect 5108 15200 5124 15264
rect 5188 15200 5196 15264
rect 4876 14176 5196 15200
rect 4876 14112 4884 14176
rect 4948 14112 4964 14176
rect 5028 14112 5044 14176
rect 5108 14112 5124 14176
rect 5188 14112 5196 14176
rect 4876 13088 5196 14112
rect 4876 13024 4884 13088
rect 4948 13024 4964 13088
rect 5028 13024 5044 13088
rect 5108 13024 5124 13088
rect 5188 13024 5196 13088
rect 4876 12000 5196 13024
rect 4876 11936 4884 12000
rect 4948 11936 4964 12000
rect 5028 11936 5044 12000
rect 5108 11936 5124 12000
rect 5188 11936 5196 12000
rect 4876 10912 5196 11936
rect 4876 10848 4884 10912
rect 4948 10848 4964 10912
rect 5028 10848 5044 10912
rect 5108 10848 5124 10912
rect 5188 10848 5196 10912
rect 4876 9824 5196 10848
rect 4876 9760 4884 9824
rect 4948 9760 4964 9824
rect 5028 9760 5044 9824
rect 5108 9760 5124 9824
rect 5188 9760 5196 9824
rect 4876 8736 5196 9760
rect 4876 8672 4884 8736
rect 4948 8672 4964 8736
rect 5028 8672 5044 8736
rect 5108 8672 5124 8736
rect 5188 8672 5196 8736
rect 4876 7648 5196 8672
rect 4876 7584 4884 7648
rect 4948 7584 4964 7648
rect 5028 7584 5044 7648
rect 5108 7584 5124 7648
rect 5188 7584 5196 7648
rect 4876 6560 5196 7584
rect 4876 6496 4884 6560
rect 4948 6496 4964 6560
rect 5028 6496 5044 6560
rect 5108 6496 5124 6560
rect 5188 6496 5196 6560
rect 4876 5472 5196 6496
rect 4876 5408 4884 5472
rect 4948 5408 4964 5472
rect 5028 5408 5044 5472
rect 5108 5408 5124 5472
rect 5188 5408 5196 5472
rect 4876 4384 5196 5408
rect 4876 4320 4884 4384
rect 4948 4320 4964 4384
rect 5028 4320 5044 4384
rect 5108 4320 5124 4384
rect 5188 4320 5196 4384
rect 4876 3296 5196 4320
rect 4876 3232 4884 3296
rect 4948 3232 4964 3296
rect 5028 3232 5044 3296
rect 5108 3232 5124 3296
rect 5188 3232 5196 3296
rect 4876 2208 5196 3232
rect 4876 2144 4884 2208
rect 4948 2144 4964 2208
rect 5028 2144 5044 2208
rect 5108 2144 5124 2208
rect 5188 2144 5196 2208
rect 4876 2128 5196 2144
rect 6843 15808 7163 15824
rect 6843 15744 6851 15808
rect 6915 15744 6931 15808
rect 6995 15744 7011 15808
rect 7075 15744 7091 15808
rect 7155 15744 7163 15808
rect 6843 14720 7163 15744
rect 6843 14656 6851 14720
rect 6915 14656 6931 14720
rect 6995 14656 7011 14720
rect 7075 14656 7091 14720
rect 7155 14656 7163 14720
rect 6843 13632 7163 14656
rect 6843 13568 6851 13632
rect 6915 13568 6931 13632
rect 6995 13568 7011 13632
rect 7075 13568 7091 13632
rect 7155 13568 7163 13632
rect 6843 12544 7163 13568
rect 6843 12480 6851 12544
rect 6915 12480 6931 12544
rect 6995 12480 7011 12544
rect 7075 12480 7091 12544
rect 7155 12480 7163 12544
rect 6843 11456 7163 12480
rect 6843 11392 6851 11456
rect 6915 11392 6931 11456
rect 6995 11392 7011 11456
rect 7075 11392 7091 11456
rect 7155 11392 7163 11456
rect 6843 10368 7163 11392
rect 6843 10304 6851 10368
rect 6915 10304 6931 10368
rect 6995 10304 7011 10368
rect 7075 10304 7091 10368
rect 7155 10304 7163 10368
rect 6843 9280 7163 10304
rect 6843 9216 6851 9280
rect 6915 9216 6931 9280
rect 6995 9216 7011 9280
rect 7075 9216 7091 9280
rect 7155 9216 7163 9280
rect 6843 8192 7163 9216
rect 6843 8128 6851 8192
rect 6915 8128 6931 8192
rect 6995 8128 7011 8192
rect 7075 8128 7091 8192
rect 7155 8128 7163 8192
rect 6843 7104 7163 8128
rect 6843 7040 6851 7104
rect 6915 7040 6931 7104
rect 6995 7040 7011 7104
rect 7075 7040 7091 7104
rect 7155 7040 7163 7104
rect 6843 6016 7163 7040
rect 6843 5952 6851 6016
rect 6915 5952 6931 6016
rect 6995 5952 7011 6016
rect 7075 5952 7091 6016
rect 7155 5952 7163 6016
rect 6843 4928 7163 5952
rect 6843 4864 6851 4928
rect 6915 4864 6931 4928
rect 6995 4864 7011 4928
rect 7075 4864 7091 4928
rect 7155 4864 7163 4928
rect 6843 3840 7163 4864
rect 6843 3776 6851 3840
rect 6915 3776 6931 3840
rect 6995 3776 7011 3840
rect 7075 3776 7091 3840
rect 7155 3776 7163 3840
rect 6843 2752 7163 3776
rect 6843 2688 6851 2752
rect 6915 2688 6931 2752
rect 6995 2688 7011 2752
rect 7075 2688 7091 2752
rect 7155 2688 7163 2752
rect 6843 2128 7163 2688
rect 8809 15264 9129 15824
rect 8809 15200 8817 15264
rect 8881 15200 8897 15264
rect 8961 15200 8977 15264
rect 9041 15200 9057 15264
rect 9121 15200 9129 15264
rect 8809 14176 9129 15200
rect 8809 14112 8817 14176
rect 8881 14112 8897 14176
rect 8961 14112 8977 14176
rect 9041 14112 9057 14176
rect 9121 14112 9129 14176
rect 8809 13088 9129 14112
rect 8809 13024 8817 13088
rect 8881 13024 8897 13088
rect 8961 13024 8977 13088
rect 9041 13024 9057 13088
rect 9121 13024 9129 13088
rect 8809 12000 9129 13024
rect 8809 11936 8817 12000
rect 8881 11936 8897 12000
rect 8961 11936 8977 12000
rect 9041 11936 9057 12000
rect 9121 11936 9129 12000
rect 8809 10912 9129 11936
rect 8809 10848 8817 10912
rect 8881 10848 8897 10912
rect 8961 10848 8977 10912
rect 9041 10848 9057 10912
rect 9121 10848 9129 10912
rect 8809 9824 9129 10848
rect 8809 9760 8817 9824
rect 8881 9760 8897 9824
rect 8961 9760 8977 9824
rect 9041 9760 9057 9824
rect 9121 9760 9129 9824
rect 8809 8736 9129 9760
rect 8809 8672 8817 8736
rect 8881 8672 8897 8736
rect 8961 8672 8977 8736
rect 9041 8672 9057 8736
rect 9121 8672 9129 8736
rect 8809 7648 9129 8672
rect 8809 7584 8817 7648
rect 8881 7584 8897 7648
rect 8961 7584 8977 7648
rect 9041 7584 9057 7648
rect 9121 7584 9129 7648
rect 8809 6560 9129 7584
rect 8809 6496 8817 6560
rect 8881 6496 8897 6560
rect 8961 6496 8977 6560
rect 9041 6496 9057 6560
rect 9121 6496 9129 6560
rect 8809 5472 9129 6496
rect 8809 5408 8817 5472
rect 8881 5408 8897 5472
rect 8961 5408 8977 5472
rect 9041 5408 9057 5472
rect 9121 5408 9129 5472
rect 8809 4384 9129 5408
rect 8809 4320 8817 4384
rect 8881 4320 8897 4384
rect 8961 4320 8977 4384
rect 9041 4320 9057 4384
rect 9121 4320 9129 4384
rect 8809 3296 9129 4320
rect 8809 3232 8817 3296
rect 8881 3232 8897 3296
rect 8961 3232 8977 3296
rect 9041 3232 9057 3296
rect 9121 3232 9129 3296
rect 8809 2208 9129 3232
rect 8809 2144 8817 2208
rect 8881 2144 8897 2208
rect 8961 2144 8977 2208
rect 9041 2144 9057 2208
rect 9121 2144 9129 2208
rect 8809 2128 9129 2144
rect 10776 15808 11096 15824
rect 10776 15744 10784 15808
rect 10848 15744 10864 15808
rect 10928 15744 10944 15808
rect 11008 15744 11024 15808
rect 11088 15744 11096 15808
rect 10776 14720 11096 15744
rect 10776 14656 10784 14720
rect 10848 14656 10864 14720
rect 10928 14656 10944 14720
rect 11008 14656 11024 14720
rect 11088 14656 11096 14720
rect 10776 13632 11096 14656
rect 10776 13568 10784 13632
rect 10848 13568 10864 13632
rect 10928 13568 10944 13632
rect 11008 13568 11024 13632
rect 11088 13568 11096 13632
rect 10776 12544 11096 13568
rect 10776 12480 10784 12544
rect 10848 12480 10864 12544
rect 10928 12480 10944 12544
rect 11008 12480 11024 12544
rect 11088 12480 11096 12544
rect 10776 11456 11096 12480
rect 10776 11392 10784 11456
rect 10848 11392 10864 11456
rect 10928 11392 10944 11456
rect 11008 11392 11024 11456
rect 11088 11392 11096 11456
rect 10776 10368 11096 11392
rect 12742 15264 13062 15824
rect 12742 15200 12750 15264
rect 12814 15200 12830 15264
rect 12894 15200 12910 15264
rect 12974 15200 12990 15264
rect 13054 15200 13062 15264
rect 12742 14176 13062 15200
rect 12742 14112 12750 14176
rect 12814 14112 12830 14176
rect 12894 14112 12910 14176
rect 12974 14112 12990 14176
rect 13054 14112 13062 14176
rect 12742 13088 13062 14112
rect 12742 13024 12750 13088
rect 12814 13024 12830 13088
rect 12894 13024 12910 13088
rect 12974 13024 12990 13088
rect 13054 13024 13062 13088
rect 12742 12000 13062 13024
rect 12742 11936 12750 12000
rect 12814 11936 12830 12000
rect 12894 11936 12910 12000
rect 12974 11936 12990 12000
rect 13054 11936 13062 12000
rect 11283 11116 11349 11117
rect 11283 11052 11284 11116
rect 11348 11052 11349 11116
rect 11283 11051 11349 11052
rect 10776 10304 10784 10368
rect 10848 10304 10864 10368
rect 10928 10304 10944 10368
rect 11008 10304 11024 10368
rect 11088 10304 11096 10368
rect 10776 9280 11096 10304
rect 10776 9216 10784 9280
rect 10848 9216 10864 9280
rect 10928 9216 10944 9280
rect 11008 9216 11024 9280
rect 11088 9216 11096 9280
rect 10776 8192 11096 9216
rect 10776 8128 10784 8192
rect 10848 8128 10864 8192
rect 10928 8128 10944 8192
rect 11008 8128 11024 8192
rect 11088 8128 11096 8192
rect 10776 7104 11096 8128
rect 10776 7040 10784 7104
rect 10848 7040 10864 7104
rect 10928 7040 10944 7104
rect 11008 7040 11024 7104
rect 11088 7040 11096 7104
rect 10776 6016 11096 7040
rect 10776 5952 10784 6016
rect 10848 5952 10864 6016
rect 10928 5952 10944 6016
rect 11008 5952 11024 6016
rect 11088 5952 11096 6016
rect 10776 4928 11096 5952
rect 11286 5541 11346 11051
rect 12742 10912 13062 11936
rect 14709 15808 15029 15824
rect 14709 15744 14717 15808
rect 14781 15744 14797 15808
rect 14861 15744 14877 15808
rect 14941 15744 14957 15808
rect 15021 15744 15029 15808
rect 14709 14720 15029 15744
rect 14709 14656 14717 14720
rect 14781 14656 14797 14720
rect 14861 14656 14877 14720
rect 14941 14656 14957 14720
rect 15021 14656 15029 14720
rect 14709 13632 15029 14656
rect 14709 13568 14717 13632
rect 14781 13568 14797 13632
rect 14861 13568 14877 13632
rect 14941 13568 14957 13632
rect 15021 13568 15029 13632
rect 14709 12544 15029 13568
rect 14709 12480 14717 12544
rect 14781 12480 14797 12544
rect 14861 12480 14877 12544
rect 14941 12480 14957 12544
rect 15021 12480 15029 12544
rect 14709 11456 15029 12480
rect 14709 11392 14717 11456
rect 14781 11392 14797 11456
rect 14861 11392 14877 11456
rect 14941 11392 14957 11456
rect 15021 11392 15029 11456
rect 14227 11116 14293 11117
rect 14227 11052 14228 11116
rect 14292 11052 14293 11116
rect 14227 11051 14293 11052
rect 12742 10848 12750 10912
rect 12814 10848 12830 10912
rect 12894 10848 12910 10912
rect 12974 10848 12990 10912
rect 13054 10848 13062 10912
rect 12742 9824 13062 10848
rect 12742 9760 12750 9824
rect 12814 9760 12830 9824
rect 12894 9760 12910 9824
rect 12974 9760 12990 9824
rect 13054 9760 13062 9824
rect 12742 8736 13062 9760
rect 12742 8672 12750 8736
rect 12814 8672 12830 8736
rect 12894 8672 12910 8736
rect 12974 8672 12990 8736
rect 13054 8672 13062 8736
rect 12742 7648 13062 8672
rect 12742 7584 12750 7648
rect 12814 7584 12830 7648
rect 12894 7584 12910 7648
rect 12974 7584 12990 7648
rect 13054 7584 13062 7648
rect 12742 6560 13062 7584
rect 12742 6496 12750 6560
rect 12814 6496 12830 6560
rect 12894 6496 12910 6560
rect 12974 6496 12990 6560
rect 13054 6496 13062 6560
rect 11283 5540 11349 5541
rect 11283 5476 11284 5540
rect 11348 5476 11349 5540
rect 11283 5475 11349 5476
rect 10776 4864 10784 4928
rect 10848 4864 10864 4928
rect 10928 4864 10944 4928
rect 11008 4864 11024 4928
rect 11088 4864 11096 4928
rect 10776 3840 11096 4864
rect 10776 3776 10784 3840
rect 10848 3776 10864 3840
rect 10928 3776 10944 3840
rect 11008 3776 11024 3840
rect 11088 3776 11096 3840
rect 10776 2752 11096 3776
rect 10776 2688 10784 2752
rect 10848 2688 10864 2752
rect 10928 2688 10944 2752
rect 11008 2688 11024 2752
rect 11088 2688 11096 2752
rect 10776 2128 11096 2688
rect 12742 5472 13062 6496
rect 12742 5408 12750 5472
rect 12814 5408 12830 5472
rect 12894 5408 12910 5472
rect 12974 5408 12990 5472
rect 13054 5408 13062 5472
rect 12742 4384 13062 5408
rect 12742 4320 12750 4384
rect 12814 4320 12830 4384
rect 12894 4320 12910 4384
rect 12974 4320 12990 4384
rect 13054 4320 13062 4384
rect 12742 3296 13062 4320
rect 12742 3232 12750 3296
rect 12814 3232 12830 3296
rect 12894 3232 12910 3296
rect 12974 3232 12990 3296
rect 13054 3232 13062 3296
rect 12742 2208 13062 3232
rect 14230 2685 14290 11051
rect 14411 10572 14477 10573
rect 14411 10508 14412 10572
rect 14476 10508 14477 10572
rect 14411 10507 14477 10508
rect 14414 4045 14474 10507
rect 14709 10368 15029 11392
rect 14709 10304 14717 10368
rect 14781 10304 14797 10368
rect 14861 10304 14877 10368
rect 14941 10304 14957 10368
rect 15021 10304 15029 10368
rect 14709 9280 15029 10304
rect 16675 15264 16995 15824
rect 16675 15200 16683 15264
rect 16747 15200 16763 15264
rect 16827 15200 16843 15264
rect 16907 15200 16923 15264
rect 16987 15200 16995 15264
rect 16675 14176 16995 15200
rect 16675 14112 16683 14176
rect 16747 14112 16763 14176
rect 16827 14112 16843 14176
rect 16907 14112 16923 14176
rect 16987 14112 16995 14176
rect 16675 13088 16995 14112
rect 16675 13024 16683 13088
rect 16747 13024 16763 13088
rect 16827 13024 16843 13088
rect 16907 13024 16923 13088
rect 16987 13024 16995 13088
rect 16675 12000 16995 13024
rect 16675 11936 16683 12000
rect 16747 11936 16763 12000
rect 16827 11936 16843 12000
rect 16907 11936 16923 12000
rect 16987 11936 16995 12000
rect 16675 10912 16995 11936
rect 16675 10848 16683 10912
rect 16747 10848 16763 10912
rect 16827 10848 16843 10912
rect 16907 10848 16923 10912
rect 16987 10848 16995 10912
rect 16675 9824 16995 10848
rect 16675 9760 16683 9824
rect 16747 9760 16763 9824
rect 16827 9760 16843 9824
rect 16907 9760 16923 9824
rect 16987 9760 16995 9824
rect 16251 9756 16317 9757
rect 16251 9692 16252 9756
rect 16316 9692 16317 9756
rect 16251 9691 16317 9692
rect 14709 9216 14717 9280
rect 14781 9216 14797 9280
rect 14861 9216 14877 9280
rect 14941 9216 14957 9280
rect 15021 9216 15029 9280
rect 14709 8192 15029 9216
rect 14709 8128 14717 8192
rect 14781 8128 14797 8192
rect 14861 8128 14877 8192
rect 14941 8128 14957 8192
rect 15021 8128 15029 8192
rect 14709 7104 15029 8128
rect 14709 7040 14717 7104
rect 14781 7040 14797 7104
rect 14861 7040 14877 7104
rect 14941 7040 14957 7104
rect 15021 7040 15029 7104
rect 14709 6016 15029 7040
rect 14709 5952 14717 6016
rect 14781 5952 14797 6016
rect 14861 5952 14877 6016
rect 14941 5952 14957 6016
rect 15021 5952 15029 6016
rect 14709 4928 15029 5952
rect 14709 4864 14717 4928
rect 14781 4864 14797 4928
rect 14861 4864 14877 4928
rect 14941 4864 14957 4928
rect 15021 4864 15029 4928
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 14709 3840 15029 4864
rect 16254 4045 16314 9691
rect 16675 8736 16995 9760
rect 16675 8672 16683 8736
rect 16747 8672 16763 8736
rect 16827 8672 16843 8736
rect 16907 8672 16923 8736
rect 16987 8672 16995 8736
rect 16675 7648 16995 8672
rect 16675 7584 16683 7648
rect 16747 7584 16763 7648
rect 16827 7584 16843 7648
rect 16907 7584 16923 7648
rect 16987 7584 16995 7648
rect 16675 6560 16995 7584
rect 16675 6496 16683 6560
rect 16747 6496 16763 6560
rect 16827 6496 16843 6560
rect 16907 6496 16923 6560
rect 16987 6496 16995 6560
rect 16675 5472 16995 6496
rect 16675 5408 16683 5472
rect 16747 5408 16763 5472
rect 16827 5408 16843 5472
rect 16907 5408 16923 5472
rect 16987 5408 16995 5472
rect 16675 4384 16995 5408
rect 16675 4320 16683 4384
rect 16747 4320 16763 4384
rect 16827 4320 16843 4384
rect 16907 4320 16923 4384
rect 16987 4320 16995 4384
rect 16251 4044 16317 4045
rect 16251 3980 16252 4044
rect 16316 3980 16317 4044
rect 16251 3979 16317 3980
rect 14709 3776 14717 3840
rect 14781 3776 14797 3840
rect 14861 3776 14877 3840
rect 14941 3776 14957 3840
rect 15021 3776 15029 3840
rect 14709 2752 15029 3776
rect 14709 2688 14717 2752
rect 14781 2688 14797 2752
rect 14861 2688 14877 2752
rect 14941 2688 14957 2752
rect 15021 2688 15029 2752
rect 14227 2684 14293 2685
rect 14227 2620 14228 2684
rect 14292 2620 14293 2684
rect 14227 2619 14293 2620
rect 12742 2144 12750 2208
rect 12814 2144 12830 2208
rect 12894 2144 12910 2208
rect 12974 2144 12990 2208
rect 13054 2144 13062 2208
rect 12742 2128 13062 2144
rect 14709 2128 15029 2688
rect 16675 3296 16995 4320
rect 16675 3232 16683 3296
rect 16747 3232 16763 3296
rect 16827 3232 16843 3296
rect 16907 3232 16923 3296
rect 16987 3232 16995 3296
rect 16675 2208 16995 3232
rect 16675 2144 16683 2208
rect 16747 2144 16763 2208
rect 16827 2144 16843 2208
rect 16907 2144 16923 2208
rect 16987 2144 16995 2208
rect 16675 2128 16995 2144
use sky130_fd_sc_hd__inv_2  _172_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1688980957
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1688980957
transform -1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1688980957
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1688980957
transform -1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1688980957
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1688980957
transform -1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1688980957
transform -1 0 15640 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1688980957
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1688980957
transform -1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1688980957
transform -1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1688980957
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1688980957
transform -1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1688980957
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1688980957
transform -1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1688980957
transform -1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1688980957
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1688980957
transform -1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1688980957
transform -1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1688980957
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1688980957
transform -1 0 6256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform -1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1688980957
transform -1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1688980957
transform -1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1688980957
transform -1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1688980957
transform -1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform -1 0 13892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1688980957
transform -1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1688980957
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1688980957
transform -1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1688980957
transform 1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1688980957
transform -1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1688980957
transform -1 0 10580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1688980957
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1688980957
transform -1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1688980957
transform -1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1688980957
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1688980957
transform -1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1688980957
transform 1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1688980957
transform -1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1688980957
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1688980957
transform -1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1688980957
transform 1 0 14352 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1688980957
transform 1 0 11592 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1688980957
transform 1 0 12144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1688980957
transform -1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1688980957
transform -1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1688980957
transform -1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1688980957
transform -1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1688980957
transform -1 0 15180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _239_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1688980957
transform -1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform -1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1688980957
transform -1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform -1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform -1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1688980957
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1688980957
transform -1 0 6256 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1688980957
transform -1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1688980957
transform -1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1688980957
transform -1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1688980957
transform -1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1688980957
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1688980957
transform -1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1688980957
transform -1 0 4508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1688980957
transform -1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1688980957
transform -1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1688980957
transform -1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1688980957
transform -1 0 8740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _267_
timestamp 1688980957
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1688980957
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1688980957
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1688980957
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1688980957
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1688980957
transform -1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _273_
timestamp 1688980957
transform -1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1688980957
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1688980957
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1688980957
transform -1 0 9200 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1688980957
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1688980957
transform -1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1688980957
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1688980957
transform 1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1688980957
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1688980957
transform -1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1688980957
transform -1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1688980957
transform 1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1688980957
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1688980957
transform -1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1688980957
transform -1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1688980957
transform -1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1688980957
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1688980957
transform -1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1688980957
transform -1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1688980957
transform -1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1688980957
transform -1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1688980957
transform -1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1688980957
transform -1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1688980957
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1688980957
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1688980957
transform -1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1688980957
transform -1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1688980957
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1688980957
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1688980957
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1688980957
transform -1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1688980957
transform -1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1688980957
transform -1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1688980957
transform -1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1688980957
transform -1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1688980957
transform -1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1688980957
transform -1 0 14720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1688980957
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1688980957
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1688980957
transform -1 0 11408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1688980957
transform -1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1688980957
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1688980957
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform -1 0 2668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1688980957
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1688980957
transform -1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1688980957
transform -1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1688980957
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform -1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1688980957
transform -1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1688980957
transform 1 0 4508 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform -1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1688980957
transform 1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1688980957
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1688980957
transform -1 0 13432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1688980957
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1688980957
transform 1 0 15640 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1688980957
transform -1 0 14904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1688980957
transform 1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1688980957
transform -1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1688980957
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1688980957
transform -1 0 15640 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1688980957
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1688980957
transform 1 0 9936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1688980957
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1688980957
transform -1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _376_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1688980957
transform -1 0 11960 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _378_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1688980957
transform -1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _381_
timestamp 1688980957
transform -1 0 13800 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1688980957
transform 1 0 9108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _384_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1688980957
transform -1 0 3864 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _387_
timestamp 1688980957
transform -1 0 10488 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1688980957
transform 1 0 14628 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1688980957
transform 1 0 12512 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1688980957
transform 1 0 9936 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1688980957
transform -1 0 8924 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1688980957
transform 1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1688980957
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1688980957
transform 1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1688980957
transform -1 0 13708 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1688980957
transform -1 0 16100 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1688980957
transform -1 0 12880 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1688980957
transform -1 0 13524 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1688980957
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1688980957
transform -1 0 7820 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _422_
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _423_
timestamp 1688980957
transform -1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _427_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1688980957
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _430_
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1688980957
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _435_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _436_
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _437_
timestamp 1688980957
transform -1 0 15456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _438_
timestamp 1688980957
transform -1 0 11224 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _439_
timestamp 1688980957
transform -1 0 14260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _440__63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _440_
timestamp 1688980957
transform -1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _441_
timestamp 1688980957
transform 1 0 10212 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _442_
timestamp 1688980957
transform -1 0 13524 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _443_
timestamp 1688980957
transform 1 0 11224 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _444_
timestamp 1688980957
transform -1 0 13340 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _445_
timestamp 1688980957
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _446_
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _447_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _448__64
timestamp 1688980957
transform -1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _448_
timestamp 1688980957
transform 1 0 4600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _449_
timestamp 1688980957
transform -1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _450_
timestamp 1688980957
transform -1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _451_
timestamp 1688980957
transform -1 0 15640 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _452_
timestamp 1688980957
transform -1 0 13248 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _453_
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _454_
timestamp 1688980957
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _455_
timestamp 1688980957
transform 1 0 4048 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _456_
timestamp 1688980957
transform -1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _457_
timestamp 1688980957
transform -1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _458_
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _459_
timestamp 1688980957
transform -1 0 11316 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _460__65
timestamp 1688980957
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _460_
timestamp 1688980957
transform -1 0 11316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _461_
timestamp 1688980957
transform -1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _462_
timestamp 1688980957
transform 1 0 14996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _463_
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _464_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _465_
timestamp 1688980957
transform -1 0 11316 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _466_
timestamp 1688980957
transform -1 0 11408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _467_
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _468_
timestamp 1688980957
transform -1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _469_
timestamp 1688980957
transform 1 0 15456 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _470_
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _471_
timestamp 1688980957
transform -1 0 5704 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _472__66
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _472_
timestamp 1688980957
transform 1 0 4048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _473_
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _474_
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _475_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _476_
timestamp 1688980957
transform -1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _477_
timestamp 1688980957
transform 1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _478_
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _479_
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _480_
timestamp 1688980957
transform -1 0 4600 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _481_
timestamp 1688980957
transform -1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _482_
timestamp 1688980957
transform -1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _483_
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _484__67
timestamp 1688980957
transform 1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _484_
timestamp 1688980957
transform -1 0 8280 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _485_
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _486_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _487_
timestamp 1688980957
transform -1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _488_
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _489_
timestamp 1688980957
transform -1 0 8648 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _490_
timestamp 1688980957
transform -1 0 8188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _491_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _492_
timestamp 1688980957
transform -1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _493_
timestamp 1688980957
transform -1 0 16468 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _494_
timestamp 1688980957
transform -1 0 16100 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _494__68
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _495_
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _496_
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _497_
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _498_
timestamp 1688980957
transform -1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _499_
timestamp 1688980957
transform -1 0 15364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _500_
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _501_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _502_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _503_
timestamp 1688980957
transform 1 0 9844 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _504__69
timestamp 1688980957
transform -1 0 9568 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _504_
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _505_
timestamp 1688980957
transform 1 0 7636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _506_
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _507_
timestamp 1688980957
transform -1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _508_
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _509_
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _510_
timestamp 1688980957
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _510__70
timestamp 1688980957
transform -1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _511_
timestamp 1688980957
transform -1 0 11316 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _512_
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _513_
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _514_
timestamp 1688980957
transform 1 0 10120 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _515_
timestamp 1688980957
transform 1 0 14444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _516__71
timestamp 1688980957
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _516_
timestamp 1688980957
transform 1 0 12696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _517_
timestamp 1688980957
transform -1 0 14720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _518_
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _519_
timestamp 1688980957
transform 1 0 11776 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _520_
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _521_
timestamp 1688980957
transform -1 0 13984 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _522__72
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _522_
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _523_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _524_
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _525_
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _526_
timestamp 1688980957
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _527_
timestamp 1688980957
transform 1 0 13156 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _528_
timestamp 1688980957
transform -1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _528__73
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _529_
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _530_
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _531_
timestamp 1688980957
transform -1 0 13524 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _532_
timestamp 1688980957
transform -1 0 12512 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _533__74
timestamp 1688980957
transform -1 0 15824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _533_
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _534_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _535_
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _536_
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _537__75
timestamp 1688980957
transform -1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _537_
timestamp 1688980957
transform 1 0 9016 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _538_
timestamp 1688980957
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _539_
timestamp 1688980957
transform 1 0 8188 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _540_
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1688980957
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1688980957
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1688980957
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_61
timestamp 1688980957
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_132
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_155
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_159
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1688980957
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_12
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_18
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_22
timestamp 1688980957
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_34
timestamp 1688980957
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_46
timestamp 1688980957
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_65
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_80
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 1688980957
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_136
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_150
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_163
timestamp 1688980957
transform 1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_32
timestamp 1688980957
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_44
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_56
timestamp 1688980957
transform 1 0 6256 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_107
timestamp 1688980957
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_124
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_150
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_160
timestamp 1688980957
transform 1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_21
timestamp 1688980957
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_33
timestamp 1688980957
transform 1 0 4140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_41
timestamp 1688980957
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_48
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_52
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp 1688980957
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_98
timestamp 1688980957
transform 1 0 10120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_154
timestamp 1688980957
transform 1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_55
timestamp 1688980957
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_80
timestamp 1688980957
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_167
timestamp 1688980957
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_103
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_119
timestamp 1688980957
transform 1 0 12052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_12
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_24
timestamp 1688980957
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_68
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_99
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_25
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_31
timestamp 1688980957
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_143
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_162
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_89
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_99
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_120
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_135
timestamp 1688980957
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_147
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_158
timestamp 1688980957
transform 1 0 15640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_167
timestamp 1688980957
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_17
timestamp 1688980957
transform 1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_41
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_12
timestamp 1688980957
transform 1 0 2208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_20
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_68
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_166
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_25
timestamp 1688980957
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_48
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_119
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_36
timestamp 1688980957
transform 1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_50
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_88
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_11
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_84
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_143
timestamp 1688980957
transform 1 0 14260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_163
timestamp 1688980957
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_55
timestamp 1688980957
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_99
timestamp 1688980957
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_167
timestamp 1688980957
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_68
timestamp 1688980957
transform 1 0 7360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_85
timestamp 1688980957
transform 1 0 8924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_117
timestamp 1688980957
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_121
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_140
timestamp 1688980957
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_157
timestamp 1688980957
transform 1 0 15548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_78
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_88
timestamp 1688980957
transform 1 0 9200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_104
timestamp 1688980957
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_108
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_112
timestamp 1688980957
transform 1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_116
timestamp 1688980957
transform 1 0 11776 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_126
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_166
timestamp 1688980957
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_83
timestamp 1688980957
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_127
timestamp 1688980957
transform 1 0 12788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_135
timestamp 1688980957
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_156
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_24
timestamp 1688980957
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_104
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_108
timestamp 1688980957
transform 1 0 11040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_112
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_12
timestamp 1688980957
transform 1 0 2208 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_24
timestamp 1688980957
transform 1 0 3312 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_36
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_40
timestamp 1688980957
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_44
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp 1688980957
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_153
timestamp 1688980957
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_124
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_167
timestamp 1688980957
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 1688980957
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_139
timestamp 1688980957
transform 1 0 13892 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_160
timestamp 1688980957
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_92
timestamp 1688980957
transform 1 0 9568 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_106
timestamp 1688980957
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_129
timestamp 1688980957
transform 1 0 12972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_161
timestamp 1688980957
transform 1 0 15916 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_9
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_17
timestamp 1688980957
transform 1 0 2668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_29
timestamp 1688980957
transform 1 0 3772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_41
timestamp 1688980957
transform 1 0 4876 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_45
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_72
timestamp 1688980957
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_84
timestamp 1688980957
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_99
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_129
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_141
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_17
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_24
timestamp 1688980957
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_38
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_50
timestamp 1688980957
transform 1 0 5704 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp 1688980957
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_57
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_72
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_101
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_106
timestamp 1688980957
transform 1 0 10856 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_113
timestamp 1688980957
transform 1 0 11500 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_119
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_123
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_135
timestamp 1688980957
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1688980957
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_166
timestamp 1688980957
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 6808 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 11040 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 6440 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 16376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 10212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 7176 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 4968 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 8464 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 12788 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 14260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 8280 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 14260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform -1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform -1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 2760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform -1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 9016 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform -1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 14996 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform -1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 14720 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 15548 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 15916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 15824 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 15824 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform -1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform -1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform -1 0 1932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 1688980957
transform -1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1688980957
transform -1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output49
timestamp 1688980957
transform -1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 1688980957
transform -1 0 2668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 1688980957
transform -1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 1688980957
transform -1 0 1932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output53
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output57
timestamp 1688980957
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sb_0__1__62
timestamp 1688980957
transform 1 0 15088 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
<< labels >>
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
flabel metal3 s 17200 8440 18000 8560 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 17200 9256 18000 9376 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 17200 1096 18000 1216 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 17200 1912 18000 2032 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 5 nsew signal input
flabel metal3 s 17200 2728 18000 2848 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 6 nsew signal input
flabel metal3 s 17200 3544 18000 3664 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 7 nsew signal input
flabel metal3 s 17200 4360 18000 4480 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 8 nsew signal input
flabel metal3 s 17200 5176 18000 5296 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 9 nsew signal input
flabel metal3 s 17200 5992 18000 6112 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 10 nsew signal input
flabel metal3 s 17200 6808 18000 6928 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 11 nsew signal input
flabel metal3 s 17200 7624 18000 7744 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 12 nsew signal input
flabel metal3 s 17200 10888 18000 11008 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 13 nsew signal tristate
flabel metal3 s 17200 11704 18000 11824 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 14 nsew signal tristate
flabel metal3 s 17200 12520 18000 12640 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 15 nsew signal tristate
flabel metal3 s 17200 13336 18000 13456 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 16 nsew signal tristate
flabel metal3 s 17200 14152 18000 14272 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 17 nsew signal tristate
flabel metal3 s 17200 14968 18000 15088 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 18 nsew signal tristate
flabel metal3 s 17200 15784 18000 15904 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 19 nsew signal tristate
flabel metal3 s 17200 16600 18000 16720 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 20 nsew signal tristate
flabel metal3 s 17200 17416 18000 17536 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 21 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 22 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 23 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 24 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 25 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 26 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 27 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 28 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 29 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 30 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 31 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 32 nsew signal tristate
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 33 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 34 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 35 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 36 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 37 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 38 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 39 nsew signal tristate
flabel metal2 s 2686 17200 2742 18000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 4250 17200 4306 18000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 41 nsew signal input
flabel metal2 s 5814 17200 5870 18000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 42 nsew signal input
flabel metal2 s 7378 17200 7434 18000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 43 nsew signal input
flabel metal2 s 8942 17200 8998 18000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 44 nsew signal input
flabel metal2 s 10506 17200 10562 18000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 45 nsew signal input
flabel metal2 s 12070 17200 12126 18000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 46 nsew signal input
flabel metal2 s 13634 17200 13690 18000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 47 nsew signal input
flabel metal2 s 15198 17200 15254 18000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 48 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chany_top_out[0]
port 49 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chany_top_out[1]
port 50 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chany_top_out[2]
port 51 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chany_top_out[3]
port 52 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chany_top_out[4]
port 53 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chany_top_out[5]
port 54 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_out[6]
port 55 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chany_top_out[7]
port 56 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chany_top_out[8]
port 57 nsew signal tristate
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 prog_clk
port 58 nsew signal input
flabel metal3 s 17200 10072 18000 10192 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 59 nsew signal input
flabel metal3 s 17200 280 18000 400 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 60 nsew signal input
flabel metal2 s 16762 17200 16818 18000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 61 nsew signal input
flabel metal2 s 1122 17200 1178 18000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 62 nsew signal input
flabel metal4 s 2910 2128 3230 15824 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 6843 2128 7163 15824 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 10776 2128 11096 15824 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 14709 2128 15029 15824 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 4876 2128 5196 15824 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 8809 2128 9129 15824 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 12742 2128 13062 15824 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 16675 2128 16995 15824 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
rlabel metal1 8970 15776 8970 15776 0 vdd
rlabel via1 9049 15232 9049 15232 0 vss
rlabel metal1 7176 3026 7176 3026 0 _000_
rlabel metal1 7912 4114 7912 4114 0 _001_
rlabel metal1 11270 11118 11270 11118 0 _002_
rlabel metal1 16054 12274 16054 12274 0 _003_
rlabel metal1 12512 6630 12512 6630 0 _004_
rlabel metal1 16698 6290 16698 6290 0 _005_
rlabel metal1 14306 6766 14306 6766 0 _006_
rlabel metal1 6302 10234 6302 10234 0 _007_
rlabel metal1 12926 10676 12926 10676 0 _008_
rlabel metal1 12972 10778 12972 10778 0 _009_
rlabel metal1 13616 13906 13616 13906 0 _010_
rlabel metal1 14950 12818 14950 12818 0 _011_
rlabel metal1 13248 13498 13248 13498 0 _012_
rlabel metal1 10304 14042 10304 14042 0 _013_
rlabel metal1 10810 14008 10810 14008 0 _014_
rlabel metal1 8924 13498 8924 13498 0 _015_
rlabel metal1 6900 11730 6900 11730 0 _016_
rlabel metal1 9614 11152 9614 11152 0 _017_
rlabel metal1 9660 10234 9660 10234 0 _018_
rlabel metal1 11868 8602 11868 8602 0 _019_
rlabel metal1 15226 6256 15226 6256 0 _020_
rlabel metal1 13386 5882 13386 5882 0 _021_
rlabel metal1 16836 3502 16836 3502 0 _022_
rlabel metal1 15364 5542 15364 5542 0 _023_
rlabel metal1 7038 6290 7038 6290 0 _024_
rlabel metal1 9062 8500 9062 8500 0 _025_
rlabel metal1 5980 7378 5980 7378 0 _026_
rlabel metal1 8050 9554 8050 9554 0 _027_
rlabel metal1 7222 8058 7222 8058 0 _028_
rlabel metal1 4508 10642 4508 10642 0 _029_
rlabel metal1 4232 7854 4232 7854 0 _030_
rlabel metal1 7590 6324 7590 6324 0 _031_
rlabel metal1 6026 8602 6026 8602 0 _032_
rlabel metal1 3128 7514 3128 7514 0 _033_
rlabel metal1 3496 7854 3496 7854 0 _034_
rlabel metal1 9752 8602 9752 8602 0 _035_
rlabel metal1 12466 5710 12466 5710 0 _036_
rlabel metal1 14398 3578 14398 3578 0 _037_
rlabel metal1 11316 6766 11316 6766 0 _038_
rlabel metal1 14766 3026 14766 3026 0 _039_
rlabel metal2 10350 5508 10350 5508 0 _040_
rlabel metal1 12604 5678 12604 5678 0 _041_
rlabel metal1 4416 6766 4416 6766 0 _042_
rlabel metal2 13754 5882 13754 5882 0 _043_
rlabel metal1 5014 5134 5014 5134 0 _044_
rlabel metal1 8418 5338 8418 5338 0 _045_
rlabel metal1 4278 4114 4278 4114 0 _046_
rlabel metal1 10810 2006 10810 2006 0 _047_
rlabel metal2 13754 4284 13754 4284 0 _048_
rlabel metal1 14444 4590 14444 4590 0 _049_
rlabel metal2 12558 2516 12558 2516 0 _050_
rlabel metal1 10902 3978 10902 3978 0 _051_
rlabel metal1 11592 2414 11592 2414 0 _052_
rlabel metal1 16008 4046 16008 4046 0 _053_
rlabel metal1 12512 2618 12512 2618 0 _054_
rlabel metal1 14950 4794 14950 4794 0 _055_
rlabel metal1 11270 4114 11270 4114 0 _056_
rlabel metal1 13984 4114 13984 4114 0 _057_
rlabel metal1 11960 2618 11960 2618 0 _058_
rlabel metal1 10396 3570 10396 3570 0 _059_
rlabel metal1 13340 4114 13340 4114 0 _060_
rlabel metal1 11776 3502 11776 3502 0 _061_
rlabel metal1 13156 3162 13156 3162 0 _062_
rlabel metal1 14674 4250 14674 4250 0 _063_
rlabel metal2 15962 4964 15962 4964 0 _064_
rlabel metal2 5566 4760 5566 4760 0 _065_
rlabel metal1 4692 4250 4692 4250 0 _066_
rlabel metal1 5474 6732 5474 6732 0 _067_
rlabel metal1 9062 5134 9062 5134 0 _068_
rlabel metal1 13938 5576 13938 5576 0 _069_
rlabel metal1 12880 5882 12880 5882 0 _070_
rlabel via1 5474 5253 5474 5253 0 _071_
rlabel metal1 5934 4046 5934 4046 0 _072_
rlabel metal2 4462 5508 4462 5508 0 _073_
rlabel metal1 7774 5202 7774 5202 0 _074_
rlabel metal1 15226 5338 15226 5338 0 _075_
rlabel metal1 3174 6426 3174 6426 0 _076_
rlabel metal1 11132 6970 11132 6970 0 _077_
rlabel metal1 11638 5066 11638 5066 0 _078_
rlabel metal1 12144 5882 12144 5882 0 _079_
rlabel metal1 15226 2924 15226 2924 0 _080_
rlabel metal2 14582 3791 14582 3791 0 _081_
rlabel metal1 9936 8466 9936 8466 0 _082_
rlabel metal1 11086 7752 11086 7752 0 _083_
rlabel metal1 11362 5202 11362 5202 0 _084_
rlabel metal1 11224 8398 11224 8398 0 _085_
rlabel metal2 15686 4692 15686 4692 0 _086_
rlabel metal1 15272 3706 15272 3706 0 _087_
rlabel metal1 9430 9452 9430 9452 0 _088_
rlabel metal1 5474 8840 5474 8840 0 _089_
rlabel metal1 3956 8058 3956 8058 0 _090_
rlabel metal1 4738 7786 4738 7786 0 _091_
rlabel metal1 3358 7446 3358 7446 0 _092_
rlabel metal1 8004 6154 8004 6154 0 _093_
rlabel metal2 4738 10948 4738 10948 0 _094_
rlabel metal1 5658 9622 5658 9622 0 _095_
rlabel metal1 4232 7990 4232 7990 0 _096_
rlabel metal2 4738 9588 4738 9588 0 _097_
rlabel metal1 4554 7378 4554 7378 0 _098_
rlabel metal1 8372 6290 8372 6290 0 _099_
rlabel metal1 5474 10642 5474 10642 0 _100_
rlabel metal1 8326 9452 8326 9452 0 _101_
rlabel metal1 8050 10132 8050 10132 0 _102_
rlabel metal1 7314 8432 7314 8432 0 _103_
rlabel metal1 6440 6290 6440 6290 0 _104_
rlabel metal1 7636 6426 7636 6426 0 _105_
rlabel metal1 8050 8500 8050 8500 0 _106_
rlabel metal1 8418 8908 8418 8908 0 _107_
rlabel metal1 8142 7922 8142 7922 0 _108_
rlabel metal1 5704 7514 5704 7514 0 _109_
rlabel metal1 7774 5882 7774 5882 0 _110_
rlabel metal2 16330 3859 16330 3859 0 _111_
rlabel metal1 15870 7276 15870 7276 0 _112_
rlabel metal1 15456 6426 15456 6426 0 _113_
rlabel metal1 15042 5780 15042 5780 0 _114_
rlabel metal1 14030 8840 14030 8840 0 _115_
rlabel metal1 16376 5338 16376 5338 0 _116_
rlabel metal1 16146 5032 16146 5032 0 _117_
rlabel metal1 14766 9690 14766 9690 0 _118_
rlabel metal1 13708 5746 13708 5746 0 _119_
rlabel metal2 13386 8908 13386 8908 0 _120_
rlabel metal1 10074 11016 10074 11016 0 _121_
rlabel metal1 10534 10676 10534 10676 0 _122_
rlabel metal2 6946 12036 6946 12036 0 _123_
rlabel metal2 9062 11560 9062 11560 0 _124_
rlabel metal1 10074 10540 10074 10540 0 _125_
rlabel metal1 7820 11186 7820 11186 0 _126_
rlabel metal1 11086 13192 11086 13192 0 _127_
rlabel metal1 9476 13906 9476 13906 0 _128_
rlabel metal1 10810 13906 10810 13906 0 _129_
rlabel metal1 11546 12954 11546 12954 0 _130_
rlabel metal1 9154 12818 9154 12818 0 _131_
rlabel metal1 10396 13362 10396 13362 0 _132_
rlabel metal1 14996 12954 14996 12954 0 _133_
rlabel metal1 12880 13362 12880 13362 0 _134_
rlabel metal1 14168 13906 14168 13906 0 _135_
rlabel metal1 15364 13362 15364 13362 0 _136_
rlabel metal2 12006 12036 12006 12036 0 _137_
rlabel metal1 13892 12818 13892 12818 0 _138_
rlabel metal1 13110 10540 13110 10540 0 _139_
rlabel metal1 13432 10642 13432 10642 0 _140_
rlabel metal1 6578 10540 6578 10540 0 _141_
rlabel metal2 12098 10914 12098 10914 0 _142_
rlabel metal1 14122 10234 14122 10234 0 _143_
rlabel metal1 7084 10778 7084 10778 0 _144_
rlabel metal1 15548 6086 15548 6086 0 _145_
rlabel metal1 14076 6630 14076 6630 0 _146_
rlabel metal2 12466 7820 12466 7820 0 _147_
rlabel metal1 13754 6834 13754 6834 0 _148_
rlabel metal1 13432 6834 13432 6834 0 _149_
rlabel metal2 12282 8772 12282 8772 0 _150_
rlabel metal1 16100 10710 16100 10710 0 _151_
rlabel metal1 11362 11016 11362 11016 0 _152_
rlabel metal1 15962 12886 15962 12886 0 _153_
rlabel metal1 10902 11764 10902 11764 0 _154_
rlabel metal1 9108 4182 9108 4182 0 _155_
rlabel metal2 7498 3298 7498 3298 0 _156_
rlabel metal1 8418 4216 8418 4216 0 _157_
rlabel metal1 7406 3570 7406 3570 0 _158_
rlabel metal2 874 1588 874 1588 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 15594 823 15594 823 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 16514 3060 16514 3060 0 ccff_head
rlabel metal1 16606 9146 16606 9146 0 ccff_tail
rlabel metal1 15318 2380 15318 2380 0 chanx_right_in[0]
rlabel metal1 15042 2448 15042 2448 0 chanx_right_in[1]
rlabel metal3 16522 2788 16522 2788 0 chanx_right_in[2]
rlabel metal2 14306 3315 14306 3315 0 chanx_right_in[3]
rlabel metal2 12374 3485 12374 3485 0 chanx_right_in[4]
rlabel metal2 13754 3689 13754 3689 0 chanx_right_in[5]
rlabel metal2 10396 2414 10396 2414 0 chanx_right_in[6]
rlabel metal1 15606 6294 15606 6294 0 chanx_right_in[7]
rlabel metal1 15686 5236 15686 5236 0 chanx_right_in[8]
rlabel via2 14582 11067 14582 11067 0 chanx_right_out[0]
rlabel metal3 16246 11764 16246 11764 0 chanx_right_out[1]
rlabel metal1 16514 13294 16514 13294 0 chanx_right_out[2]
rlabel metal2 16514 13651 16514 13651 0 chanx_right_out[3]
rlabel via2 16514 14331 16514 14331 0 chanx_right_out[4]
rlabel metal2 15594 15181 15594 15181 0 chanx_right_out[5]
rlabel metal1 16468 15674 16468 15674 0 chanx_right_out[6]
rlabel metal1 16468 15130 16468 15130 0 chanx_right_out[7]
rlabel metal2 2346 1027 2346 1027 0 chany_bottom_in[0]
rlabel metal2 3818 1027 3818 1027 0 chany_bottom_in[1]
rlabel metal2 5290 1027 5290 1027 0 chany_bottom_in[2]
rlabel metal2 6762 891 6762 891 0 chany_bottom_in[3]
rlabel metal2 8234 1588 8234 1588 0 chany_bottom_in[4]
rlabel metal2 9706 1588 9706 1588 0 chany_bottom_in[5]
rlabel metal2 11178 1554 11178 1554 0 chany_bottom_in[6]
rlabel metal2 12650 1027 12650 1027 0 chany_bottom_in[7]
rlabel metal2 14122 1588 14122 1588 0 chany_bottom_in[8]
rlabel metal3 820 10132 820 10132 0 chany_bottom_out[0]
rlabel metal3 1050 10948 1050 10948 0 chany_bottom_out[1]
rlabel metal3 820 11764 820 11764 0 chany_bottom_out[2]
rlabel metal3 820 12580 820 12580 0 chany_bottom_out[3]
rlabel metal3 1096 13396 1096 13396 0 chany_bottom_out[4]
rlabel metal3 820 14212 820 14212 0 chany_bottom_out[5]
rlabel metal3 935 15028 935 15028 0 chany_bottom_out[6]
rlabel metal3 820 15844 820 15844 0 chany_bottom_out[7]
rlabel metal3 1096 16660 1096 16660 0 chany_bottom_out[8]
rlabel metal2 2714 16943 2714 16943 0 chany_top_in[0]
rlabel metal2 4278 16943 4278 16943 0 chany_top_in[1]
rlabel metal2 5842 16943 5842 16943 0 chany_top_in[2]
rlabel metal2 7406 16943 7406 16943 0 chany_top_in[3]
rlabel metal2 8970 16943 8970 16943 0 chany_top_in[4]
rlabel metal1 10672 15470 10672 15470 0 chany_top_in[5]
rlabel metal1 12236 15470 12236 15470 0 chany_top_in[6]
rlabel metal1 13938 15504 13938 15504 0 chany_top_in[7]
rlabel metal2 15226 16398 15226 16398 0 chany_top_in[8]
rlabel metal3 820 1972 820 1972 0 chany_top_out[0]
rlabel metal3 820 2788 820 2788 0 chany_top_out[1]
rlabel metal3 820 3604 820 3604 0 chany_top_out[2]
rlabel metal3 820 4420 820 4420 0 chany_top_out[3]
rlabel metal3 751 5236 751 5236 0 chany_top_out[4]
rlabel metal3 820 6052 820 6052 0 chany_top_out[5]
rlabel metal3 1096 6868 1096 6868 0 chany_top_out[6]
rlabel metal3 820 7684 820 7684 0 chany_top_out[7]
rlabel metal3 820 8500 820 8500 0 chany_top_out[8]
rlabel metal1 7038 5712 7038 5712 0 clknet_0_prog_clk
rlabel metal1 9200 6290 9200 6290 0 clknet_2_0__leaf_prog_clk
rlabel metal1 6440 9554 6440 9554 0 clknet_2_1__leaf_prog_clk
rlabel metal1 12604 8942 12604 8942 0 clknet_2_2__leaf_prog_clk
rlabel metal1 9660 12818 9660 12818 0 clknet_2_3__leaf_prog_clk
rlabel metal1 8556 4454 8556 4454 0 mem_bottom_track_1.DFF_0_.D
rlabel metal2 9614 7735 9614 7735 0 mem_bottom_track_1.DFF_0_.Q
rlabel metal1 10304 6086 10304 6086 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal1 10074 7174 10074 7174 0 mem_bottom_track_1.DFF_2_.Q
rlabel metal1 5520 9350 5520 9350 0 mem_bottom_track_17.DFF_0_.D
rlabel metal1 13294 9690 13294 9690 0 mem_bottom_track_17.DFF_0_.Q
rlabel metal1 16514 5644 16514 5644 0 mem_bottom_track_17.DFF_1_.Q
rlabel metal1 4278 10540 4278 10540 0 mem_bottom_track_9.DFF_0_.Q
rlabel metal1 3312 10030 3312 10030 0 mem_bottom_track_9.DFF_1_.Q
rlabel metal1 15824 11730 15824 11730 0 mem_right_track_10.DFF_0_.D
rlabel metal1 7820 10642 7820 10642 0 mem_right_track_10.DFF_0_.Q
rlabel metal2 12282 9945 12282 9945 0 mem_right_track_10.DFF_1_.Q
rlabel metal1 13938 7412 13938 7412 0 mem_right_track_12.DFF_0_.Q
rlabel metal1 13938 6834 13938 6834 0 mem_right_track_12.DFF_1_.Q
rlabel metal2 6394 4420 6394 4420 0 mem_right_track_14.DFF_0_.Q
rlabel metal1 6900 9350 6900 9350 0 mem_right_track_2.DFF_0_.D
rlabel metal1 9108 10642 9108 10642 0 mem_right_track_2.DFF_0_.Q
rlabel metal1 10212 11730 10212 11730 0 mem_right_track_2.DFF_1_.Q
rlabel metal1 9384 13294 9384 13294 0 mem_right_track_4.DFF_0_.Q
rlabel metal2 11546 14110 11546 14110 0 mem_right_track_4.DFF_1_.Q
rlabel metal1 12788 12614 12788 12614 0 mem_right_track_6.DFF_0_.Q
rlabel metal1 14214 13260 14214 13260 0 mem_right_track_6.DFF_1_.Q
rlabel metal1 14628 12750 14628 12750 0 mem_right_track_8.DFF_0_.Q
rlabel metal2 14122 6494 14122 6494 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 12742 4148 12742 4148 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 13570 4794 13570 4794 0 mem_top_track_0.DFF_2_.Q
rlabel metal1 6440 6766 6440 6766 0 mem_top_track_16.DFF_0_.D
rlabel metal1 7222 6766 7222 6766 0 mem_top_track_16.DFF_0_.Q
rlabel metal1 6026 8500 6026 8500 0 mem_top_track_16.DFF_1_.Q
rlabel metal1 8188 5746 8188 5746 0 mem_top_track_8.DFF_0_.Q
rlabel metal1 4600 5134 4600 5134 0 mem_top_track_8.DFF_1_.Q
rlabel metal1 6624 11118 6624 11118 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 9752 14246 9752 14246 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 15226 2618 15226 2618 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 13800 4046 13800 4046 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 16192 5678 16192 5678 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 14766 2958 14766 2958 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 10212 8602 10212 8602 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14950 4182 14950 4182 0 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 15548 5678 15548 5678 0 mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 11178 7667 11178 7667 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10672 6426 10672 6426 0 mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 8326 7752 8326 7752 0 mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 13202 12818 13202 12818 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 12282 14246 12282 14246 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 13110 6154 13110 6154 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 14674 5678 14674 5678 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 15548 6698 15548 6698 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal2 14490 9350 14490 9350 0 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 15318 7140 15318 7140 0 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 15686 9010 15686 9010 0 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 15548 7446 15548 7446 0 mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 8142 12512 8142 12512 0 mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 5773 12886 5773 12886 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 5658 11254 5658 11254 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal2 8510 5967 8510 5967 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal2 7958 4930 7958 4930 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 9614 2448 9614 2448 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 3128 3162 3128 3162 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal2 4830 10880 4830 10880 0 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 7866 6800 7866 6800 0 mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4370 7514 4370 7514 0 mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 5382 9486 5382 9486 0 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 4968 8330 4968 8330 0 mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 2760 12818 2760 12818 0 mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 6394 8398 6394 8398 0 mux_right_track_10.INVTX1_1_.out
rlabel metal2 13938 3587 13938 3587 0 mux_right_track_10.INVTX1_2_.out
rlabel metal1 7636 10710 7636 10710 0 mux_right_track_10.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14582 10438 14582 10438 0 mux_right_track_10.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 13754 11186 13754 11186 0 mux_right_track_10.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10810 5304 10810 5304 0 mux_right_track_12.INVTX1_1_.out
rlabel metal2 13478 4964 13478 4964 0 mux_right_track_12.INVTX1_2_.out
rlabel metal1 12788 8534 12788 8534 0 mux_right_track_12.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13156 7514 13156 7514 0 mux_right_track_12.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 14214 14994 14214 14994 0 mux_right_track_12.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7728 3502 7728 3502 0 mux_right_track_14.INVTX1_0_.out
rlabel metal1 7912 3162 7912 3162 0 mux_right_track_14.INVTX1_1_.out
rlabel metal1 8280 3638 8280 3638 0 mux_right_track_14.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9890 4046 9890 4046 0 mux_right_track_14.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 7590 13605 7590 13605 0 mux_right_track_2.INVTX1_1_.out
rlabel metal1 16376 9690 16376 9690 0 mux_right_track_2.INVTX1_2_.out
rlabel metal1 7912 12070 7912 12070 0 mux_right_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 10304 10438 10304 10438 0 mux_right_track_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 13846 8670 13846 8670 0 mux_right_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11362 13838 11362 13838 0 mux_right_track_4.INVTX1_1_.out
rlabel metal1 8694 12750 8694 12750 0 mux_right_track_4.INVTX1_2_.out
rlabel metal2 10718 13600 10718 13600 0 mux_right_track_4.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 9706 13328 9706 13328 0 mux_right_track_4.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 11960 13430 11960 13430 0 mux_right_track_4.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 14674 13940 14674 13940 0 mux_right_track_6.INVTX1_1_.out
rlabel metal1 9936 6834 9936 6834 0 mux_right_track_6.INVTX1_2_.out
rlabel metal2 14306 13192 14306 13192 0 mux_right_track_6.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 12972 13158 12972 13158 0 mux_right_track_6.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 15686 13940 15686 13940 0 mux_right_track_6.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11224 4046 11224 4046 0 mux_right_track_8.INVTX1_1_.out
rlabel metal1 15456 12750 15456 12750 0 mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 15916 12750 15916 12750 0 mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 14766 14790 14766 14790 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 16330 4114 16330 4114 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14490 4998 14490 4998 0 mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 10718 3808 10718 3808 0 mux_top_track_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 13340 3910 13340 3910 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11776 3162 11776 3162 0 mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 12834 3162 12834 3162 0 mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 8004 7514 8004 7514 0 mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7222 8330 7222 8330 0 mux_top_track_16.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 7682 8160 7682 8160 0 mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7866 9486 7866 9486 0 mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 8510 8976 8510 8976 0 mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3128 14790 3128 14790 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 4094 6188 4094 6188 0 mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel via2 14858 6851 14858 6851 0 mux_top_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 7268 5202 7268 5202 0 mux_top_track_8.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 4692 6426 4692 6426 0 mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5934 4658 5934 4658 0 mux_top_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 2162 5780 2162 5780 0 mux_top_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 2484 2618 2484 2618 0 net1
rlabel metal1 10718 1904 10718 1904 0 net10
rlabel via1 9885 12818 9885 12818 0 net100
rlabel metal1 5704 9146 5704 9146 0 net101
rlabel metal1 9885 7446 9885 7446 0 net102
rlabel metal2 7590 11526 7590 11526 0 net103
rlabel metal1 13570 4556 13570 4556 0 net104
rlabel metal2 9890 5814 9890 5814 0 net105
rlabel viali 13406 10028 13406 10028 0 net106
rlabel metal1 15962 3502 15962 3502 0 net11
rlabel metal1 15502 4182 15502 4182 0 net12
rlabel metal2 2622 2754 2622 2754 0 net13
rlabel metal1 4002 3536 4002 3536 0 net14
rlabel metal1 5520 4114 5520 4114 0 net15
rlabel metal1 7314 2618 7314 2618 0 net16
rlabel metal1 8924 2618 8924 2618 0 net17
rlabel metal1 9062 6188 9062 6188 0 net18
rlabel metal2 11914 2397 11914 2397 0 net19
rlabel metal1 14030 2550 14030 2550 0 net2
rlabel metal1 13294 2618 13294 2618 0 net20
rlabel metal1 14122 2618 14122 2618 0 net21
rlabel metal1 2898 15334 2898 15334 0 net22
rlabel metal1 4554 12886 4554 12886 0 net23
rlabel metal2 6210 13396 6210 13396 0 net24
rlabel metal1 7590 14994 7590 14994 0 net25
rlabel metal1 9292 14382 9292 14382 0 net26
rlabel metal1 5474 14994 5474 14994 0 net27
rlabel metal1 12006 14994 12006 14994 0 net28
rlabel metal1 13570 14382 13570 14382 0 net29
rlabel metal1 16790 3162 16790 3162 0 net3
rlabel metal1 14858 14416 14858 14416 0 net30
rlabel metal1 16284 8602 16284 8602 0 net31
rlabel metal1 10948 2414 10948 2414 0 net32
rlabel metal1 14812 14994 14812 14994 0 net33
rlabel metal1 2852 14994 2852 14994 0 net34
rlabel metal2 16146 8602 16146 8602 0 net35
rlabel metal1 11270 2550 11270 2550 0 net36
rlabel metal1 15916 13906 15916 13906 0 net37
rlabel metal1 15778 13294 15778 13294 0 net38
rlabel metal1 15962 13974 15962 13974 0 net39
rlabel metal1 8418 3060 8418 3060 0 net4
rlabel metal1 16146 14484 16146 14484 0 net40
rlabel metal2 15778 15266 15778 15266 0 net41
rlabel metal1 15226 14926 15226 14926 0 net42
rlabel metal1 16146 14926 16146 14926 0 net43
rlabel metal2 1794 9622 1794 9622 0 net44
rlabel metal1 2024 11118 2024 11118 0 net45
rlabel metal1 1886 12138 1886 12138 0 net46
rlabel metal1 1794 12784 1794 12784 0 net47
rlabel metal1 1932 12954 1932 12954 0 net48
rlabel metal1 4347 14314 4347 14314 0 net49
rlabel metal1 14812 2414 14812 2414 0 net5
rlabel metal1 4416 15130 4416 15130 0 net50
rlabel metal1 1978 15504 1978 15504 0 net51
rlabel metal1 2024 14994 2024 14994 0 net52
rlabel metal1 10074 2414 10074 2414 0 net53
rlabel metal1 1886 3094 1886 3094 0 net54
rlabel metal2 3818 3944 3818 3944 0 net55
rlabel metal2 5290 4386 5290 4386 0 net56
rlabel metal1 1932 5610 1932 5610 0 net57
rlabel metal1 6302 5814 6302 5814 0 net58
rlabel metal2 1794 7174 1794 7174 0 net59
rlabel metal1 11408 2414 11408 2414 0 net6
rlabel metal1 1886 7786 1886 7786 0 net60
rlabel metal1 1794 9010 1794 9010 0 net61
rlabel metal1 15180 14994 15180 14994 0 net62
rlabel metal1 12282 3094 12282 3094 0 net63
rlabel metal1 4462 4658 4462 4658 0 net64
rlabel metal1 11270 6324 11270 6324 0 net65
rlabel metal1 4140 8466 4140 8466 0 net66
rlabel metal1 8280 10030 8280 10030 0 net67
rlabel metal1 16146 4658 16146 4658 0 net68
rlabel metal1 10028 10642 10028 10642 0 net69
rlabel metal1 8142 2958 8142 2958 0 net7
rlabel metal1 9154 13838 9154 13838 0 net70
rlabel metal2 12742 13600 12742 13600 0 net71
rlabel metal2 13294 11152 13294 11152 0 net72
rlabel metal2 14122 7072 14122 7072 0 net73
rlabel metal2 15778 12274 15778 12274 0 net74
rlabel metal1 9200 4046 9200 4046 0 net75
rlabel metal2 10350 12002 10350 12002 0 net76
rlabel metal2 8970 10438 8970 10438 0 net77
rlabel metal1 9460 9622 9460 9622 0 net78
rlabel metal2 10350 7378 10350 7378 0 net79
rlabel metal1 11914 2550 11914 2550 0 net8
rlabel metal3 13662 9588 13662 9588 0 net80
rlabel metal2 9614 4114 9614 4114 0 net81
rlabel metal1 7114 4522 7114 4522 0 net82
rlabel via1 5938 6290 5938 6290 0 net83
rlabel metal1 12001 12886 12001 12886 0 net84
rlabel metal1 13580 5202 13580 5202 0 net85
rlabel metal1 15425 12138 15425 12138 0 net86
rlabel metal1 15690 11050 15690 11050 0 net87
rlabel metal1 14393 11798 14393 11798 0 net88
rlabel via1 7502 4114 7502 4114 0 net89
rlabel metal1 15318 3536 15318 3536 0 net9
rlabel metal2 15226 9078 15226 9078 0 net90
rlabel metal1 6578 6970 6578 6970 0 net91
rlabel metal2 4278 5474 4278 5474 0 net92
rlabel metal1 4012 5202 4012 5202 0 net93
rlabel metal1 4319 9622 4319 9622 0 net94
rlabel metal1 12803 7786 12803 7786 0 net95
rlabel metal1 12921 12138 12921 12138 0 net96
rlabel metal2 7222 9350 7222 9350 0 net97
rlabel metal2 12098 4386 12098 4386 0 net98
rlabel metal1 13197 8942 13197 8942 0 net99
rlabel metal3 1671 9316 1671 9316 0 prog_clk
rlabel metal1 16054 8432 16054 8432 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 13938 1377 13938 1377 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 14950 15504 14950 15504 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 2024 15062 2024 15062 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
