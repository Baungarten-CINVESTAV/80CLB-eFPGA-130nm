* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt sb_1__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
+ prog_clk right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
+ vdd vss
XFILLER_0_27_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_294_ _044_ vss vss vdd vdd _061_ sky130_fd_sc_hd__clkbuf_1
X_363_ clknet_2_0__leaf_prog_clk net75 vss vss vdd vdd mem_left_track_17.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_501_ net73 _139_ vss vss vdd vdd mux_left_track_9.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_39 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_432_ mux_left_track_17.mux_l2_in_1_.TGATE_0_.out _070_ vss vss vdd vdd mux_left_track_17.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_346_ net30 vss vss vdd vdd mux_left_track_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_415_ mux_left_track_9.INVTX1_3_.out _053_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_24_72 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_277_ mem_left_track_17.DFF_1_.Q vss vss vdd vdd _076_ sky130_fd_sc_hd__inv_2
X_200_ _012_ vss vss vdd vdd _119_ sky130_fd_sc_hd__clkbuf_1
X_329_ mux_top_track_16.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net62 sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_452__68 vss vss vdd vdd net68 _452__68/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_117 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_16_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_9 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput53 net53 vss vss vdd vdd chanx_right_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 vss vss vdd vdd chanx_left_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_123 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_293_ mem_right_track_16.DFF_1_.Q vss vss vdd vdd _044_ sky130_fd_sc_hd__clkbuf_1
X_500_ mux_left_track_9.mux_l2_in_1_.TGATE_0_.out _138_ vss vss vdd vdd mux_left_track_9.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_431_ mux_left_track_17.INVTX1_0_.out _069_ vss vss vdd vdd mux_right_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_362_ clknet_2_2__leaf_prog_clk net89 vss vss vdd vdd mem_left_track_17.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_120 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_414_ mux_top_track_0.mux_l1_in_1_.TGATE_0_.out _052_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_345_ net20 vss vss vdd vdd mux_left_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_276_ _038_ vss vss vdd vdd _070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_61 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_259_ _032_ vss vss vdd vdd _082_ sky130_fd_sc_hd__clkbuf_1
X_328_ net10 vss vss vdd vdd mux_top_track_14.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_21_52 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold20 mem_right_track_16.DFF_0_.Q vss vss vdd vdd net93 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_62 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_21_132 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_6_18 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput54 net54 vss vss vdd vdd chany_top_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput43 net43 vss vss vdd vdd chanx_left_out[7] sky130_fd_sc_hd__clkbuf_4
XTAP_124 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ mem_right_track_16.DFF_1_.Q vss vss vdd vdd _066_ sky130_fd_sc_hd__inv_2
X_430_ mux_left_track_17.INVTX1_2_.out _068_ vss vss vdd vdd mux_right_track_16.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_361_ clknet_2_2__leaf_prog_clk net99 vss vss vdd vdd net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_413_ mux_top_track_0.mux_l2_in_1_.TGATE_0_.out _051_ vss vss vdd vdd mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_344_ net23 vss vss vdd vdd mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_275_ net35 vss vss vdd vdd _038_ sky130_fd_sc_hd__clkbuf_1
X_258_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _032_ sky130_fd_sc_hd__clkbuf_1
X_327_ mux_top_track_14.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net61 sky130_fd_sc_hd__inv_2
XFILLER_0_19_116 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_189_ _009_ vss vss vdd vdd _126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_97 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_42 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_74 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold21 mem_top_track_0.DFF_1_.Q vss vss vdd vdd net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 mem_top_track_2.DFF_1_.Q vss vss vdd vdd net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput55 net55 vss vss vdd vdd chany_top_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 vss vss vdd vdd chanx_left_out[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_125 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_85 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_114 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ _043_ vss vss vdd vdd _060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_141 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_360_ clknet_2_2__leaf_prog_clk net78 vss vss vdd vdd mem_right_track_16.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_489_ net72 _127_ vss vss vdd vdd mux_left_track_1.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_412_ net63 _050_ vss vss vdd vdd mux_top_track_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_343_ net26 vss vss vdd vdd mux_left_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_274_ _037_ vss vss vdd vdd _073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_257_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _085_ sky130_fd_sc_hd__inv_2
X_326_ mux_top_track_8.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net58 sky130_fd_sc_hd__inv_2
X_188_ mem_left_track_1.DFF_2_.Q vss vss vdd vdd _009_ sky130_fd_sc_hd__clkbuf_1
X_309_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _055_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_109 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_21_76 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold11 mem_top_track_8.DFF_0_.Q vss vss vdd vdd net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 mem_left_track_1.DFF_0_.Q vss vss vdd vdd net95 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput56 net56 vss vss vdd vdd chany_top_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput45 net45 vss vss vdd vdd chanx_right_out[0] sky130_fd_sc_hd__clkbuf_4
XTAP_126 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412__63 vss vss vdd vdd net63 _412__63/LO sky130_fd_sc_hd__conb_1
X_290_ mem_left_track_1.DFF_0_.D vss vss vdd vdd _043_ sky130_fd_sc_hd__clkbuf_1
X_488_ mux_left_track_1.mux_l2_in_1_.TGATE_0_.out _126_ vss vss vdd vdd mux_left_track_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_1_101 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_411_ net15 vss vss vdd vdd net56 sky130_fd_sc_hd__clkbuf_1
X_273_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _037_ sky130_fd_sc_hd__clkbuf_1
X_342_ net11 vss vss vdd vdd mux_left_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_4_53 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_4_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_325_ net19 vss vss vdd vdd mux_top_track_2.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_256_ mem_top_track_2.DFF_1_.Q vss vss vdd vdd _083_ sky130_fd_sc_hd__inv_2
X_187_ _008_ vss vss vdd vdd _130_ sky130_fd_sc_hd__clkbuf_1
X_308_ _049_ vss vss vdd vdd _050_ sky130_fd_sc_hd__clkbuf_1
X_239_ mem_right_track_0.DFF_0_.D vss vss vdd vdd _026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_87 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_43 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold12 mem_top_track_16.DFF_0_.Q vss vss vdd vdd net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 mem_left_track_9.DFF_0_.Q vss vss vdd vdd net96 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_3__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_44 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput57 net57 vss vss vdd vdd chany_top_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput46 net46 vss vss vdd vdd chanx_right_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_0_7_140 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_127 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_34 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_487_ mux_left_track_1.INVTX1_0_.out _125_ vss vss vdd vdd mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_410_ net16 vss vss vdd vdd net57 sky130_fd_sc_hd__clkbuf_1
X_272_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _078_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_341_ net15 vss vss vdd vdd mux_left_track_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_0_24_44 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_324_ net34 vss vss vdd vdd mux_top_track_2.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_255_ _031_ vss vss vdd vdd _086_ sky130_fd_sc_hd__clkbuf_1
X_186_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_130 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_307_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _049_ sky130_fd_sc_hd__clkbuf_1
X_169_ _002_ vss vss vdd vdd _142_ sky130_fd_sc_hd__clkbuf_1
X_238_ _025_ vss vss vdd vdd _096_ sky130_fd_sc_hd__clkbuf_1
Xhold24 mem_right_track_0.DFF_1_.Q vss vss vdd vdd net97 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold13 mem_left_track_1.DFF_2_.Q vss vss vdd vdd net86 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput58 net58 vss vss vdd vdd chany_top_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput47 net47 vss vss vdd vdd chanx_right_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput36 net36 vss vss vdd vdd chanx_left_out[0] sky130_fd_sc_hd__clkbuf_4
XTAP_128 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_7_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_68 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_486_ mux_left_track_1.INVTX1_2_.out _124_ vss vss vdd vdd mux_right_track_8.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_271_ _036_ vss vss vdd vdd _072_ sky130_fd_sc_hd__clkbuf_1
X_340_ mux_left_track_1.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net36 sky130_fd_sc_hd__inv_2
X_469_ mux_left_track_9.INVTX1_1_.out _107_ vss vss vdd vdd mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_323_ mux_top_track_2.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net55 sky130_fd_sc_hd__inv_2
X_254_ mem_top_track_14.DFF_0_.D vss vss vdd vdd _031_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_185_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _136_ sky130_fd_sc_hd__inv_2
X_306_ _048_ vss vss vdd vdd _051_ sky130_fd_sc_hd__clkbuf_1
X_168_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _002_ sky130_fd_sc_hd__clkbuf_1
X_237_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _025_ sky130_fd_sc_hd__clkbuf_1
Xhold14 mem_top_track_2.DFF_0_.Q vss vss vdd vdd net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 mem_left_track_9.DFF_1_.Q vss vss vdd vdd net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_12 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput59 net59 vss vss vdd vdd chany_top_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput48 net48 vss vss vdd vdd chanx_right_out[3] sky130_fd_sc_hd__clkbuf_4
Xoutput37 net37 vss vss vdd vdd chanx_left_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_120 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_129 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_22 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_47 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_126 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_485_ mux_right_track_8.INVTX1_4_.out _123_ vss vss vdd vdd mux_right_track_8.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xclkbuf_2_0__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_2_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_270_ mem_left_track_17.DFF_1_.Q vss vss vdd vdd _036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_468_ mux_right_track_0.INVTX1_3_.out _106_ vss vss vdd vdd mux_right_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_399_ net13 vss vss vdd vdd net39 sky130_fd_sc_hd__clkbuf_1
X_322_ net17 vss vss vdd vdd mux_left_track_17.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_253_ _030_ vss vss vdd vdd _087_ sky130_fd_sc_hd__clkbuf_1
X_184_ _007_ vss vss vdd vdd _128_ sky130_fd_sc_hd__clkbuf_1
X_305_ mem_top_track_0.DFF_2_.Q vss vss vdd vdd _048_ sky130_fd_sc_hd__clkbuf_1
X_167_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _148_ sky130_fd_sc_hd__inv_2
X_236_ _024_ vss vss vdd vdd _097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_135 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_1_79 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_35 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_1_24 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xhold26 mem_left_track_17.DFF_1_.Q vss vss vdd vdd net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 mem_right_track_8.DFF_1_.Q vss vss vdd vdd net88 sky130_fd_sc_hd__dlygate4sd3_1
X_219_ mem_right_track_0.DFF_1_.Q vss vss vdd vdd _019_ sky130_fd_sc_hd__clkbuf_1
Xoutput49 net49 vss vss vdd vdd chanx_right_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput38 net38 vss vss vdd vdd chanx_left_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_132 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_27_46 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_119 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_7_34 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_484_ mux_right_track_8.mux_l1_in_0_.TGATE_0_.out _122_ vss vss vdd vdd mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_467_ mux_right_track_0.INVTX1_5_.out _105_ vss vss vdd vdd mux_right_track_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_398_ net15 vss vss vdd vdd net41 sky130_fd_sc_hd__clkbuf_1
X_252_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _030_ sky130_fd_sc_hd__clkbuf_1
X_321_ net21 vss vss vdd vdd mux_left_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_183_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_133 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_304_ _047_ vss vss vdd vdd _054_ sky130_fd_sc_hd__clkbuf_1
X_235_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _024_ sky130_fd_sc_hd__clkbuf_1
X_166_ _001_ vss vss vdd vdd _140_ sky130_fd_sc_hd__clkbuf_1
Xhold27 mem_right_track_0.DFF_0_.Q vss vss vdd vdd net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 mem_left_track_17.DFF_0_.Q vss vss vdd vdd net89 sky130_fd_sc_hd__dlygate4sd3_1
X_218_ _018_ vss vss vdd vdd _107_ sky130_fd_sc_hd__clkbuf_1
X_433__65 vss vss vdd vdd net65 _433__65/LO sky130_fd_sc_hd__conb_1
XFILLER_0_12_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput39 net39 vss vss vdd vdd chanx_left_out[3] sky130_fd_sc_hd__clkbuf_4
XTAP_109 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_46 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_7_79 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_483_ mux_right_track_8.mux_l1_in_2_.TGATE_0_.out _121_ vss vss vdd vdd mux_right_track_8.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_24_15 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_466_ mux_right_track_0.mux_l1_in_1_.TGATE_0_.out _104_ vss vss vdd vdd mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_397_ net16 vss vss vdd vdd net42 sky130_fd_sc_hd__buf_1
XFILLER_0_5_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_320_ net24 vss vss vdd vdd mux_left_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_251_ mem_top_track_8.DFF_0_.Q vss vss vdd vdd _089_ sky130_fd_sc_hd__inv_2
X_182_ _006_ vss vss vdd vdd _131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_449_ mux_right_track_16.INVTX1_4_.out _087_ vss vss vdd vdd mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_25_91 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_303_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_38 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_165_ mem_left_track_9.DFF_1_.Q vss vss vdd vdd _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_48 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_234_ mem_top_track_16.DFF_0_.Q vss vss vdd vdd _101_ sky130_fd_sc_hd__inv_2
Xhold17 mem_top_track_16.DFF_1_.Q vss vss vdd vdd net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 mem_left_track_1.DFF_1_.Q vss vss vdd vdd net101 sky130_fd_sc_hd__dlygate4sd3_1
X_217_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_118 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_11_140 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_482_ mux_right_track_8.mux_l2_in_0_.TGATE_0_.out _120_ vss vss vdd vdd mux_right_track_8.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_24_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_465_ net70 _103_ vss vss vdd vdd mux_right_track_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_396_ net17 vss vss vdd vdd net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_4_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_250_ mem_top_track_14.DFF_0_.D vss vss vdd vdd _088_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_181_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _006_ sky130_fd_sc_hd__clkbuf_1
X_448_ net67 _086_ vss vss vdd vdd mux_top_track_8.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_379_ clknet_2_0__leaf_prog_clk net101 vss vss vdd vdd mem_left_track_1.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_302_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _058_ sky130_fd_sc_hd__inv_2
X_164_ _000_ vss vss vdd vdd _143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_17 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_233_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _100_ sky130_fd_sc_hd__inv_2
Xhold29 mem_top_track_0.DFF_0_.Q vss vss vdd vdd net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 mem_right_track_16.DFF_1_.Q vss vss vdd vdd net91 sky130_fd_sc_hd__dlygate4sd3_1
X_216_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _113_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_18_8 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_8 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_481_ mux_left_track_1.INVTX1_1_.out _119_ vss vss vdd vdd mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_0_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_464_ mux_right_track_0.mux_l2_in_1_.TGATE_0_.out _102_ vss vss vdd vdd mux_right_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_180_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _137_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_125 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_447_ mux_top_track_2.INVTX1_0_.out _085_ vss vss vdd vdd mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_378_ clknet_2_2__leaf_prog_clk net74 vss vss vdd vdd mem_right_track_8.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_301_ _046_ vss vss vdd vdd _052_ sky130_fd_sc_hd__clkbuf_1
X_163_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _000_ sky130_fd_sc_hd__clkbuf_1
X_232_ mem_right_track_0.DFF_0_.D vss vss vdd vdd _098_ sky130_fd_sc_hd__inv_2
Xhold19 mem_right_track_8.DFF_0_.Q vss vss vdd vdd net92 sky130_fd_sc_hd__dlygate4sd3_1
X_215_ mem_right_track_0.DFF_1_.Q vss vss vdd vdd _110_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_71 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_480_ mux_right_track_8.INVTX1_3_.out _118_ vss vss vdd vdd mux_right_track_8.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_24_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_463_ mux_left_track_1.INVTX1_3_.out _101_ vss vss vdd vdd mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_446_ mux_top_track_2.INVTX1_2_.out _084_ vss vss vdd vdd mux_top_track_2.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_377_ clknet_2_0__leaf_prog_clk net92 vss vss vdd vdd mem_right_track_8.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_24_118 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_300_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _046_ sky130_fd_sc_hd__clkbuf_1
X_162_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _149_ sky130_fd_sc_hd__inv_2
X_231_ _023_ vss vss vdd vdd _103_ sky130_fd_sc_hd__clkbuf_1
X_429_ mux_right_track_16.mux_l1_in_0_.TGATE_0_.out _067_ vss vss vdd vdd mux_right_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
Xinput1 ccff_head vss vss vdd vdd net1 sky130_fd_sc_hd__buf_1
XTAP_90 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ mem_right_track_0.DFF_2_.Q vss vss vdd vdd _108_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_27_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_462_ mux_top_track_16.mux_l1_in_0_.TGATE_0_.out _100_ vss vss vdd vdd mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_4_18 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_96 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_445_ mux_top_track_2.mux_l1_in_0_.TGATE_0_.out _083_ vss vss vdd vdd mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_376_ clknet_2_2__leaf_prog_clk net88 vss vss vdd vdd mem_right_track_16.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
X_230_ mem_right_track_0.DFF_1_.Q vss vss vdd vdd _023_ sky130_fd_sc_hd__clkbuf_1
X_161_ mem_left_track_9.DFF_1_.Q vss vss vdd vdd _146_ sky130_fd_sc_hd__inv_2
X_428_ mux_right_track_16.INVTX1_4_.out _066_ vss vss vdd vdd mux_right_track_16.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_359_ clknet_2_3__leaf_prog_clk net93 vss vss vdd vdd mem_right_track_16.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_91 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 chanx_left_in[0] vss vss vdd vdd net2 sky130_fd_sc_hd__buf_1
XTAP_80 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _017_ vss vss vdd vdd _115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_122 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_461_ mux_top_track_16.INVTX1_3_.out _099_ vss vss vdd vdd mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_444_ mux_left_track_17.INVTX1_3_.out _082_ vss vss vdd vdd mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_375_ clknet_2_3__leaf_prog_clk net81 vss vss vdd vdd mem_right_track_0.DFF_0_.Q
+ sky130_fd_sc_hd__dfxtp_2
X_427_ mux_right_track_16.mux_l2_in_0_.TGATE_0_.out _065_ vss vss vdd vdd mux_right_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_358_ clknet_2_2__leaf_prog_clk net91 vss vss vdd vdd mem_left_track_1.DFF_0_.D sky130_fd_sc_hd__dfxtp_1
X_289_ _042_ vss vss vdd vdd _063_ sky130_fd_sc_hd__clkbuf_1
XTAP_92 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[1] vss vss vdd vdd net3 sky130_fd_sc_hd__buf_1
XTAP_70 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ mem_right_track_8.DFF_1_.Q vss vss vdd vdd _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_134 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_460_ mux_top_track_16.mux_l2_in_0_.TGATE_0_.out _098_ vss vss vdd vdd mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_443_ net66 _081_ vss vss vdd vdd mux_top_track_2.mux_l1_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_374_ clknet_2_1__leaf_prog_clk net100 vss vss vdd vdd mem_right_track_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_74 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_357_ clknet_2_3__leaf_prog_clk net1 vss vss vdd vdd mem_top_track_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
X_288_ mem_right_track_16.DFF_0_.Q vss vss vdd vdd _042_ sky130_fd_sc_hd__clkbuf_1
X_426_ mux_left_track_17.INVTX1_1_.out _064_ vss vss vdd vdd mux_right_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_93 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 chanx_left_in[2] vss vss vdd vdd net4 sky130_fd_sc_hd__buf_1
XTAP_82 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _016_ vss vss vdd vdd _117_ sky130_fd_sc_hd__clkbuf_1
X_409_ net7 vss vss vdd vdd net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_17_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_14_7 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_0_135 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_8_41 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_14_88 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_14_22 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_448__67 vss vss vdd vdd net67 _448__67/LO sky130_fd_sc_hd__conb_1
X_442_ mux_top_track_2.mux_l1_in_1_.TGATE_0_.out _080_ vss vss vdd vdd mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_511_ mux_left_track_9.INVTX1_0_.out _149_ vss vss vdd vdd mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_373_ clknet_2_1__leaf_prog_clk net97 vss vss vdd vdd mem_right_track_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_87 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_356_ clknet_2_1__leaf_prog_clk net102 vss vss vdd vdd mem_top_track_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_425_ mux_right_track_16.INVTX1_3_.out _063_ vss vss vdd vdd mux_right_track_16.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_287_ mem_right_track_16.DFF_0_.Q vss vss vdd vdd _068_ sky130_fd_sc_hd__inv_2
Xinput5 chanx_left_in[3] vss vss vdd vdd net5 sky130_fd_sc_hd__clkbuf_1
XTAP_94 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ net6 vss vss vdd vdd net60 sky130_fd_sc_hd__clkbuf_1
X_210_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_77 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_339_ net7 vss vss vdd vdd mux_right_track_8.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_0_6_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xinput30 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_ vss vss vdd vdd
+ net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_100 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_78 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_27_109 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_372_ clknet_2_3__leaf_prog_clk net82 vss vss vdd vdd mem_top_track_16.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_510_ mux_left_track_9.INVTX1_2_.out _148_ vss vss vdd vdd mux_left_track_9.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_441_ mux_left_track_17.INVTX1_0_.out _079_ vss vss vdd vdd mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_25_66 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_355_ clknet_2_1__leaf_prog_clk net94 vss vss vdd vdd mem_top_track_0.DFF_2_.Q sky130_fd_sc_hd__dfxtp_1
X_424_ mux_right_track_16.mux_l1_in_1_.TGATE_0_.out _062_ vss vss vdd vdd mux_right_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_286_ _041_ vss vss vdd vdd _062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_95 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 chanx_left_in[4] vss vss vdd vdd net6 sky130_fd_sc_hd__clkbuf_2
X_269_ _035_ vss vss vdd vdd _074_ sky130_fd_sc_hd__clkbuf_1
X_407_ net2 vss vss vdd vdd net46 sky130_fd_sc_hd__clkbuf_1
X_338_ net31 vss vss vdd vdd mux_right_track_8.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_7_109 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput20 chany_top_in[0] vss vss vdd vdd net20 sky130_fd_sc_hd__buf_1
XFILLER_0_17_34 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput31 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net31 sky130_fd_sc_hd__buf_1
XFILLER_0_3_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_126 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_457__69 vss vss vdd vdd net69 _457__69/LO sky130_fd_sc_hd__conb_1
X_371_ clknet_2_2__leaf_prog_clk net85 vss vss vdd vdd mem_top_track_16.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_440_ mux_left_track_17.INVTX1_2_.out _078_ vss vss vdd vdd mux_left_track_17.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_132 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_88 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_423_ net64 _061_ vss vss vdd vdd mux_right_track_16.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_354_ mem_left_track_17.DFF_0_.D vss vss vdd vdd _144_ sky130_fd_sc_hd__inv_2
X_285_ mem_right_track_16.DFF_1_.Q vss vss vdd vdd _041_ sky130_fd_sc_hd__clkbuf_1
XTAP_96 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_left_in[5] vss vss vdd vdd net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_22_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_423__64 vss vss vdd vdd net64 _423__64/LO sky130_fd_sc_hd__conb_1
X_268_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _035_ sky130_fd_sc_hd__clkbuf_1
X_406_ net3 vss vss vdd vdd net47 sky130_fd_sc_hd__clkbuf_1
X_337_ net3 vss vss vdd vdd mux_right_track_8.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_199_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_57 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_17_46 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xinput21 chany_top_in[1] vss vss vdd vdd net21 sky130_fd_sc_hd__buf_1
Xinput32 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_ vss vss vdd vdd
+ net32 sky130_fd_sc_hd__clkbuf_1
Xinput10 chanx_left_in[8] vss vss vdd vdd net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_66 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_465__70 vss vss vdd vdd net70 _465__70/LO sky130_fd_sc_hd__conb_1
XFILLER_0_12_7 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_370_ clknet_2_3__leaf_prog_clk net90 vss vss vdd vdd mem_right_track_0.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_499_ mux_left_track_1.INVTX1_0_.out _137_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_353_ net29 vss vss vdd vdd mux_left_track_9.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_0_17_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_422_ mux_right_track_16.mux_l2_in_1_.TGATE_0_.out _060_ vss vss vdd vdd mux_right_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_284_ _040_ vss vss vdd vdd _064_ sky130_fd_sc_hd__clkbuf_1
Xinput8 chanx_left_in[6] vss vss vdd vdd net8 sky130_fd_sc_hd__buf_1
XTAP_97 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_117 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_267_ mem_left_track_17.DFF_0_.Q vss vss vdd vdd _079_ sky130_fd_sc_hd__inv_2
X_336_ mux_right_track_8.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net49 sky130_fd_sc_hd__inv_2
X_405_ net4 vss vss vdd vdd net48 sky130_fd_sc_hd__clkbuf_1
X_198_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _125_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_100 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_319_ net27 vss vss vdd vdd mux_left_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
Xinput22 chany_top_in[2] vss vss vdd vdd net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ vss vss vdd vdd
+ net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput11 chanx_right_in[0] vss vss vdd vdd net11 sky130_fd_sc_hd__buf_1
XFILLER_0_0_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_498_ mux_left_track_1.INVTX1_2_.out _136_ vss vss vdd vdd mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_421_ mux_top_track_0.mux_l1_in_0_.TGATE_0_.out _059_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_352_ net22 vss vss vdd vdd mux_left_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
Xinput9 chanx_left_in[7] vss vss vdd vdd net9 sky130_fd_sc_hd__clkbuf_1
XTAP_98 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ mem_right_track_16.DFF_0_.Q vss vss vdd vdd _040_ sky130_fd_sc_hd__clkbuf_1
XTAP_65 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ net6 vss vss vdd vdd mux_right_track_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_266_ mem_left_track_17.DFF_1_.Q vss vss vdd vdd _077_ sky130_fd_sc_hd__inv_2
X_404_ net6 vss vss vdd vdd net50 sky130_fd_sc_hd__clkbuf_1
X_197_ mem_right_track_8.DFF_1_.Q vss vss vdd vdd _122_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_47 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_112 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_6_123 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput34 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_ vss vss vdd vdd
+ net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 chany_top_in[3] vss vss vdd vdd net23 sky130_fd_sc_hd__clkbuf_1
X_249_ _029_ vss vss vdd vdd _090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xinput12 chanx_right_in[1] vss vss vdd vdd net12 sky130_fd_sc_hd__buf_1
X_318_ net13 vss vss vdd vdd mux_left_track_17.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_18_91 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold1 mem_right_track_0.DFF_2_.Q vss vss vdd vdd net74 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_91 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_47 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_497_ mux_left_track_1.INVTX1_4_.out _135_ vss vss vdd vdd mux_left_track_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_17_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_420_ mux_top_track_0.INVTX1_2_.out _058_ vss vss vdd vdd mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_351_ net25 vss vss vdd vdd mux_left_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_282_ mem_right_track_16.DFF_0_.Q vss vss vdd vdd _069_ sky130_fd_sc_hd__inv_2
XTAP_99 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_334_ net32 vss vss vdd vdd mux_right_track_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_22_38 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_403_ net7 vss vss vdd vdd net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_59 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_196_ mem_right_track_16.DFF_0_.D vss vss vdd vdd _120_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_135 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_265_ net35 vss vss vdd vdd _075_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_60 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xinput24 chany_top_in[4] vss vss vdd vdd net24 sky130_fd_sc_hd__clkbuf_1
X_248_ mem_top_track_14.DFF_1_.Q vss vss vdd vdd _029_ sky130_fd_sc_hd__clkbuf_1
X_317_ mux_left_track_17.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net44 sky130_fd_sc_hd__inv_2
X_179_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _134_ sky130_fd_sc_hd__inv_2
Xinput13 chanx_right_in[2] vss vss vdd vdd net13 sky130_fd_sc_hd__buf_1
XFILLER_0_23_70 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_119 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_108 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_19_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold2 mem_left_track_17.DFF_0_.D vss vss vdd vdd net75 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_496_ mux_left_track_1.mux_l1_in_0_.TGATE_0_.out _134_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_5_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_350_ net28 vss vss vdd vdd mux_left_track_9.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_281_ mem_right_track_16.DFF_1_.Q vss vss vdd vdd _067_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_106 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_56 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_479_ mux_right_track_8.INVTX1_5_.out _117_ vss vss vdd vdd mux_right_track_8.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_78 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_51 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_264_ _034_ vss vss vdd vdd _081_ sky130_fd_sc_hd__clkbuf_1
XPHY_40 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_402_ net8 vss vss vdd vdd net52 sky130_fd_sc_hd__clkbuf_1
X_333_ net2 vss vss vdd vdd mux_right_track_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_195_ _011_ vss vss vdd vdd _127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput25 chany_top_in[5] vss vss vdd vdd net25 sky130_fd_sc_hd__buf_1
X_247_ _028_ vss vss vdd vdd _091_ sky130_fd_sc_hd__clkbuf_1
X_316_ net8 vss vss vdd vdd mux_right_track_16.INVTX1_4_.out sky130_fd_sc_hd__inv_2
Xinput14 chanx_right_in[3] vss vss vdd vdd net14 sky130_fd_sc_hd__clkbuf_1
X_178_ mem_left_track_1.DFF_2_.Q vss vss vdd vdd _132_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_81 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_477__71 vss vss vdd vdd net71 _477__71/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold3 mem_top_track_14.DFF_0_.D vss vss vdd vdd net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_495_ mux_left_track_1.mux_l1_in_2_.TGATE_0_.out _133_ vss vss vdd vdd mux_left_track_1.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_94 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_280_ mem_left_track_1.DFF_0_.D vss vss vdd vdd _065_ sky130_fd_sc_hd__inv_2
XTAP_57 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_478_ mux_right_track_8.mux_l1_in_1_.TGATE_0_.out _116_ vss vss vdd vdd mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_79 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_263_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_22_18 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_30 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_332_ mux_right_track_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net45 sky130_fd_sc_hd__inv_2
X_194_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _011_ sky130_fd_sc_hd__clkbuf_1
X_401_ net11 vss vss vdd vdd net37 sky130_fd_sc_hd__buf_1
X_501__73 vss vss vdd vdd net73 _501__73/LO sky130_fd_sc_hd__conb_1
XFILLER_0_12_95 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xinput26 chany_top_in[6] vss vss vdd vdd net26 sky130_fd_sc_hd__clkbuf_1
X_246_ mem_top_track_14.DFF_0_.Q vss vss vdd vdd _028_ sky130_fd_sc_hd__clkbuf_1
Xinput15 chanx_right_in[4] vss vss vdd vdd net15 sky130_fd_sc_hd__dlymetal6s2s_1
X_177_ _005_ vss vss vdd vdd _139_ sky130_fd_sc_hd__clkbuf_1
X_315_ net4 vss vss vdd vdd mux_right_track_16.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_229_ _022_ vss vss vdd vdd _105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold4 mem_top_track_0.DFF_2_.Q vss vss vdd vdd net77 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_0_72 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_494_ mux_left_track_1.mux_l2_in_0_.TGATE_0_.out _132_ vss vss vdd vdd mux_left_track_1.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XTAP_58 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_477_ net71 _115_ vss vss vdd vdd mux_right_track_8.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_22_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_130 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_262_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _084_ sky130_fd_sc_hd__inv_2
XPHY_42 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_331_ net9 vss vss vdd vdd mux_top_track_16.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XPHY_31 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_400_ net12 vss vss vdd vdd net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_93 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_193_ _010_ vss vss vdd vdd _129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_18 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput27 chany_top_in[7] vss vss vdd vdd net27 sky130_fd_sc_hd__clkbuf_1
X_245_ mem_top_track_14.DFF_0_.Q vss vss vdd vdd _093_ sky130_fd_sc_hd__inv_2
Xinput16 chanx_right_in[5] vss vss vdd vdd net16 sky130_fd_sc_hd__dlymetal6s2s_1
X_176_ mem_left_track_9.DFF_1_.Q vss vss vdd vdd _005_ sky130_fd_sc_hd__clkbuf_1
X_314_ mux_right_track_16.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net53 sky130_fd_sc_hd__inv_2
XFILLER_0_2_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_228_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _022_ sky130_fd_sc_hd__clkbuf_1
Xhold5 mem_right_track_16.DFF_0_.D vss vss vdd vdd net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_493_ mux_left_track_1.INVTX1_1_.out _131_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_59 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ mux_right_track_8.mux_l2_in_1_.TGATE_0_.out _114_ vss vss vdd vdd mux_right_track_8.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_9_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_54 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_261_ _033_ vss vss vdd vdd _080_ sky130_fd_sc_hd__clkbuf_1
XPHY_43 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_32 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_330_ net14 vss vss vdd vdd mux_top_track_16.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_192_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _010_ sky130_fd_sc_hd__clkbuf_1
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_459_ mux_top_track_16.INVTX1_1_.out _097_ vss vss vdd vdd mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput28 chany_top_in[8] vss vss vdd vdd net28 sky130_fd_sc_hd__clkbuf_1
X_244_ mem_top_track_14.DFF_1_.Q vss vss vdd vdd _092_ sky130_fd_sc_hd__inv_2
Xinput17 chanx_right_in[6] vss vss vdd vdd net17 sky130_fd_sc_hd__dlymetal6s2s_1
X_175_ _004_ vss vss vdd vdd _141_ sky130_fd_sc_hd__clkbuf_1
X_313_ net5 vss vss vdd vdd mux_top_track_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_0_3_51 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_227_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _111_ sky130_fd_sc_hd__inv_2
Xhold6 mem_left_track_1.DFF_0_.D vss vss vdd vdd net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_63 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_26_129 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_492_ mux_left_track_1.INVTX1_3_.out _130_ vss vss vdd vdd mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_475_ mux_left_track_9.INVTX1_0_.out _113_ vss vss vdd vdd mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_55 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_260_ mem_top_track_2.DFF_1_.Q vss vss vdd vdd _033_ sky130_fd_sc_hd__clkbuf_1
XPHY_44 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_33 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_458_ mux_right_track_8.INVTX1_4_.out _096_ vss vss vdd vdd mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_12_21 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_191_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _135_ sky130_fd_sc_hd__inv_2
X_489__72 vss vss vdd vdd net72 _489__72/LO sky130_fd_sc_hd__conb_1
X_312_ net33 vss vss vdd vdd mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
Xinput29 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net29 sky130_fd_sc_hd__clkbuf_1
Xinput18 chanx_right_in[7] vss vss vdd vdd net18 sky130_fd_sc_hd__clkbuf_1
X_174_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _004_ sky130_fd_sc_hd__clkbuf_1
X_243_ _027_ vss vss vdd vdd _095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_226_ mem_right_track_0.DFF_1_.Q vss vss vdd vdd _109_ sky130_fd_sc_hd__inv_2
Xhold7 mem_top_track_14.DFF_0_.Q vss vss vdd vdd net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_54 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_209_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _123_ sky130_fd_sc_hd__inv_2
X_491_ mux_left_track_1.INVTX1_5_.out _129_ vss vss vdd vdd mux_left_track_1.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_25_130 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_474_ mux_left_track_9.INVTX1_2_.out _112_ vss vss vdd vdd mux_right_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_63 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_45 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_34 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_190_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _133_ sky130_fd_sc_hd__inv_2
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_457_ net69 _095_ vss vss vdd vdd mux_top_track_16.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_103 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xinput19 chanx_right_in[8] vss vss vdd vdd net19 sky130_fd_sc_hd__clkbuf_1
X_311_ net18 vss vss vdd vdd mux_top_track_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_173_ mem_left_track_9.DFF_0_.Q vss vss vdd vdd _147_ sky130_fd_sc_hd__inv_2
X_242_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _027_ sky130_fd_sc_hd__clkbuf_1
X_509_ mux_left_track_9.INVTX1_4_.out _147_ vss vss vdd vdd mux_left_track_9.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_225_ _021_ vss vss vdd vdd _102_ sky130_fd_sc_hd__clkbuf_1
Xhold8 mem_right_track_0.DFF_0_.D vss vss vdd vdd net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_44 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_17_6 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_208_ mem_right_track_8.DFF_1_.Q vss vss vdd vdd _121_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_41 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_490_ mux_left_track_1.mux_l1_in_1_.TGATE_0_.out _128_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_3 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_473_ mux_right_track_0.INVTX1_4_.out _111_ vss vss vdd vdd mux_right_track_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_6 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_6_75 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_46 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_456_ mux_top_track_16.mux_l2_in_1_.TGATE_0_.out _094_ vss vss vdd vdd mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_10_115 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_310_ mux_top_track_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net54 sky130_fd_sc_hd__inv_2
XFILLER_0_23_99 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_241_ mem_top_track_16.DFF_1_.Q vss vss vdd vdd _099_ sky130_fd_sc_hd__inv_2
X_508_ mux_left_track_9.mux_l1_in_0_.TGATE_0_.out _146_ vss vss vdd vdd mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_172_ mem_left_track_9.DFF_1_.Q vss vss vdd vdd _145_ sky130_fd_sc_hd__inv_2
X_439_ mux_left_track_17.mux_l1_in_0_.TGATE_0_.out _077_ vss vss vdd vdd mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_224_ mem_right_track_0.DFF_2_.Q vss vss vdd vdd _021_ sky130_fd_sc_hd__clkbuf_1
Xhold9 mem_top_track_14.DFF_1_.Q vss vss vdd vdd net82 sky130_fd_sc_hd__dlygate4sd3_1
X_207_ _015_ vss vss vdd vdd _114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_99 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_25_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_472_ mux_right_track_0.mux_l1_in_0_.TGATE_0_.out _110_ vss vss vdd vdd mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XPHY_47 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_455_ mux_right_track_16.INVTX1_3_.out _093_ vss vss vdd vdd mux_top_track_14.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_127 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_240_ _026_ vss vss vdd vdd _094_ sky130_fd_sc_hd__clkbuf_1
X_171_ _003_ vss vss vdd vdd _138_ sky130_fd_sc_hd__clkbuf_1
X_369_ clknet_2_3__leaf_prog_clk net76 vss vss vdd vdd mem_top_track_14.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_507_ mux_left_track_9.mux_l1_in_2_.TGATE_0_.out _145_ vss vss vdd vdd mux_left_track_9.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_438_ mux_left_track_17.INVTX1_4_.out _076_ vss vss vdd vdd mux_left_track_17.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_88 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_223_ _020_ vss vss vdd vdd _106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_56 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_206_ mem_right_track_16.DFF_0_.D vss vss vdd vdd _015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_45 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_22_6 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_471_ mux_right_track_0.mux_l1_in_2_.TGATE_0_.out _109_ vss vss vdd vdd mux_right_track_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_16_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_48 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_37 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_454_ mux_top_track_14.mux_l1_in_0_.TGATE_0_.out _092_ vss vss vdd vdd mux_top_track_14.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_10_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_100 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_170_ mem_left_track_17.DFF_0_.D vss vss vdd vdd _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_23_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_299_ _045_ vss vss vdd vdd _053_ sky130_fd_sc_hd__clkbuf_1
X_368_ clknet_2_3__leaf_prog_clk net80 vss vss vdd vdd mem_top_track_14.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_506_ mux_left_track_9.mux_l2_in_0_.TGATE_0_.out _144_ vss vss vdd vdd mux_left_track_9.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_437_ mux_left_track_17.mux_l2_in_0_.TGATE_0_.out _075_ vss vss vdd vdd mux_left_track_17.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_222_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_24 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_205_ _014_ vss vss vdd vdd _118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_79 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_22_137 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_470_ mux_right_track_0.mux_l2_in_0_.TGATE_0_.out _108_ vss vss vdd vdd mux_right_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XPHY_49 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_38 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_453_ mux_top_track_14.INVTX1_1_.out _091_ vss vss vdd vdd mux_top_track_14.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_384_ clknet_2_0__leaf_prog_clk net86 vss vss vdd vdd mem_left_track_9.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_6 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_23_47 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_298_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_36 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_505_ mux_left_track_9.INVTX1_1_.out _143_ vss vss vdd vdd mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_367_ clknet_2_3__leaf_prog_clk net83 vss vss vdd vdd mem_top_track_8.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_436_ mux_left_track_17.INVTX1_1_.out _074_ vss vss vdd vdd mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_221_ mem_right_track_0.DFF_0_.Q vss vss vdd vdd _112_ sky130_fd_sc_hd__inv_2
X_419_ mux_top_track_0.INVTX1_0_.out _057_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_204_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_36 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_7 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_28 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_452_ net68 _090_ vss vss vdd vdd mux_top_track_14.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XPHY_39 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_383_ clknet_2_0__leaf_prog_clk net96 vss vss vdd vdd mem_left_track_9.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput60 net60 vss vss vdd vdd chany_top_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_130 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_297_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _057_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_366_ clknet_2_3__leaf_prog_clk net84 vss vss vdd vdd mem_top_track_14.DFF_0_.D sky130_fd_sc_hd__dfxtp_1
X_504_ mux_left_track_9.INVTX1_3_.out _142_ vss vss vdd vdd mux_left_track_9.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_435_ mux_left_track_17.INVTX1_3_.out _073_ vss vss vdd vdd mux_left_track_17.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_220_ _019_ vss vss vdd vdd _104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_37 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_418_ mux_top_track_0.mux_l2_in_0_.TGATE_0_.out _056_ vss vss vdd vdd mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_349_ net12 vss vss vdd vdd mux_left_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_203_ mem_right_track_8.DFF_0_.Q vss vss vdd vdd _124_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_125 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_15_49 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_26_15 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput61 net61 vss vss vdd vdd chany_top_out[7] sky130_fd_sc_hd__clkbuf_4
X_451_ mux_left_track_17.INVTX1_4_.out _089_ vss vss vdd vdd mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_382_ clknet_2_0__leaf_prog_clk net98 vss vss vdd vdd mem_left_track_17.DFF_0_.D
+ sky130_fd_sc_hd__dfxtp_1
Xoutput50 net50 vss vss vdd vdd chanx_right_out[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_17 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_120 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_296_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _059_ sky130_fd_sc_hd__inv_2
X_365_ clknet_2_1__leaf_prog_clk net77 vss vss vdd vdd mem_top_track_2.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_503_ mux_left_track_9.INVTX1_5_.out _141_ vss vss vdd vdd mux_left_track_9.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_434_ mux_left_track_17.mux_l1_in_1_.TGATE_0_.out _072_ vss vss vdd vdd mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_417_ mux_top_track_0.INVTX1_4_.out _055_ vss vss vdd vdd mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_348_ net16 vss vss vdd vdd mux_left_track_9.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_279_ _039_ vss vss vdd vdd _071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_80 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_202_ _013_ vss vss vdd vdd _116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_36 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_72 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_443__66 vss vss vdd vdd net66 _443__66/LO sky130_fd_sc_hd__conb_1
XFILLER_0_21_93 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_26_38 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_6_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput62 net62 vss vss vdd vdd chany_top_out[8] sky130_fd_sc_hd__clkbuf_4
X_450_ mux_top_track_8.mux_l1_in_0_.TGATE_0_.out _088_ vss vss vdd vdd mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xoutput51 net51 vss vss vdd vdd chanx_right_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput40 net40 vss vss vdd vdd chanx_left_out[4] sky130_fd_sc_hd__clkbuf_4
X_381_ clknet_2_2__leaf_prog_clk net79 vss vss vdd vdd mem_left_track_1.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
XTAP_121 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_502_ mux_left_track_9.mux_l1_in_1_.TGATE_0_.out _140_ vss vss vdd vdd mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_2_6 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_433_ net65 _071_ vss vss vdd vdd mux_left_track_17.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_295_ mem_top_track_0.DFF_2_.Q vss vss vdd vdd _056_ sky130_fd_sc_hd__inv_2
X_364_ clknet_2_3__leaf_prog_clk net87 vss vss vdd vdd mem_top_track_2.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_27 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_416_ mux_right_track_0.INVTX1_4_.out _054_ vss vss vdd vdd mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_347_ mux_left_track_9.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net40 sky130_fd_sc_hd__inv_2
X_278_ mem_left_track_17.DFF_1_.Q vss vss vdd vdd _039_ sky130_fd_sc_hd__clkbuf_1
X_201_ mem_right_track_8.DFF_1_.Q vss vss vdd vdd _013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_102 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_25_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xoutput52 net52 vss vss vdd vdd chanx_right_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 vss vss vdd vdd chanx_left_out[5] sky130_fd_sc_hd__clkbuf_4
X_380_ clknet_2_0__leaf_prog_clk net95 vss vss vdd vdd mem_left_track_1.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XTAP_122 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

