magic
tech sky130A
magscale 1 2
timestamp 1708041115
<< viali >>
rect 2053 11305 2087 11339
rect 2513 11305 2547 11339
rect 12449 11305 12483 11339
rect 3617 11237 3651 11271
rect 8401 11237 8435 11271
rect 9873 11237 9907 11271
rect 11345 11237 11379 11271
rect 11713 11237 11747 11271
rect 8953 11169 8987 11203
rect 1501 11101 1535 11135
rect 1777 11101 1811 11135
rect 2237 11101 2271 11135
rect 2605 11095 2639 11129
rect 2881 11101 2915 11135
rect 3433 11101 3467 11135
rect 4629 11101 4663 11135
rect 5825 11101 5859 11135
rect 7021 11101 7055 11135
rect 8217 11101 8251 11135
rect 9137 11101 9171 11135
rect 9689 11101 9723 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 11161 11097 11195 11131
rect 11529 11101 11563 11135
rect 11989 11101 12023 11135
rect 12265 11101 12299 11135
rect 1685 10965 1719 10999
rect 1961 10965 1995 10999
rect 2697 10965 2731 10999
rect 4813 10965 4847 10999
rect 6009 10965 6043 10999
rect 7205 10965 7239 10999
rect 9597 10965 9631 10999
rect 10425 10965 10459 10999
rect 10793 10965 10827 10999
rect 11805 10965 11839 10999
rect 1685 10761 1719 10795
rect 9229 10761 9263 10795
rect 9505 10761 9539 10795
rect 10333 10693 10367 10727
rect 10425 10693 10459 10727
rect 11161 10693 11195 10727
rect 1409 10625 1443 10659
rect 1869 10625 1903 10659
rect 8861 10625 8895 10659
rect 9137 10625 9171 10659
rect 11253 10625 11287 10659
rect 11897 10625 11931 10659
rect 12173 10625 12207 10659
rect 12265 10625 12299 10659
rect 9965 10557 9999 10591
rect 10149 10557 10183 10591
rect 10977 10557 11011 10591
rect 11989 10489 12023 10523
rect 1593 10421 1627 10455
rect 9045 10421 9079 10455
rect 11713 10421 11747 10455
rect 12449 10421 12483 10455
rect 9505 10217 9539 10251
rect 9321 10013 9355 10047
rect 12173 9673 12207 9707
rect 1409 9537 1443 9571
rect 11989 9537 12023 9571
rect 12265 9537 12299 9571
rect 9137 9469 9171 9503
rect 10885 9469 10919 9503
rect 1593 9333 1627 9367
rect 9781 9333 9815 9367
rect 12449 9333 12483 9367
rect 10333 9061 10367 9095
rect 10885 8993 10919 9027
rect 11161 8993 11195 9027
rect 7849 8925 7883 8959
rect 8953 8925 8987 8959
rect 9220 8925 9254 8959
rect 10425 8925 10459 8959
rect 10977 8857 11011 8891
rect 8493 8789 8527 8823
rect 10609 8789 10643 8823
rect 1593 8585 1627 8619
rect 10793 8585 10827 8619
rect 8686 8517 8720 8551
rect 9312 8517 9346 8551
rect 12173 8517 12207 8551
rect 1409 8449 1443 8483
rect 10609 8449 10643 8483
rect 11805 8449 11839 8483
rect 8953 8381 8987 8415
rect 9045 8381 9079 8415
rect 7573 8313 7607 8347
rect 12449 8313 12483 8347
rect 10425 8245 10459 8279
rect 11897 8245 11931 8279
rect 11069 7905 11103 7939
rect 11437 7905 11471 7939
rect 10425 7837 10459 7871
rect 11253 7837 11287 7871
rect 11345 7837 11379 7871
rect 11805 7837 11839 7871
rect 6745 7769 6779 7803
rect 8953 7769 8987 7803
rect 9505 7769 9539 7803
rect 9597 7769 9631 7803
rect 12173 7769 12207 7803
rect 8033 7701 8067 7735
rect 9873 7701 9907 7735
rect 10609 7701 10643 7735
rect 11713 7701 11747 7735
rect 12265 7701 12299 7735
rect 7757 7497 7791 7531
rect 10517 7497 10551 7531
rect 10241 7429 10275 7463
rect 10333 7429 10367 7463
rect 12173 7429 12207 7463
rect 1501 7361 1535 7395
rect 1777 7361 1811 7395
rect 5917 7361 5951 7395
rect 6644 7361 6678 7395
rect 7849 7361 7883 7395
rect 10793 7361 10827 7395
rect 11069 7361 11103 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 6377 7293 6411 7327
rect 11529 7293 11563 7327
rect 9781 7225 9815 7259
rect 1685 7157 1719 7191
rect 1961 7157 1995 7191
rect 6101 7157 6135 7191
rect 9137 7157 9171 7191
rect 10977 7157 11011 7191
rect 7205 6953 7239 6987
rect 8401 6953 8435 6987
rect 12357 6953 12391 6987
rect 9045 6817 9079 6851
rect 1685 6749 1719 6783
rect 1777 6749 1811 6783
rect 4997 6749 5031 6783
rect 5733 6749 5767 6783
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 8493 6749 8527 6783
rect 9312 6749 9346 6783
rect 11161 6749 11195 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 5641 6681 5675 6715
rect 5978 6681 6012 6715
rect 8585 6681 8619 6715
rect 1593 6613 1627 6647
rect 1961 6613 1995 6647
rect 7113 6613 7147 6647
rect 8125 6613 8159 6647
rect 10425 6613 10459 6647
rect 11345 6613 11379 6647
rect 1685 6409 1719 6443
rect 4353 6409 4387 6443
rect 6377 6409 6411 6443
rect 5488 6341 5522 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 2053 6273 2087 6307
rect 2973 6273 3007 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 8697 6273 8731 6307
rect 8953 6273 8987 6307
rect 9137 6273 9171 6307
rect 10241 6273 10275 6307
rect 10517 6273 10551 6307
rect 11713 6273 11747 6307
rect 12265 6273 12299 6307
rect 2237 6205 2271 6239
rect 2881 6205 2915 6239
rect 7021 6205 7055 6239
rect 7113 6205 7147 6239
rect 9597 6205 9631 6239
rect 10701 6205 10735 6239
rect 11529 6205 11563 6239
rect 7573 6137 7607 6171
rect 1961 6069 1995 6103
rect 2697 6069 2731 6103
rect 6101 6069 6135 6103
rect 9321 6069 9355 6103
rect 11161 6069 11195 6103
rect 11897 6069 11931 6103
rect 12449 6069 12483 6103
rect 5733 5865 5767 5899
rect 10333 5865 10367 5899
rect 10793 5865 10827 5899
rect 12357 5865 12391 5899
rect 1777 5797 1811 5831
rect 9597 5797 9631 5831
rect 10609 5797 10643 5831
rect 11253 5797 11287 5831
rect 2421 5729 2455 5763
rect 9873 5729 9907 5763
rect 11529 5729 11563 5763
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2237 5661 2271 5695
rect 7021 5661 7055 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 10425 5661 10459 5695
rect 10701 5661 10735 5695
rect 11069 5661 11103 5695
rect 12081 5661 12115 5695
rect 12173 5661 12207 5695
rect 7205 5593 7239 5627
rect 7297 5593 7331 5627
rect 7849 5593 7883 5627
rect 1593 5525 1627 5559
rect 2881 5525 2915 5559
rect 11989 5525 12023 5559
rect 1593 5321 1627 5355
rect 6653 5321 6687 5355
rect 9321 5321 9355 5355
rect 12173 5321 12207 5355
rect 5549 5253 5583 5287
rect 5641 5253 5675 5287
rect 1409 5185 1443 5219
rect 6469 5185 6503 5219
rect 9229 5185 9263 5219
rect 11989 5185 12023 5219
rect 12265 5185 12299 5219
rect 6101 5049 6135 5083
rect 12449 4981 12483 5015
rect 1409 4097 1443 4131
rect 12265 4097 12299 4131
rect 1593 3893 1627 3927
rect 12449 3893 12483 3927
rect 11989 3485 12023 3519
rect 12541 3485 12575 3519
rect 12081 3349 12115 3383
rect 12357 3349 12391 3383
rect 11805 3145 11839 3179
rect 12173 3077 12207 3111
rect 5917 3009 5951 3043
rect 11897 3009 11931 3043
rect 6101 2805 6135 2839
rect 12449 2805 12483 2839
rect 2145 2397 2179 2431
rect 2973 2397 3007 2431
rect 3341 2397 3375 2431
rect 4629 2397 4663 2431
rect 6469 2397 6503 2431
rect 7205 2397 7239 2431
rect 8493 2397 8527 2431
rect 9781 2397 9815 2431
rect 11069 2397 11103 2431
rect 11529 2397 11563 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 2053 2329 2087 2363
rect 2237 2329 2271 2363
rect 2605 2329 2639 2363
rect 2881 2329 2915 2363
rect 3893 2329 3927 2363
rect 5089 2329 5123 2363
rect 7849 2329 7883 2363
rect 9229 2329 9263 2363
rect 10609 2329 10643 2363
rect 11897 2329 11931 2363
rect 12173 2329 12207 2363
rect 3525 2261 3559 2295
rect 4169 2261 4203 2295
rect 4813 2261 4847 2295
rect 5181 2261 5215 2295
rect 6561 2261 6595 2295
rect 7389 2261 7423 2295
rect 7941 2261 7975 2295
rect 8677 2261 8711 2295
rect 9321 2261 9355 2295
rect 9965 2261 9999 2295
rect 10701 2261 10735 2295
rect 11253 2261 11287 2295
rect 12449 2261 12483 2295
<< metal1 >>
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 12894 11608 12900 11620
rect 11204 11580 12900 11608
rect 11204 11568 11210 11580
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 1104 11450 12880 11472
rect 1104 11398 2422 11450
rect 2474 11398 2486 11450
rect 2538 11398 2550 11450
rect 2602 11398 2614 11450
rect 2666 11398 2678 11450
rect 2730 11398 5366 11450
rect 5418 11398 5430 11450
rect 5482 11398 5494 11450
rect 5546 11398 5558 11450
rect 5610 11398 5622 11450
rect 5674 11398 8310 11450
rect 8362 11398 8374 11450
rect 8426 11398 8438 11450
rect 8490 11398 8502 11450
rect 8554 11398 8566 11450
rect 8618 11398 11254 11450
rect 11306 11398 11318 11450
rect 11370 11398 11382 11450
rect 11434 11398 11446 11450
rect 11498 11398 11510 11450
rect 11562 11398 12880 11450
rect 1104 11376 12880 11398
rect 1026 11296 1032 11348
rect 1084 11296 1090 11348
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2041 11339 2099 11345
rect 2041 11336 2053 11339
rect 1728 11308 2053 11336
rect 1728 11296 1734 11308
rect 2041 11305 2053 11308
rect 2087 11305 2099 11339
rect 2041 11299 2099 11305
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2547 11308 8984 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 1044 11268 1072 11296
rect 1044 11240 2268 11268
rect 934 11160 940 11212
rect 992 11200 998 11212
rect 992 11172 1808 11200
rect 992 11160 998 11172
rect 1486 11092 1492 11144
rect 1544 11092 1550 11144
rect 1780 11141 1808 11172
rect 2240 11141 2268 11240
rect 2332 11240 2774 11268
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2332 11064 2360 11240
rect 2746 11200 2774 11240
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 3605 11271 3663 11277
rect 3605 11268 3617 11271
rect 3384 11240 3617 11268
rect 3384 11228 3390 11240
rect 3605 11237 3617 11240
rect 3651 11237 3663 11271
rect 3605 11231 3663 11237
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 8662 11268 8668 11280
rect 8435 11240 8668 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 8956 11209 8984 11308
rect 12434 11296 12440 11348
rect 12492 11296 12498 11348
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11268 9919 11271
rect 10134 11268 10140 11280
rect 9907 11240 10140 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 11333 11271 11391 11277
rect 10612 11240 11284 11268
rect 8941 11203 8999 11209
rect 2746 11172 8340 11200
rect 2593 11129 2651 11135
rect 2593 11095 2605 11129
rect 2639 11095 2651 11129
rect 2593 11089 2651 11095
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 4614 11092 4620 11144
rect 4672 11092 4678 11144
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 8202 11092 8208 11144
rect 8260 11092 8266 11144
rect 8312 11132 8340 11172
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 10612 11200 10640 11240
rect 8941 11163 8999 11169
rect 9048 11172 10640 11200
rect 11256 11200 11284 11240
rect 11333 11237 11345 11271
rect 11379 11268 11391 11271
rect 11606 11268 11612 11280
rect 11379 11240 11612 11268
rect 11379 11237 11391 11240
rect 11333 11231 11391 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 11701 11271 11759 11277
rect 11701 11237 11713 11271
rect 11747 11268 11759 11271
rect 12066 11268 12072 11280
rect 11747 11240 12072 11268
rect 11747 11237 11759 11240
rect 11701 11231 11759 11237
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 11256 11172 11560 11200
rect 9048 11132 9076 11172
rect 8312 11104 9076 11132
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9456 11104 9689 11132
rect 9456 11092 9462 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 1964 11036 2360 11064
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1762 10996 1768 11008
rect 1719 10968 1768 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 1964 11005 1992 11036
rect 1949 10999 2007 11005
rect 1949 10965 1961 10999
rect 1995 10965 2007 10999
rect 2608 10996 2636 11089
rect 10520 11064 10548 11095
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 11146 11092 11152 11144
rect 11204 11128 11210 11144
rect 11532 11141 11560 11172
rect 11517 11135 11575 11141
rect 11204 11100 11245 11128
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11204 11092 11210 11100
rect 11517 11095 11575 11101
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11977 11135 12035 11141
rect 11977 11132 11989 11135
rect 11756 11104 11989 11132
rect 11756 11092 11762 11104
rect 11977 11101 11989 11104
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 11149 11091 11207 11092
rect 11054 11064 11060 11076
rect 10520 11036 11060 11064
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 12268 11064 12296 11095
rect 11388 11036 12296 11064
rect 11388 11024 11394 11036
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 2608 10968 2697 10996
rect 1949 10959 2007 10965
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 2685 10959 2743 10965
rect 4798 10956 4804 11008
rect 4856 10956 4862 11008
rect 5994 10956 6000 11008
rect 6052 10956 6058 11008
rect 7190 10956 7196 11008
rect 7248 10956 7254 11008
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10192 10968 10425 10996
rect 10192 10956 10198 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 11790 10956 11796 11008
rect 11848 10956 11854 11008
rect 1104 10906 13040 10928
rect 1104 10854 3894 10906
rect 3946 10854 3958 10906
rect 4010 10854 4022 10906
rect 4074 10854 4086 10906
rect 4138 10854 4150 10906
rect 4202 10854 6838 10906
rect 6890 10854 6902 10906
rect 6954 10854 6966 10906
rect 7018 10854 7030 10906
rect 7082 10854 7094 10906
rect 7146 10854 9782 10906
rect 9834 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 12726 10906
rect 12778 10854 12790 10906
rect 12842 10854 12854 10906
rect 12906 10854 12918 10906
rect 12970 10854 12982 10906
rect 13034 10854 13040 10906
rect 1104 10832 13040 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1673 10795 1731 10801
rect 1673 10792 1685 10795
rect 1544 10764 1685 10792
rect 1544 10752 1550 10764
rect 1673 10761 1685 10764
rect 1719 10761 1731 10795
rect 1673 10755 1731 10761
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 9180 10764 9229 10792
rect 9180 10752 9186 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 9582 10792 9588 10804
rect 9539 10764 9588 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11020 10764 11928 10792
rect 11020 10752 11026 10764
rect 9600 10724 9628 10752
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 9600 10696 10333 10724
rect 10321 10693 10333 10696
rect 10367 10693 10379 10727
rect 10321 10687 10379 10693
rect 10413 10727 10471 10733
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 11149 10727 11207 10733
rect 11149 10724 11161 10727
rect 10459 10696 11161 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 11149 10693 11161 10696
rect 11195 10693 11207 10727
rect 11149 10687 11207 10693
rect 11330 10684 11336 10736
rect 11388 10684 11394 10736
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1854 10616 1860 10668
rect 1912 10616 1918 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9122 10656 9128 10668
rect 8895 10628 9128 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11348 10656 11376 10684
rect 11900 10665 11928 10764
rect 11287 10628 11376 10656
rect 11885 10659 11943 10665
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 9950 10548 9956 10600
rect 10008 10548 10014 10600
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 10962 10548 10968 10600
rect 11020 10548 11026 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11256 10588 11284 10619
rect 12158 10616 12164 10668
rect 12216 10616 12222 10668
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 11204 10560 11284 10588
rect 11204 10548 11210 10560
rect 11977 10523 12035 10529
rect 11977 10520 11989 10523
rect 10980 10492 11989 10520
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 9030 10412 9036 10464
rect 9088 10412 9094 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10980 10452 11008 10492
rect 11977 10489 11989 10492
rect 12023 10489 12035 10523
rect 11977 10483 12035 10489
rect 10560 10424 11008 10452
rect 10560 10412 10566 10424
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11112 10424 11713 10452
rect 11112 10412 11118 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 1104 10362 12880 10384
rect 1104 10310 2422 10362
rect 2474 10310 2486 10362
rect 2538 10310 2550 10362
rect 2602 10310 2614 10362
rect 2666 10310 2678 10362
rect 2730 10310 5366 10362
rect 5418 10310 5430 10362
rect 5482 10310 5494 10362
rect 5546 10310 5558 10362
rect 5610 10310 5622 10362
rect 5674 10310 8310 10362
rect 8362 10310 8374 10362
rect 8426 10310 8438 10362
rect 8490 10310 8502 10362
rect 8554 10310 8566 10362
rect 8618 10310 11254 10362
rect 11306 10310 11318 10362
rect 11370 10310 11382 10362
rect 11434 10310 11446 10362
rect 11498 10310 11510 10362
rect 11562 10310 12880 10362
rect 1104 10288 12880 10310
rect 9030 10208 9036 10260
rect 9088 10208 9094 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9950 10248 9956 10260
rect 9539 10220 9956 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 9048 10044 9076 10208
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9048 10016 9321 10044
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 1104 9818 13040 9840
rect 1104 9766 3894 9818
rect 3946 9766 3958 9818
rect 4010 9766 4022 9818
rect 4074 9766 4086 9818
rect 4138 9766 4150 9818
rect 4202 9766 6838 9818
rect 6890 9766 6902 9818
rect 6954 9766 6966 9818
rect 7018 9766 7030 9818
rect 7082 9766 7094 9818
rect 7146 9766 9782 9818
rect 9834 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 12726 9818
rect 12778 9766 12790 9818
rect 12842 9766 12854 9818
rect 12906 9766 12918 9818
rect 12970 9766 12982 9818
rect 13034 9766 13040 9818
rect 1104 9744 13040 9766
rect 12161 9707 12219 9713
rect 12161 9673 12173 9707
rect 12207 9704 12219 9707
rect 12250 9704 12256 9716
rect 12207 9676 12256 9704
rect 12207 9673 12219 9676
rect 12161 9667 12219 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 934 9528 940 9580
rect 992 9568 998 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 992 9540 1409 9568
rect 992 9528 998 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11940 9540 11989 9568
rect 11940 9528 11946 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 12124 9540 12265 9568
rect 12124 9528 12130 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10744 9472 10885 9500
rect 10744 9460 10750 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 2746 9404 12204 9432
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2746 9364 2774 9404
rect 12176 9376 12204 9404
rect 1627 9336 2774 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 12158 9324 12164 9376
rect 12216 9324 12222 9376
rect 12434 9324 12440 9376
rect 12492 9324 12498 9376
rect 1104 9274 12880 9296
rect 1104 9222 2422 9274
rect 2474 9222 2486 9274
rect 2538 9222 2550 9274
rect 2602 9222 2614 9274
rect 2666 9222 2678 9274
rect 2730 9222 5366 9274
rect 5418 9222 5430 9274
rect 5482 9222 5494 9274
rect 5546 9222 5558 9274
rect 5610 9222 5622 9274
rect 5674 9222 8310 9274
rect 8362 9222 8374 9274
rect 8426 9222 8438 9274
rect 8490 9222 8502 9274
rect 8554 9222 8566 9274
rect 8618 9222 11254 9274
rect 11306 9222 11318 9274
rect 11370 9222 11382 9274
rect 11434 9222 11446 9274
rect 11498 9222 11510 9274
rect 11562 9222 12880 9274
rect 1104 9200 12880 9222
rect 11146 9120 11152 9172
rect 11204 9120 11210 9172
rect 10321 9095 10379 9101
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 11164 9092 11192 9120
rect 10367 9064 11192 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 7834 8916 7840 8968
rect 7892 8916 7898 8968
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 9030 8956 9036 8968
rect 8987 8928 9036 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9208 8959 9266 8965
rect 9208 8925 9220 8959
rect 9254 8956 9266 8959
rect 9766 8956 9772 8968
rect 9254 8928 9772 8956
rect 9254 8925 9266 8928
rect 9208 8919 9266 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10428 8965 10456 9064
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10744 8996 10885 9024
rect 10744 8984 10750 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11020 8996 11161 9024
rect 11020 8984 11026 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 1820 8860 10916 8888
rect 1820 8848 1826 8860
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 10594 8780 10600 8832
rect 10652 8780 10658 8832
rect 10888 8820 10916 8860
rect 10962 8848 10968 8900
rect 11020 8848 11026 8900
rect 11698 8820 11704 8832
rect 10888 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 1104 8730 13040 8752
rect 1104 8678 3894 8730
rect 3946 8678 3958 8730
rect 4010 8678 4022 8730
rect 4074 8678 4086 8730
rect 4138 8678 4150 8730
rect 4202 8678 6838 8730
rect 6890 8678 6902 8730
rect 6954 8678 6966 8730
rect 7018 8678 7030 8730
rect 7082 8678 7094 8730
rect 7146 8678 9782 8730
rect 9834 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 12726 8730
rect 12778 8678 12790 8730
rect 12842 8678 12854 8730
rect 12906 8678 12918 8730
rect 12970 8678 12982 8730
rect 13034 8678 13040 8730
rect 1104 8656 13040 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1627 8588 9260 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 8674 8551 8732 8557
rect 8674 8548 8686 8551
rect 8536 8520 8686 8548
rect 8536 8508 8542 8520
rect 8674 8517 8686 8520
rect 8720 8517 8732 8551
rect 8674 8511 8732 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 9122 8480 9128 8492
rect 7576 8452 9128 8480
rect 7576 8353 7604 8452
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9232 8480 9260 8588
rect 10594 8576 10600 8628
rect 10652 8576 10658 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11606 8576 11612 8628
rect 11664 8576 11670 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 9300 8551 9358 8557
rect 9300 8517 9312 8551
rect 9346 8548 9358 8551
rect 10502 8548 10508 8560
rect 9346 8520 10508 8548
rect 9346 8517 9358 8520
rect 9300 8511 9358 8517
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10612 8489 10640 8576
rect 10597 8483 10655 8489
rect 9232 8452 10088 8480
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9030 8412 9036 8424
rect 8987 8384 9036 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8313 7619 8347
rect 10060 8344 10088 8452
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 11624 8480 11652 8576
rect 11716 8548 11744 8576
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 11716 8520 12173 8548
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11624 8452 11805 8480
rect 10597 8443 10655 8449
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11698 8344 11704 8356
rect 10060 8316 11704 8344
rect 7561 8307 7619 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12437 8347 12495 8353
rect 12437 8344 12449 8347
rect 12400 8316 12449 8344
rect 12400 8304 12406 8316
rect 12437 8313 12449 8316
rect 12483 8313 12495 8347
rect 12437 8307 12495 8313
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10192 8248 10425 8276
rect 10192 8236 10198 8248
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 10413 8239 10471 8245
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11885 8279 11943 8285
rect 11885 8276 11897 8279
rect 11204 8248 11897 8276
rect 11204 8236 11210 8248
rect 11885 8245 11897 8248
rect 11931 8245 11943 8279
rect 11885 8239 11943 8245
rect 1104 8186 12880 8208
rect 1104 8134 2422 8186
rect 2474 8134 2486 8186
rect 2538 8134 2550 8186
rect 2602 8134 2614 8186
rect 2666 8134 2678 8186
rect 2730 8134 5366 8186
rect 5418 8134 5430 8186
rect 5482 8134 5494 8186
rect 5546 8134 5558 8186
rect 5610 8134 5622 8186
rect 5674 8134 8310 8186
rect 8362 8134 8374 8186
rect 8426 8134 8438 8186
rect 8490 8134 8502 8186
rect 8554 8134 8566 8186
rect 8618 8134 11254 8186
rect 11306 8134 11318 8186
rect 11370 8134 11382 8186
rect 11434 8134 11446 8186
rect 11498 8134 11510 8186
rect 11562 8134 12880 8186
rect 1104 8112 12880 8134
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 6696 7976 12204 8004
rect 6696 7964 6702 7976
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11425 7939 11483 7945
rect 11425 7936 11437 7939
rect 11103 7908 11437 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 11425 7905 11437 7908
rect 11471 7905 11483 7939
rect 11425 7899 11483 7905
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10192 7840 10425 7868
rect 10192 7828 10198 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 6730 7760 6736 7812
rect 6788 7760 6794 7812
rect 8938 7760 8944 7812
rect 8996 7760 9002 7812
rect 9214 7760 9220 7812
rect 9272 7800 9278 7812
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 9272 7772 9505 7800
rect 9272 7760 9278 7772
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 9493 7763 9551 7769
rect 9582 7760 9588 7812
rect 9640 7760 9646 7812
rect 10428 7800 10456 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11204 7840 11253 7868
rect 11204 7828 11210 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11348 7800 11376 7831
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 12176 7809 12204 7976
rect 10428 7772 11376 7800
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7769 12219 7803
rect 12161 7763 12219 7769
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7708 7704 8033 7732
rect 7708 7692 7714 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 9732 7704 9873 7732
rect 9732 7692 9738 7704
rect 9861 7701 9873 7704
rect 9907 7701 9919 7735
rect 9861 7695 9919 7701
rect 10594 7692 10600 7744
rect 10652 7692 10658 7744
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11664 7704 11713 7732
rect 11664 7692 11670 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11701 7695 11759 7701
rect 12250 7692 12256 7744
rect 12308 7692 12314 7744
rect 1104 7642 13040 7664
rect 1104 7590 3894 7642
rect 3946 7590 3958 7642
rect 4010 7590 4022 7642
rect 4074 7590 4086 7642
rect 4138 7590 4150 7642
rect 4202 7590 6838 7642
rect 6890 7590 6902 7642
rect 6954 7590 6966 7642
rect 7018 7590 7030 7642
rect 7082 7590 7094 7642
rect 7146 7590 9782 7642
rect 9834 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 12726 7642
rect 12778 7590 12790 7642
rect 12842 7590 12854 7642
rect 12906 7590 12918 7642
rect 12970 7590 12982 7642
rect 13034 7590 13040 7642
rect 1104 7568 13040 7590
rect 1578 7488 1584 7540
rect 1636 7488 1642 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 7834 7528 7840 7540
rect 7791 7500 7840 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 9640 7500 10517 7528
rect 9640 7488 9646 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 1596 7392 1624 7488
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10229 7463 10287 7469
rect 10229 7460 10241 7463
rect 10100 7432 10241 7460
rect 10100 7420 10106 7432
rect 10229 7429 10241 7432
rect 10275 7429 10287 7463
rect 10229 7423 10287 7429
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 10367 7432 12173 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 12161 7429 12173 7432
rect 12207 7460 12219 7463
rect 12434 7460 12440 7472
rect 12207 7432 12440 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 1535 7364 1624 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6632 7395 6690 7401
rect 6632 7361 6644 7395
rect 6678 7392 6690 7395
rect 7190 7392 7196 7404
rect 6678 7364 7196 7392
rect 6678 7361 6690 7364
rect 6632 7355 6690 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7708 7364 7849 7392
rect 7708 7352 7714 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 10827 7364 11069 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11195 7364 11713 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 5776 7296 6377 7324
rect 5776 7284 5782 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 10796 7324 10824 7355
rect 6365 7287 6423 7293
rect 8864 7296 10824 7324
rect 11517 7327 11575 7333
rect 8864 7200 8892 7296
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 11606 7324 11612 7336
rect 11563 7296 11612 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 8996 7228 9781 7256
rect 8996 7216 9002 7228
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 1854 7188 1860 7200
rect 1719 7160 1860 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 1946 7148 1952 7200
rect 2004 7148 2010 7200
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 6270 7188 6276 7200
rect 6135 7160 6276 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 8846 7148 8852 7200
rect 8904 7148 8910 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 9088 7160 9137 7188
rect 9088 7148 9094 7160
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11054 7188 11060 7200
rect 11011 7160 11060 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 1104 7098 12880 7120
rect 1104 7046 2422 7098
rect 2474 7046 2486 7098
rect 2538 7046 2550 7098
rect 2602 7046 2614 7098
rect 2666 7046 2678 7098
rect 2730 7046 5366 7098
rect 5418 7046 5430 7098
rect 5482 7046 5494 7098
rect 5546 7046 5558 7098
rect 5610 7046 5622 7098
rect 5674 7046 8310 7098
rect 8362 7046 8374 7098
rect 8426 7046 8438 7098
rect 8490 7046 8502 7098
rect 8554 7046 8566 7098
rect 8618 7046 11254 7098
rect 11306 7046 11318 7098
rect 11370 7046 11382 7098
rect 11434 7046 11446 7098
rect 11498 7046 11510 7098
rect 11562 7046 12880 7098
rect 1104 7024 12880 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 6638 6984 6644 6996
rect 1912 6956 6644 6984
rect 1912 6944 1918 6956
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 7190 6944 7196 6996
rect 7248 6944 7254 6996
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 9214 6984 9220 6996
rect 8435 6956 9220 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12434 6984 12440 6996
rect 12391 6956 12440 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 8846 6916 8852 6928
rect 7852 6888 8852 6916
rect 7852 6848 7880 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 7760 6820 7880 6848
rect 7944 6820 8524 6848
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 1946 6780 1952 6792
rect 1811 6752 1952 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4356 6752 4997 6780
rect 4356 6656 4384 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 7760 6789 7788 6820
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7116 6752 7757 6780
rect 5629 6715 5687 6721
rect 5629 6681 5641 6715
rect 5675 6712 5687 6715
rect 5966 6715 6024 6721
rect 5966 6712 5978 6715
rect 5675 6684 5978 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 5966 6681 5978 6684
rect 6012 6681 6024 6715
rect 5966 6675 6024 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1854 6644 1860 6656
rect 1627 6616 1860 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 1946 6604 1952 6656
rect 2004 6604 2010 6656
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 7116 6653 7144 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7944 6789 7972 6820
rect 8496 6789 8524 6820
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7892 6752 7941 6780
rect 7892 6740 7898 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7929 6743 7987 6749
rect 8128 6752 8217 6780
rect 8128 6653 8156 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 9300 6783 9358 6789
rect 9300 6749 9312 6783
rect 9346 6780 9358 6783
rect 9674 6780 9680 6792
rect 9346 6752 9680 6780
rect 9346 6749 9358 6752
rect 9300 6743 9358 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 8573 6715 8631 6721
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 10060 6712 10088 6808
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 11112 6752 11161 6780
rect 11112 6740 11118 6752
rect 11149 6749 11161 6752
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12084 6712 12112 6743
rect 8619 6684 10088 6712
rect 11348 6684 12112 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6613 7159 6647
rect 7101 6607 7159 6613
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 11348 6653 11376 6684
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 1104 6554 13040 6576
rect 1104 6502 3894 6554
rect 3946 6502 3958 6554
rect 4010 6502 4022 6554
rect 4074 6502 4086 6554
rect 4138 6502 4150 6554
rect 4202 6502 6838 6554
rect 6890 6502 6902 6554
rect 6954 6502 6966 6554
rect 7018 6502 7030 6554
rect 7082 6502 7094 6554
rect 7146 6502 9782 6554
rect 9834 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 12726 6554
rect 12778 6502 12790 6554
rect 12842 6502 12854 6554
rect 12906 6502 12918 6554
rect 12970 6502 12982 6554
rect 13034 6502 13040 6554
rect 1104 6480 13040 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6409 1731 6443
rect 1673 6403 1731 6409
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6273 1547 6307
rect 1688 6304 1716 6403
rect 1854 6400 1860 6452
rect 1912 6400 1918 6452
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 2004 6412 3096 6440
rect 2004 6400 2010 6412
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1688 6276 1777 6304
rect 1489 6267 1547 6273
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1872 6304 1900 6400
rect 2041 6307 2099 6313
rect 2041 6304 2053 6307
rect 1872 6276 2053 6304
rect 1765 6267 1823 6273
rect 2041 6273 2053 6276
rect 2087 6273 2099 6307
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2041 6267 2099 6273
rect 2148 6276 2973 6304
rect 1504 6236 1532 6267
rect 2148 6236 2176 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 1504 6208 2176 6236
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2271 6208 2881 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 2866 6100 2872 6112
rect 2731 6072 2872 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 2976 6100 3004 6267
rect 3068 6168 3096 6412
rect 4338 6400 4344 6452
rect 4396 6400 4402 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5644 6412 6377 6440
rect 4356 6304 4384 6400
rect 5476 6375 5534 6381
rect 5476 6341 5488 6375
rect 5522 6372 5534 6375
rect 5644 6372 5672 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 5522 6344 5672 6372
rect 5736 6344 8984 6372
rect 5522 6341 5534 6344
rect 5476 6335 5534 6341
rect 5736 6316 5764 6344
rect 4356 6276 5672 6304
rect 5644 6236 5672 6276
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 8956 6313 8984 6344
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 8685 6307 8743 6313
rect 8685 6273 8697 6307
rect 8731 6304 8743 6307
rect 8941 6307 8999 6313
rect 8731 6276 8892 6304
rect 8731 6273 8743 6276
rect 8685 6267 8743 6273
rect 5902 6236 5908 6248
rect 5644 6208 5908 6236
rect 5902 6196 5908 6208
rect 5960 6236 5966 6248
rect 6012 6236 6040 6267
rect 5960 6208 6040 6236
rect 7009 6239 7067 6245
rect 5960 6196 5966 6208
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7190 6236 7196 6248
rect 7147 6208 7196 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 4706 6168 4712 6180
rect 3068 6140 4712 6168
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 7024 6168 7052 6199
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 8864 6236 8892 6276
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 10134 6304 10140 6316
rect 9171 6276 10140 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6304 10287 6307
rect 10428 6304 10456 6400
rect 10275 6276 10456 6304
rect 10505 6307 10563 6313
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10594 6304 10600 6316
rect 10551 6276 10600 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 8864 6208 9597 6236
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10520 6236 10548 6267
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11204 6276 11713 6304
rect 11204 6264 11210 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 12250 6264 12256 6316
rect 12308 6264 12314 6316
rect 10376 6208 10548 6236
rect 10376 6196 10382 6208
rect 10686 6196 10692 6248
rect 10744 6196 10750 6248
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 11606 6236 11612 6248
rect 11563 6208 11612 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 5736 6140 7573 6168
rect 5736 6100 5764 6140
rect 7561 6137 7573 6140
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 2976 6072 5764 6100
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 11149 6103 11207 6109
rect 11149 6069 11161 6103
rect 11195 6100 11207 6103
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11195 6072 11897 6100
rect 11195 6069 11207 6072
rect 11149 6063 11207 6069
rect 11885 6069 11897 6072
rect 11931 6100 11943 6103
rect 11974 6100 11980 6112
rect 11931 6072 11980 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12434 6060 12440 6112
rect 12492 6060 12498 6112
rect 1104 6010 12880 6032
rect 1104 5958 2422 6010
rect 2474 5958 2486 6010
rect 2538 5958 2550 6010
rect 2602 5958 2614 6010
rect 2666 5958 2678 6010
rect 2730 5958 5366 6010
rect 5418 5958 5430 6010
rect 5482 5958 5494 6010
rect 5546 5958 5558 6010
rect 5610 5958 5622 6010
rect 5674 5958 8310 6010
rect 8362 5958 8374 6010
rect 8426 5958 8438 6010
rect 8490 5958 8502 6010
rect 8554 5958 8566 6010
rect 8618 5958 11254 6010
rect 11306 5958 11318 6010
rect 11370 5958 11382 6010
rect 11434 5958 11446 6010
rect 11498 5958 11510 6010
rect 11562 5958 12880 6010
rect 1104 5936 12880 5958
rect 1946 5856 1952 5908
rect 2004 5856 2010 5908
rect 5718 5856 5724 5908
rect 5776 5856 5782 5908
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 10410 5856 10416 5908
rect 10468 5856 10474 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10744 5868 10793 5896
rect 10744 5856 10750 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 10781 5859 10839 5865
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 12308 5868 12357 5896
rect 12308 5856 12314 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5797 1823 5831
rect 1765 5791 1823 5797
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 1780 5692 1808 5791
rect 1964 5760 1992 5856
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 1964 5732 2421 5760
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 7650 5760 7656 5772
rect 2409 5723 2467 5729
rect 7024 5732 7656 5760
rect 7024 5701 7052 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 1719 5664 1808 5692
rect 1949 5695 2007 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 9324 5692 9352 5856
rect 9585 5831 9643 5837
rect 9585 5797 9597 5831
rect 9631 5828 9643 5831
rect 9631 5800 9904 5828
rect 9631 5797 9643 5800
rect 9585 5791 9643 5797
rect 9876 5769 9904 5800
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9324 5664 9413 5692
rect 7009 5655 7067 5661
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 1026 5584 1032 5636
rect 1084 5624 1090 5636
rect 1964 5624 1992 5655
rect 1084 5596 1992 5624
rect 1084 5584 1090 5596
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 2240 5556 2268 5655
rect 9674 5652 9680 5704
rect 9732 5652 9738 5704
rect 10428 5701 10456 5856
rect 10597 5831 10655 5837
rect 10597 5797 10609 5831
rect 10643 5797 10655 5831
rect 11164 5828 11192 5856
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 11164 5800 11253 5828
rect 10597 5791 10655 5797
rect 11241 5797 11253 5800
rect 11287 5797 11299 5831
rect 11241 5791 11299 5797
rect 10612 5760 10640 5791
rect 11517 5763 11575 5769
rect 10612 5732 11100 5760
rect 11072 5701 11100 5732
rect 11517 5729 11529 5763
rect 11563 5760 11575 5763
rect 11624 5760 11652 5856
rect 11563 5732 11652 5760
rect 11563 5729 11575 5732
rect 11517 5723 11575 5729
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10459 5664 10701 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11992 5692 12020 5856
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11992 5664 12081 5692
rect 11057 5655 11115 5661
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 4764 5596 5672 5624
rect 4764 5584 4770 5596
rect 1627 5528 2268 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 5534 5556 5540 5568
rect 2924 5528 5540 5556
rect 2924 5516 2930 5528
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5644 5556 5672 5596
rect 7190 5584 7196 5636
rect 7248 5584 7254 5636
rect 7285 5627 7343 5633
rect 7285 5593 7297 5627
rect 7331 5624 7343 5627
rect 7374 5624 7380 5636
rect 7331 5596 7380 5624
rect 7331 5593 7343 5596
rect 7285 5587 7343 5593
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 7834 5584 7840 5636
rect 7892 5584 7898 5636
rect 11054 5556 11060 5568
rect 5644 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11974 5516 11980 5568
rect 12032 5516 12038 5568
rect 1104 5466 13040 5488
rect 1104 5414 3894 5466
rect 3946 5414 3958 5466
rect 4010 5414 4022 5466
rect 4074 5414 4086 5466
rect 4138 5414 4150 5466
rect 4202 5414 6838 5466
rect 6890 5414 6902 5466
rect 6954 5414 6966 5466
rect 7018 5414 7030 5466
rect 7082 5414 7094 5466
rect 7146 5414 9782 5466
rect 9834 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 12726 5466
rect 12778 5414 12790 5466
rect 12842 5414 12854 5466
rect 12906 5414 12918 5466
rect 12970 5414 12982 5466
rect 13034 5414 13040 5466
rect 1104 5392 13040 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1627 5324 2774 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2746 5080 2774 5324
rect 6086 5312 6092 5364
rect 6144 5312 6150 5364
rect 6270 5312 6276 5364
rect 6328 5312 6334 5364
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 7374 5352 7380 5364
rect 6687 5324 7380 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 9309 5355 9367 5361
rect 9309 5321 9321 5355
rect 9355 5352 9367 5355
rect 9674 5352 9680 5364
rect 9355 5324 9680 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 5534 5244 5540 5296
rect 5592 5244 5598 5296
rect 5629 5287 5687 5293
rect 5629 5253 5641 5287
rect 5675 5284 5687 5287
rect 6104 5284 6132 5312
rect 5675 5256 6132 5284
rect 5675 5253 5687 5256
rect 5629 5247 5687 5253
rect 6288 5216 6316 5312
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6288 5188 6469 5216
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9232 5148 9260 5179
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11756 5188 11989 5216
rect 11756 5176 11762 5188
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 12176 5216 12204 5315
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12176 5188 12265 5216
rect 11977 5179 12035 5185
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 5644 5120 9260 5148
rect 5644 5080 5672 5120
rect 2746 5052 5672 5080
rect 6089 5083 6147 5089
rect 6089 5049 6101 5083
rect 6135 5080 6147 5083
rect 7834 5080 7840 5092
rect 6135 5052 7840 5080
rect 6135 5049 6147 5052
rect 6089 5043 6147 5049
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 12434 4972 12440 5024
rect 12492 4972 12498 5024
rect 1104 4922 12880 4944
rect 1104 4870 2422 4922
rect 2474 4870 2486 4922
rect 2538 4870 2550 4922
rect 2602 4870 2614 4922
rect 2666 4870 2678 4922
rect 2730 4870 5366 4922
rect 5418 4870 5430 4922
rect 5482 4870 5494 4922
rect 5546 4870 5558 4922
rect 5610 4870 5622 4922
rect 5674 4870 8310 4922
rect 8362 4870 8374 4922
rect 8426 4870 8438 4922
rect 8490 4870 8502 4922
rect 8554 4870 8566 4922
rect 8618 4870 11254 4922
rect 11306 4870 11318 4922
rect 11370 4870 11382 4922
rect 11434 4870 11446 4922
rect 11498 4870 11510 4922
rect 11562 4870 12880 4922
rect 1104 4848 12880 4870
rect 1104 4378 13040 4400
rect 1104 4326 3894 4378
rect 3946 4326 3958 4378
rect 4010 4326 4022 4378
rect 4074 4326 4086 4378
rect 4138 4326 4150 4378
rect 4202 4326 6838 4378
rect 6890 4326 6902 4378
rect 6954 4326 6966 4378
rect 7018 4326 7030 4378
rect 7082 4326 7094 4378
rect 7146 4326 9782 4378
rect 9834 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 12726 4378
rect 12778 4326 12790 4378
rect 12842 4326 12854 4378
rect 12906 4326 12918 4378
rect 12970 4326 12982 4378
rect 13034 4326 13040 4378
rect 1104 4304 13040 4326
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 992 4100 1409 4128
rect 992 4088 998 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 11112 4100 12265 4128
rect 11112 4088 11118 4100
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 11790 3924 11796 3936
rect 1627 3896 11796 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12434 3884 12440 3936
rect 12492 3884 12498 3936
rect 1104 3834 12880 3856
rect 1104 3782 2422 3834
rect 2474 3782 2486 3834
rect 2538 3782 2550 3834
rect 2602 3782 2614 3834
rect 2666 3782 2678 3834
rect 2730 3782 5366 3834
rect 5418 3782 5430 3834
rect 5482 3782 5494 3834
rect 5546 3782 5558 3834
rect 5610 3782 5622 3834
rect 5674 3782 8310 3834
rect 8362 3782 8374 3834
rect 8426 3782 8438 3834
rect 8490 3782 8502 3834
rect 8554 3782 8566 3834
rect 8618 3782 11254 3834
rect 11306 3782 11318 3834
rect 11370 3782 11382 3834
rect 11434 3782 11446 3834
rect 11498 3782 11510 3834
rect 11562 3782 12880 3834
rect 1104 3760 12880 3782
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 7892 3488 11989 3516
rect 7892 3476 7898 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12575 3488 12664 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12636 3392 12664 3488
rect 12066 3340 12072 3392
rect 12124 3340 12130 3392
rect 12342 3340 12348 3392
rect 12400 3340 12406 3392
rect 12618 3340 12624 3392
rect 12676 3340 12682 3392
rect 1104 3290 13040 3312
rect 1104 3238 3894 3290
rect 3946 3238 3958 3290
rect 4010 3238 4022 3290
rect 4074 3238 4086 3290
rect 4138 3238 4150 3290
rect 4202 3238 6838 3290
rect 6890 3238 6902 3290
rect 6954 3238 6966 3290
rect 7018 3238 7030 3290
rect 7082 3238 7094 3290
rect 7146 3238 9782 3290
rect 9834 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 12726 3290
rect 12778 3238 12790 3290
rect 12842 3238 12854 3290
rect 12906 3238 12918 3290
rect 12970 3238 12982 3290
rect 13034 3238 13040 3290
rect 1104 3216 13040 3238
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 11882 3176 11888 3188
rect 11839 3148 11888 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12124 3148 12204 3176
rect 12124 3136 12130 3148
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6012 3040 6040 3136
rect 12176 3117 12204 3148
rect 12342 3136 12348 3188
rect 12400 3136 12406 3188
rect 12161 3111 12219 3117
rect 12161 3077 12173 3111
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 5951 3012 6040 3040
rect 11885 3043 11943 3049
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12360 3040 12388 3136
rect 11931 3012 12388 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 6086 2796 6092 2848
rect 6144 2796 6150 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 12400 2808 12449 2836
rect 12400 2796 12406 2808
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 1104 2746 12880 2768
rect 1104 2694 2422 2746
rect 2474 2694 2486 2746
rect 2538 2694 2550 2746
rect 2602 2694 2614 2746
rect 2666 2694 2678 2746
rect 2730 2694 5366 2746
rect 5418 2694 5430 2746
rect 5482 2694 5494 2746
rect 5546 2694 5558 2746
rect 5610 2694 5622 2746
rect 5674 2694 8310 2746
rect 8362 2694 8374 2746
rect 8426 2694 8438 2746
rect 8490 2694 8502 2746
rect 8554 2694 8566 2746
rect 8618 2694 11254 2746
rect 11306 2694 11318 2746
rect 11370 2694 11382 2746
rect 11434 2694 11446 2746
rect 11498 2694 11510 2746
rect 11562 2694 12880 2746
rect 1104 2672 12880 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 6730 2632 6736 2644
rect 3476 2604 6736 2632
rect 3476 2592 3482 2604
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 10870 2564 10876 2576
rect 2976 2536 10876 2564
rect 2976 2437 3004 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 8938 2496 8944 2508
rect 3436 2468 8944 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 750 2320 756 2372
rect 808 2360 814 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 808 2332 1409 2360
rect 808 2320 814 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 2041 2363 2099 2369
rect 2041 2360 2053 2363
rect 1811 2332 2053 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 2041 2329 2053 2332
rect 2087 2329 2099 2363
rect 2041 2323 2099 2329
rect 2148 2292 2176 2391
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 2222 2320 2228 2372
rect 2280 2320 2286 2372
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 2869 2363 2927 2369
rect 2869 2360 2881 2363
rect 2639 2332 2881 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 2869 2329 2881 2332
rect 2915 2329 2927 2363
rect 2869 2323 2927 2329
rect 3436 2292 3464 2468
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 6144 2400 6469 2428
rect 6144 2388 6150 2400
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 10318 2428 10324 2440
rect 9815 2400 10324 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 10836 2400 11069 2428
rect 10836 2388 10842 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2428 11575 2431
rect 12434 2428 12440 2440
rect 11563 2400 12440 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3528 2332 3893 2360
rect 3528 2301 3556 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2329 5135 2363
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 5077 2323 5135 2329
rect 7392 2332 7849 2360
rect 2148 2264 3464 2292
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2261 3571 2295
rect 3513 2255 3571 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3844 2264 4169 2292
rect 3844 2252 3850 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 5092 2292 5120 2323
rect 4847 2264 5120 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 5166 2252 5172 2304
rect 5224 2252 5230 2304
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 7392 2301 7420 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 7837 2323 7895 2329
rect 8680 2332 9229 2360
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6328 2264 6561 2292
rect 6328 2252 6334 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 7377 2295 7435 2301
rect 7377 2261 7389 2295
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 8680 2301 8708 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 10597 2363 10655 2369
rect 10597 2329 10609 2363
rect 10643 2329 10655 2363
rect 10597 2323 10655 2329
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7708 2264 7941 2292
rect 7708 2252 7714 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 10612 2292 10640 2323
rect 11882 2320 11888 2372
rect 11940 2320 11946 2372
rect 12161 2363 12219 2369
rect 12161 2360 12173 2363
rect 11992 2332 12173 2360
rect 9999 2264 10640 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 10686 2252 10692 2304
rect 10744 2252 10750 2304
rect 11241 2295 11299 2301
rect 11241 2261 11253 2295
rect 11287 2292 11299 2295
rect 11992 2292 12020 2332
rect 12161 2329 12173 2332
rect 12207 2329 12219 2363
rect 12161 2323 12219 2329
rect 11287 2264 12020 2292
rect 11287 2261 11299 2264
rect 11241 2255 11299 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12124 2264 12449 2292
rect 12124 2252 12130 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 1104 2202 13040 2224
rect 1104 2150 3894 2202
rect 3946 2150 3958 2202
rect 4010 2150 4022 2202
rect 4074 2150 4086 2202
rect 4138 2150 4150 2202
rect 4202 2150 6838 2202
rect 6890 2150 6902 2202
rect 6954 2150 6966 2202
rect 7018 2150 7030 2202
rect 7082 2150 7094 2202
rect 7146 2150 9782 2202
rect 9834 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 12726 2202
rect 12778 2150 12790 2202
rect 12842 2150 12854 2202
rect 12906 2150 12918 2202
rect 12970 2150 12982 2202
rect 13034 2150 13040 2202
rect 1104 2128 13040 2150
<< via1 >>
rect 11152 11568 11204 11620
rect 12900 11568 12952 11620
rect 2422 11398 2474 11450
rect 2486 11398 2538 11450
rect 2550 11398 2602 11450
rect 2614 11398 2666 11450
rect 2678 11398 2730 11450
rect 5366 11398 5418 11450
rect 5430 11398 5482 11450
rect 5494 11398 5546 11450
rect 5558 11398 5610 11450
rect 5622 11398 5674 11450
rect 8310 11398 8362 11450
rect 8374 11398 8426 11450
rect 8438 11398 8490 11450
rect 8502 11398 8554 11450
rect 8566 11398 8618 11450
rect 11254 11398 11306 11450
rect 11318 11398 11370 11450
rect 11382 11398 11434 11450
rect 11446 11398 11498 11450
rect 11510 11398 11562 11450
rect 1032 11296 1084 11348
rect 1676 11296 1728 11348
rect 940 11160 992 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 3332 11228 3384 11280
rect 8668 11228 8720 11280
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 10140 11228 10192 11280
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 11612 11228 11664 11280
rect 12072 11228 12124 11280
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9404 11092 9456 11144
rect 1768 10956 1820 11008
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 11152 11131 11204 11144
rect 11152 11097 11161 11131
rect 11161 11097 11195 11131
rect 11195 11097 11204 11131
rect 11152 11092 11204 11097
rect 11704 11092 11756 11144
rect 11060 11024 11112 11076
rect 11336 11024 11388 11076
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 9588 10999 9640 11008
rect 9588 10965 9597 10999
rect 9597 10965 9631 10999
rect 9631 10965 9640 10999
rect 9588 10956 9640 10965
rect 10140 10956 10192 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 11796 10999 11848 11008
rect 11796 10965 11805 10999
rect 11805 10965 11839 10999
rect 11839 10965 11848 10999
rect 11796 10956 11848 10965
rect 3894 10854 3946 10906
rect 3958 10854 4010 10906
rect 4022 10854 4074 10906
rect 4086 10854 4138 10906
rect 4150 10854 4202 10906
rect 6838 10854 6890 10906
rect 6902 10854 6954 10906
rect 6966 10854 7018 10906
rect 7030 10854 7082 10906
rect 7094 10854 7146 10906
rect 9782 10854 9834 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 12726 10854 12778 10906
rect 12790 10854 12842 10906
rect 12854 10854 12906 10906
rect 12918 10854 12970 10906
rect 12982 10854 13034 10906
rect 1492 10752 1544 10804
rect 9128 10752 9180 10804
rect 9588 10752 9640 10804
rect 10968 10752 11020 10804
rect 11336 10684 11388 10736
rect 940 10616 992 10668
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11152 10548 11204 10600
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 10508 10412 10560 10464
rect 11060 10412 11112 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 2422 10310 2474 10362
rect 2486 10310 2538 10362
rect 2550 10310 2602 10362
rect 2614 10310 2666 10362
rect 2678 10310 2730 10362
rect 5366 10310 5418 10362
rect 5430 10310 5482 10362
rect 5494 10310 5546 10362
rect 5558 10310 5610 10362
rect 5622 10310 5674 10362
rect 8310 10310 8362 10362
rect 8374 10310 8426 10362
rect 8438 10310 8490 10362
rect 8502 10310 8554 10362
rect 8566 10310 8618 10362
rect 11254 10310 11306 10362
rect 11318 10310 11370 10362
rect 11382 10310 11434 10362
rect 11446 10310 11498 10362
rect 11510 10310 11562 10362
rect 9036 10208 9088 10260
rect 9956 10208 10008 10260
rect 3894 9766 3946 9818
rect 3958 9766 4010 9818
rect 4022 9766 4074 9818
rect 4086 9766 4138 9818
rect 4150 9766 4202 9818
rect 6838 9766 6890 9818
rect 6902 9766 6954 9818
rect 6966 9766 7018 9818
rect 7030 9766 7082 9818
rect 7094 9766 7146 9818
rect 9782 9766 9834 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 12726 9766 12778 9818
rect 12790 9766 12842 9818
rect 12854 9766 12906 9818
rect 12918 9766 12970 9818
rect 12982 9766 13034 9818
rect 12256 9664 12308 9716
rect 940 9528 992 9580
rect 11888 9528 11940 9580
rect 12072 9528 12124 9580
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 10692 9460 10744 9512
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 12164 9324 12216 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 2422 9222 2474 9274
rect 2486 9222 2538 9274
rect 2550 9222 2602 9274
rect 2614 9222 2666 9274
rect 2678 9222 2730 9274
rect 5366 9222 5418 9274
rect 5430 9222 5482 9274
rect 5494 9222 5546 9274
rect 5558 9222 5610 9274
rect 5622 9222 5674 9274
rect 8310 9222 8362 9274
rect 8374 9222 8426 9274
rect 8438 9222 8490 9274
rect 8502 9222 8554 9274
rect 8566 9222 8618 9274
rect 11254 9222 11306 9274
rect 11318 9222 11370 9274
rect 11382 9222 11434 9274
rect 11446 9222 11498 9274
rect 11510 9222 11562 9274
rect 11152 9120 11204 9172
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 9036 8916 9088 8968
rect 9772 8916 9824 8968
rect 10692 8984 10744 9036
rect 10968 8984 11020 9036
rect 1768 8848 1820 8900
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 10968 8891 11020 8900
rect 10968 8857 10977 8891
rect 10977 8857 11011 8891
rect 11011 8857 11020 8891
rect 10968 8848 11020 8857
rect 11704 8780 11756 8832
rect 3894 8678 3946 8730
rect 3958 8678 4010 8730
rect 4022 8678 4074 8730
rect 4086 8678 4138 8730
rect 4150 8678 4202 8730
rect 6838 8678 6890 8730
rect 6902 8678 6954 8730
rect 6966 8678 7018 8730
rect 7030 8678 7082 8730
rect 7094 8678 7146 8730
rect 9782 8678 9834 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 12726 8678 12778 8730
rect 12790 8678 12842 8730
rect 12854 8678 12906 8730
rect 12918 8678 12970 8730
rect 12982 8678 13034 8730
rect 8484 8508 8536 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 9128 8440 9180 8492
rect 10600 8576 10652 8628
rect 10968 8576 11020 8628
rect 11612 8576 11664 8628
rect 11704 8576 11756 8628
rect 10508 8508 10560 8560
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 11704 8304 11756 8356
rect 12348 8304 12400 8356
rect 10140 8236 10192 8288
rect 11152 8236 11204 8288
rect 2422 8134 2474 8186
rect 2486 8134 2538 8186
rect 2550 8134 2602 8186
rect 2614 8134 2666 8186
rect 2678 8134 2730 8186
rect 5366 8134 5418 8186
rect 5430 8134 5482 8186
rect 5494 8134 5546 8186
rect 5558 8134 5610 8186
rect 5622 8134 5674 8186
rect 8310 8134 8362 8186
rect 8374 8134 8426 8186
rect 8438 8134 8490 8186
rect 8502 8134 8554 8186
rect 8566 8134 8618 8186
rect 11254 8134 11306 8186
rect 11318 8134 11370 8186
rect 11382 8134 11434 8186
rect 11446 8134 11498 8186
rect 11510 8134 11562 8186
rect 6644 7964 6696 8016
rect 10140 7828 10192 7880
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 8944 7803 8996 7812
rect 8944 7769 8953 7803
rect 8953 7769 8987 7803
rect 8987 7769 8996 7803
rect 8944 7760 8996 7769
rect 9220 7760 9272 7812
rect 9588 7803 9640 7812
rect 9588 7769 9597 7803
rect 9597 7769 9631 7803
rect 9631 7769 9640 7803
rect 9588 7760 9640 7769
rect 11152 7828 11204 7880
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 7656 7692 7708 7744
rect 9680 7692 9732 7744
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 11612 7692 11664 7744
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 3894 7590 3946 7642
rect 3958 7590 4010 7642
rect 4022 7590 4074 7642
rect 4086 7590 4138 7642
rect 4150 7590 4202 7642
rect 6838 7590 6890 7642
rect 6902 7590 6954 7642
rect 6966 7590 7018 7642
rect 7030 7590 7082 7642
rect 7094 7590 7146 7642
rect 9782 7590 9834 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 12726 7590 12778 7642
rect 12790 7590 12842 7642
rect 12854 7590 12906 7642
rect 12918 7590 12970 7642
rect 12982 7590 13034 7642
rect 1584 7488 1636 7540
rect 7840 7488 7892 7540
rect 9588 7488 9640 7540
rect 10048 7420 10100 7472
rect 12440 7420 12492 7472
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 7196 7352 7248 7404
rect 7656 7352 7708 7404
rect 5724 7284 5776 7336
rect 11612 7284 11664 7336
rect 8944 7216 8996 7268
rect 1860 7148 1912 7200
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 6276 7148 6328 7200
rect 8852 7148 8904 7200
rect 9036 7148 9088 7200
rect 11060 7148 11112 7200
rect 2422 7046 2474 7098
rect 2486 7046 2538 7098
rect 2550 7046 2602 7098
rect 2614 7046 2666 7098
rect 2678 7046 2730 7098
rect 5366 7046 5418 7098
rect 5430 7046 5482 7098
rect 5494 7046 5546 7098
rect 5558 7046 5610 7098
rect 5622 7046 5674 7098
rect 8310 7046 8362 7098
rect 8374 7046 8426 7098
rect 8438 7046 8490 7098
rect 8502 7046 8554 7098
rect 8566 7046 8618 7098
rect 11254 7046 11306 7098
rect 11318 7046 11370 7098
rect 11382 7046 11434 7098
rect 11446 7046 11498 7098
rect 11510 7046 11562 7098
rect 1860 6944 1912 6996
rect 6644 6944 6696 6996
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 9220 6944 9272 6996
rect 12440 6944 12492 6996
rect 8852 6876 8904 6928
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 1952 6740 2004 6792
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 1860 6604 1912 6656
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 4344 6604 4396 6656
rect 7840 6740 7892 6792
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 10048 6808 10100 6860
rect 9680 6740 9732 6792
rect 11060 6740 11112 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 3894 6502 3946 6554
rect 3958 6502 4010 6554
rect 4022 6502 4074 6554
rect 4086 6502 4138 6554
rect 4150 6502 4202 6554
rect 6838 6502 6890 6554
rect 6902 6502 6954 6554
rect 6966 6502 7018 6554
rect 7030 6502 7082 6554
rect 7094 6502 7146 6554
rect 9782 6502 9834 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 12726 6502 12778 6554
rect 12790 6502 12842 6554
rect 12854 6502 12906 6554
rect 12918 6502 12970 6554
rect 12982 6502 13034 6554
rect 1860 6400 1912 6452
rect 1952 6400 2004 6452
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2872 6060 2924 6112
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 10416 6400 10468 6452
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5908 6196 5960 6248
rect 4712 6128 4764 6180
rect 7196 6196 7248 6248
rect 10140 6264 10192 6316
rect 10324 6196 10376 6248
rect 10600 6264 10652 6316
rect 11152 6264 11204 6316
rect 12256 6307 12308 6316
rect 12256 6273 12265 6307
rect 12265 6273 12299 6307
rect 12299 6273 12308 6307
rect 12256 6264 12308 6273
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 11612 6196 11664 6248
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 11980 6060 12032 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 2422 5958 2474 6010
rect 2486 5958 2538 6010
rect 2550 5958 2602 6010
rect 2614 5958 2666 6010
rect 2678 5958 2730 6010
rect 5366 5958 5418 6010
rect 5430 5958 5482 6010
rect 5494 5958 5546 6010
rect 5558 5958 5610 6010
rect 5622 5958 5674 6010
rect 8310 5958 8362 6010
rect 8374 5958 8426 6010
rect 8438 5958 8490 6010
rect 8502 5958 8554 6010
rect 8566 5958 8618 6010
rect 11254 5958 11306 6010
rect 11318 5958 11370 6010
rect 11382 5958 11434 6010
rect 11446 5958 11498 6010
rect 11510 5958 11562 6010
rect 1952 5856 2004 5908
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 9312 5856 9364 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 10416 5856 10468 5908
rect 10692 5856 10744 5908
rect 11152 5856 11204 5908
rect 11612 5856 11664 5908
rect 11980 5856 12032 5908
rect 12256 5856 12308 5908
rect 7656 5720 7708 5772
rect 1032 5584 1084 5636
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 4712 5584 4764 5636
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 5540 5516 5592 5568
rect 7196 5627 7248 5636
rect 7196 5593 7205 5627
rect 7205 5593 7239 5627
rect 7239 5593 7248 5627
rect 7196 5584 7248 5593
rect 7380 5584 7432 5636
rect 7840 5627 7892 5636
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 11060 5516 11112 5568
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 3894 5414 3946 5466
rect 3958 5414 4010 5466
rect 4022 5414 4074 5466
rect 4086 5414 4138 5466
rect 4150 5414 4202 5466
rect 6838 5414 6890 5466
rect 6902 5414 6954 5466
rect 6966 5414 7018 5466
rect 7030 5414 7082 5466
rect 7094 5414 7146 5466
rect 9782 5414 9834 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 12726 5414 12778 5466
rect 12790 5414 12842 5466
rect 12854 5414 12906 5466
rect 12918 5414 12970 5466
rect 12982 5414 13034 5466
rect 940 5176 992 5228
rect 6092 5312 6144 5364
rect 6276 5312 6328 5364
rect 7380 5312 7432 5364
rect 9680 5312 9732 5364
rect 5540 5287 5592 5296
rect 5540 5253 5549 5287
rect 5549 5253 5583 5287
rect 5583 5253 5592 5287
rect 5540 5244 5592 5253
rect 11704 5176 11756 5228
rect 7840 5040 7892 5092
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 2422 4870 2474 4922
rect 2486 4870 2538 4922
rect 2550 4870 2602 4922
rect 2614 4870 2666 4922
rect 2678 4870 2730 4922
rect 5366 4870 5418 4922
rect 5430 4870 5482 4922
rect 5494 4870 5546 4922
rect 5558 4870 5610 4922
rect 5622 4870 5674 4922
rect 8310 4870 8362 4922
rect 8374 4870 8426 4922
rect 8438 4870 8490 4922
rect 8502 4870 8554 4922
rect 8566 4870 8618 4922
rect 11254 4870 11306 4922
rect 11318 4870 11370 4922
rect 11382 4870 11434 4922
rect 11446 4870 11498 4922
rect 11510 4870 11562 4922
rect 3894 4326 3946 4378
rect 3958 4326 4010 4378
rect 4022 4326 4074 4378
rect 4086 4326 4138 4378
rect 4150 4326 4202 4378
rect 6838 4326 6890 4378
rect 6902 4326 6954 4378
rect 6966 4326 7018 4378
rect 7030 4326 7082 4378
rect 7094 4326 7146 4378
rect 9782 4326 9834 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 12726 4326 12778 4378
rect 12790 4326 12842 4378
rect 12854 4326 12906 4378
rect 12918 4326 12970 4378
rect 12982 4326 13034 4378
rect 940 4088 992 4140
rect 11060 4088 11112 4140
rect 11796 3884 11848 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 2422 3782 2474 3834
rect 2486 3782 2538 3834
rect 2550 3782 2602 3834
rect 2614 3782 2666 3834
rect 2678 3782 2730 3834
rect 5366 3782 5418 3834
rect 5430 3782 5482 3834
rect 5494 3782 5546 3834
rect 5558 3782 5610 3834
rect 5622 3782 5674 3834
rect 8310 3782 8362 3834
rect 8374 3782 8426 3834
rect 8438 3782 8490 3834
rect 8502 3782 8554 3834
rect 8566 3782 8618 3834
rect 11254 3782 11306 3834
rect 11318 3782 11370 3834
rect 11382 3782 11434 3834
rect 11446 3782 11498 3834
rect 11510 3782 11562 3834
rect 7840 3476 7892 3528
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 12348 3383 12400 3392
rect 12348 3349 12357 3383
rect 12357 3349 12391 3383
rect 12391 3349 12400 3383
rect 12348 3340 12400 3349
rect 12624 3340 12676 3392
rect 3894 3238 3946 3290
rect 3958 3238 4010 3290
rect 4022 3238 4074 3290
rect 4086 3238 4138 3290
rect 4150 3238 4202 3290
rect 6838 3238 6890 3290
rect 6902 3238 6954 3290
rect 6966 3238 7018 3290
rect 7030 3238 7082 3290
rect 7094 3238 7146 3290
rect 9782 3238 9834 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 12726 3238 12778 3290
rect 12790 3238 12842 3290
rect 12854 3238 12906 3290
rect 12918 3238 12970 3290
rect 12982 3238 13034 3290
rect 6000 3136 6052 3188
rect 11888 3136 11940 3188
rect 12072 3136 12124 3188
rect 12348 3136 12400 3188
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 12348 2796 12400 2848
rect 2422 2694 2474 2746
rect 2486 2694 2538 2746
rect 2550 2694 2602 2746
rect 2614 2694 2666 2746
rect 2678 2694 2730 2746
rect 5366 2694 5418 2746
rect 5430 2694 5482 2746
rect 5494 2694 5546 2746
rect 5558 2694 5610 2746
rect 5622 2694 5674 2746
rect 8310 2694 8362 2746
rect 8374 2694 8426 2746
rect 8438 2694 8490 2746
rect 8502 2694 8554 2746
rect 8566 2694 8618 2746
rect 11254 2694 11306 2746
rect 11318 2694 11370 2746
rect 11382 2694 11434 2746
rect 11446 2694 11498 2746
rect 11510 2694 11562 2746
rect 3424 2592 3476 2644
rect 6736 2592 6788 2644
rect 10876 2524 10928 2576
rect 756 2320 808 2372
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 8944 2456 8996 2508
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 6092 2388 6144 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 10324 2388 10376 2440
rect 10784 2388 10836 2440
rect 12440 2388 12492 2440
rect 3792 2252 3844 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 6276 2252 6328 2304
rect 7656 2252 7708 2304
rect 9036 2252 9088 2304
rect 11888 2363 11940 2372
rect 11888 2329 11897 2363
rect 11897 2329 11931 2363
rect 11931 2329 11940 2363
rect 11888 2320 11940 2329
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 12072 2252 12124 2304
rect 3894 2150 3946 2202
rect 3958 2150 4010 2202
rect 4022 2150 4074 2202
rect 4086 2150 4138 2202
rect 4150 2150 4202 2202
rect 6838 2150 6890 2202
rect 6902 2150 6954 2202
rect 6966 2150 7018 2202
rect 7030 2150 7082 2202
rect 7094 2150 7146 2202
rect 9782 2150 9834 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 12726 2150 12778 2202
rect 12790 2150 12842 2202
rect 12854 2150 12906 2202
rect 12918 2150 12970 2202
rect 12982 2150 13034 2202
<< metal2 >>
rect 938 13200 994 14000
rect 2134 13200 2190 14000
rect 2240 13246 2728 13274
rect 952 12458 980 13200
rect 2148 13138 2176 13200
rect 2240 13138 2268 13246
rect 2148 13110 2268 13138
rect 952 12430 1072 12458
rect 938 12336 994 12345
rect 938 12271 994 12280
rect 952 11218 980 12271
rect 1044 11354 1072 12430
rect 2700 11642 2728 13246
rect 3330 13200 3386 14000
rect 4526 13200 4582 14000
rect 5722 13200 5778 14000
rect 6918 13200 6974 14000
rect 8114 13200 8170 14000
rect 9310 13200 9366 14000
rect 10506 13200 10562 14000
rect 10966 13424 11022 13433
rect 10966 13359 11022 13368
rect 3344 12434 3372 13200
rect 4540 12434 4568 13200
rect 5736 12434 5764 13200
rect 6932 12434 6960 13200
rect 8128 12434 8156 13200
rect 3344 12406 3464 12434
rect 4540 12406 4660 12434
rect 5736 12406 5856 12434
rect 6932 12406 7052 12434
rect 8128 12406 8248 12434
rect 2700 11614 2912 11642
rect 2422 11452 2730 11461
rect 2422 11450 2428 11452
rect 2484 11450 2508 11452
rect 2564 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2730 11452
rect 2484 11398 2486 11450
rect 2666 11398 2668 11450
rect 2422 11396 2428 11398
rect 2484 11396 2508 11398
rect 2564 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2730 11398
rect 2422 11387 2730 11396
rect 1032 11348 1084 11354
rect 1032 11290 1084 11296
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 940 11212 992 11218
rect 940 11154 992 11160
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10810 1532 11086
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10169 980 10610
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 952 9081 980 9522
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1596 7546 1624 10406
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 6798 1716 11290
rect 2884 11150 2912 11614
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 2872 11144 2924 11150
rect 1858 11112 1914 11121
rect 2872 11086 2924 11092
rect 1858 11047 1914 11056
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 8906 1808 10950
rect 1872 10674 1900 11047
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2422 10364 2730 10373
rect 2422 10362 2428 10364
rect 2484 10362 2508 10364
rect 2564 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2730 10364
rect 2484 10310 2486 10362
rect 2666 10310 2668 10362
rect 2422 10308 2428 10310
rect 2484 10308 2508 10310
rect 2564 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2730 10310
rect 2422 10299 2730 10308
rect 2422 9276 2730 9285
rect 2422 9274 2428 9276
rect 2484 9274 2508 9276
rect 2564 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2730 9276
rect 2484 9222 2486 9274
rect 2666 9222 2668 9274
rect 2422 9220 2428 9222
rect 2484 9220 2508 9222
rect 2564 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2730 9222
rect 2422 9211 2730 9220
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 2422 8188 2730 8197
rect 2422 8186 2428 8188
rect 2484 8186 2508 8188
rect 2564 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2730 8188
rect 2484 8134 2486 8186
rect 2666 8134 2668 8186
rect 2422 8132 2428 8134
rect 2484 8132 2508 8134
rect 2564 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2730 8134
rect 2422 8123 2730 8132
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 6905 1808 7346
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1872 7002 1900 7142
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1964 6798 1992 7142
rect 2422 7100 2730 7109
rect 2422 7098 2428 7100
rect 2484 7098 2508 7100
rect 2564 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2730 7100
rect 2484 7046 2486 7098
rect 2666 7046 2668 7098
rect 2422 7044 2428 7046
rect 2484 7044 2508 7046
rect 2564 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2730 7046
rect 2422 7035 2730 7044
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1872 6458 1900 6598
rect 1964 6458 1992 6598
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 1964 5914 1992 6054
rect 2422 6012 2730 6021
rect 2422 6010 2428 6012
rect 2484 6010 2508 6012
rect 2564 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2730 6012
rect 2484 5958 2486 6010
rect 2666 5958 2668 6010
rect 2422 5956 2428 5958
rect 2484 5956 2508 5958
rect 2564 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2730 5958
rect 2422 5947 2730 5956
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1030 5808 1086 5817
rect 1030 5743 1086 5752
rect 1044 5642 1072 5743
rect 1032 5636 1084 5642
rect 1032 5578 1084 5584
rect 2884 5574 2912 6054
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4729 980 5170
rect 2422 4924 2730 4933
rect 2422 4922 2428 4924
rect 2484 4922 2508 4924
rect 2564 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2730 4924
rect 2484 4870 2486 4922
rect 2666 4870 2668 4922
rect 2422 4868 2428 4870
rect 2484 4868 2508 4870
rect 2564 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2730 4870
rect 2422 4859 2730 4868
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3641 980 4082
rect 2422 3836 2730 3845
rect 2422 3834 2428 3836
rect 2484 3834 2508 3836
rect 2564 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2730 3836
rect 2484 3782 2486 3834
rect 2666 3782 2668 3834
rect 2422 3780 2428 3782
rect 2484 3780 2508 3782
rect 2564 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2730 3782
rect 2422 3771 2730 3780
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 2422 2748 2730 2757
rect 2422 2746 2428 2748
rect 2484 2746 2508 2748
rect 2564 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2730 2748
rect 2484 2694 2486 2746
rect 2666 2694 2668 2746
rect 2422 2692 2428 2694
rect 2484 2692 2508 2694
rect 2564 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2730 2694
rect 2422 2683 2730 2692
rect 3344 2446 3372 11222
rect 3436 11150 3464 12406
rect 4632 11150 4660 12406
rect 5366 11452 5674 11461
rect 5366 11450 5372 11452
rect 5428 11450 5452 11452
rect 5508 11450 5532 11452
rect 5588 11450 5612 11452
rect 5668 11450 5674 11452
rect 5428 11398 5430 11450
rect 5610 11398 5612 11450
rect 5366 11396 5372 11398
rect 5428 11396 5452 11398
rect 5508 11396 5532 11398
rect 5588 11396 5612 11398
rect 5668 11396 5674 11398
rect 5366 11387 5674 11396
rect 5828 11150 5856 12406
rect 7024 11150 7052 12406
rect 8220 11150 8248 12406
rect 8310 11452 8618 11461
rect 8310 11450 8316 11452
rect 8372 11450 8396 11452
rect 8452 11450 8476 11452
rect 8532 11450 8556 11452
rect 8612 11450 8618 11452
rect 8372 11398 8374 11450
rect 8554 11398 8556 11450
rect 8310 11396 8316 11398
rect 8372 11396 8396 11398
rect 8452 11396 8476 11398
rect 8532 11396 8556 11398
rect 8612 11396 8618 11398
rect 8310 11387 8618 11396
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 3894 10908 4202 10917
rect 3894 10906 3900 10908
rect 3956 10906 3980 10908
rect 4036 10906 4060 10908
rect 4116 10906 4140 10908
rect 4196 10906 4202 10908
rect 3956 10854 3958 10906
rect 4138 10854 4140 10906
rect 3894 10852 3900 10854
rect 3956 10852 3980 10854
rect 4036 10852 4060 10854
rect 4116 10852 4140 10854
rect 4196 10852 4202 10854
rect 3894 10843 4202 10852
rect 3894 9820 4202 9829
rect 3894 9818 3900 9820
rect 3956 9818 3980 9820
rect 4036 9818 4060 9820
rect 4116 9818 4140 9820
rect 4196 9818 4202 9820
rect 3956 9766 3958 9818
rect 4138 9766 4140 9818
rect 3894 9764 3900 9766
rect 3956 9764 3980 9766
rect 4036 9764 4060 9766
rect 4116 9764 4140 9766
rect 4196 9764 4202 9766
rect 3894 9755 4202 9764
rect 3894 8732 4202 8741
rect 3894 8730 3900 8732
rect 3956 8730 3980 8732
rect 4036 8730 4060 8732
rect 4116 8730 4140 8732
rect 4196 8730 4202 8732
rect 3956 8678 3958 8730
rect 4138 8678 4140 8730
rect 3894 8676 3900 8678
rect 3956 8676 3980 8678
rect 4036 8676 4060 8678
rect 4116 8676 4140 8678
rect 4196 8676 4202 8678
rect 3894 8667 4202 8676
rect 3894 7644 4202 7653
rect 3894 7642 3900 7644
rect 3956 7642 3980 7644
rect 4036 7642 4060 7644
rect 4116 7642 4140 7644
rect 4196 7642 4202 7644
rect 3956 7590 3958 7642
rect 4138 7590 4140 7642
rect 3894 7588 3900 7590
rect 3956 7588 3980 7590
rect 4036 7588 4060 7590
rect 4116 7588 4140 7590
rect 4196 7588 4202 7590
rect 3894 7579 4202 7588
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 3894 6556 4202 6565
rect 3894 6554 3900 6556
rect 3956 6554 3980 6556
rect 4036 6554 4060 6556
rect 4116 6554 4140 6556
rect 4196 6554 4202 6556
rect 3956 6502 3958 6554
rect 4138 6502 4140 6554
rect 3894 6500 3900 6502
rect 3956 6500 3980 6502
rect 4036 6500 4060 6502
rect 4116 6500 4140 6502
rect 4196 6500 4202 6502
rect 3894 6491 4202 6500
rect 4356 6458 4384 6598
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5642 4752 6122
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 3894 5468 4202 5477
rect 3894 5466 3900 5468
rect 3956 5466 3980 5468
rect 4036 5466 4060 5468
rect 4116 5466 4140 5468
rect 4196 5466 4202 5468
rect 3956 5414 3958 5466
rect 4138 5414 4140 5466
rect 3894 5412 3900 5414
rect 3956 5412 3980 5414
rect 4036 5412 4060 5414
rect 4116 5412 4140 5414
rect 4196 5412 4202 5414
rect 3894 5403 4202 5412
rect 3894 4380 4202 4389
rect 3894 4378 3900 4380
rect 3956 4378 3980 4380
rect 4036 4378 4060 4380
rect 4116 4378 4140 4380
rect 4196 4378 4202 4380
rect 3956 4326 3958 4378
rect 4138 4326 4140 4378
rect 3894 4324 3900 4326
rect 3956 4324 3980 4326
rect 4036 4324 4060 4326
rect 4116 4324 4140 4326
rect 4196 4324 4202 4326
rect 3894 4315 4202 4324
rect 3894 3292 4202 3301
rect 3894 3290 3900 3292
rect 3956 3290 3980 3292
rect 4036 3290 4060 3292
rect 4116 3290 4140 3292
rect 4196 3290 4202 3292
rect 3956 3238 3958 3290
rect 4138 3238 4140 3290
rect 3894 3236 3900 3238
rect 3956 3236 3980 3238
rect 4036 3236 4060 3238
rect 4116 3236 4140 3238
rect 4196 3236 4202 3238
rect 3894 3227 4202 3236
rect 4816 2774 4844 10950
rect 5366 10364 5674 10373
rect 5366 10362 5372 10364
rect 5428 10362 5452 10364
rect 5508 10362 5532 10364
rect 5588 10362 5612 10364
rect 5668 10362 5674 10364
rect 5428 10310 5430 10362
rect 5610 10310 5612 10362
rect 5366 10308 5372 10310
rect 5428 10308 5452 10310
rect 5508 10308 5532 10310
rect 5588 10308 5612 10310
rect 5668 10308 5674 10310
rect 5366 10299 5674 10308
rect 5366 9276 5674 9285
rect 5366 9274 5372 9276
rect 5428 9274 5452 9276
rect 5508 9274 5532 9276
rect 5588 9274 5612 9276
rect 5668 9274 5674 9276
rect 5428 9222 5430 9274
rect 5610 9222 5612 9274
rect 5366 9220 5372 9222
rect 5428 9220 5452 9222
rect 5508 9220 5532 9222
rect 5588 9220 5612 9222
rect 5668 9220 5674 9222
rect 5366 9211 5674 9220
rect 5366 8188 5674 8197
rect 5366 8186 5372 8188
rect 5428 8186 5452 8188
rect 5508 8186 5532 8188
rect 5588 8186 5612 8188
rect 5668 8186 5674 8188
rect 5428 8134 5430 8186
rect 5610 8134 5612 8186
rect 5366 8132 5372 8134
rect 5428 8132 5452 8134
rect 5508 8132 5532 8134
rect 5588 8132 5612 8134
rect 5668 8132 5674 8134
rect 5366 8123 5674 8132
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5366 7100 5674 7109
rect 5366 7098 5372 7100
rect 5428 7098 5452 7100
rect 5508 7098 5532 7100
rect 5588 7098 5612 7100
rect 5668 7098 5674 7100
rect 5428 7046 5430 7098
rect 5610 7046 5612 7098
rect 5366 7044 5372 7046
rect 5428 7044 5452 7046
rect 5508 7044 5532 7046
rect 5588 7044 5612 7046
rect 5668 7044 5674 7046
rect 5366 7035 5674 7044
rect 5736 6798 5764 7278
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6322 5764 6734
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5366 6012 5674 6021
rect 5366 6010 5372 6012
rect 5428 6010 5452 6012
rect 5508 6010 5532 6012
rect 5588 6010 5612 6012
rect 5668 6010 5674 6012
rect 5428 5958 5430 6010
rect 5610 5958 5612 6010
rect 5366 5956 5372 5958
rect 5428 5956 5452 5958
rect 5508 5956 5532 5958
rect 5588 5956 5612 5958
rect 5668 5956 5674 5958
rect 5366 5947 5674 5956
rect 5736 5914 5764 6258
rect 5920 6254 5948 7346
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5302 5580 5510
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5366 4924 5674 4933
rect 5366 4922 5372 4924
rect 5428 4922 5452 4924
rect 5508 4922 5532 4924
rect 5588 4922 5612 4924
rect 5668 4922 5674 4924
rect 5428 4870 5430 4922
rect 5610 4870 5612 4922
rect 5366 4868 5372 4870
rect 5428 4868 5452 4870
rect 5508 4868 5532 4870
rect 5588 4868 5612 4870
rect 5668 4868 5674 4870
rect 5366 4859 5674 4868
rect 5366 3836 5674 3845
rect 5366 3834 5372 3836
rect 5428 3834 5452 3836
rect 5508 3834 5532 3836
rect 5588 3834 5612 3836
rect 5668 3834 5674 3836
rect 5428 3782 5430 3834
rect 5610 3782 5612 3834
rect 5366 3780 5372 3782
rect 5428 3780 5452 3782
rect 5508 3780 5532 3782
rect 5588 3780 5612 3782
rect 5668 3780 5674 3782
rect 5366 3771 5674 3780
rect 6012 3194 6040 10950
rect 6838 10908 7146 10917
rect 6838 10906 6844 10908
rect 6900 10906 6924 10908
rect 6980 10906 7004 10908
rect 7060 10906 7084 10908
rect 7140 10906 7146 10908
rect 6900 10854 6902 10906
rect 7082 10854 7084 10906
rect 6838 10852 6844 10854
rect 6900 10852 6924 10854
rect 6980 10852 7004 10854
rect 7060 10852 7084 10854
rect 7140 10852 7146 10854
rect 6838 10843 7146 10852
rect 6838 9820 7146 9829
rect 6838 9818 6844 9820
rect 6900 9818 6924 9820
rect 6980 9818 7004 9820
rect 7060 9818 7084 9820
rect 7140 9818 7146 9820
rect 6900 9766 6902 9818
rect 7082 9766 7084 9818
rect 6838 9764 6844 9766
rect 6900 9764 6924 9766
rect 6980 9764 7004 9766
rect 7060 9764 7084 9766
rect 7140 9764 7146 9766
rect 6838 9755 7146 9764
rect 6838 8732 7146 8741
rect 6838 8730 6844 8732
rect 6900 8730 6924 8732
rect 6980 8730 7004 8732
rect 7060 8730 7084 8732
rect 7140 8730 7146 8732
rect 6900 8678 6902 8730
rect 7082 8678 7084 8730
rect 6838 8676 6844 8678
rect 6900 8676 6924 8678
rect 6980 8676 7004 8678
rect 7060 8676 7084 8678
rect 7140 8676 7146 8678
rect 6838 8667 7146 8676
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5370 6132 6054
rect 6288 5370 6316 7142
rect 6656 7002 6684 7958
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 4632 2746 4844 2774
rect 5366 2748 5674 2757
rect 5366 2746 5372 2748
rect 5428 2746 5452 2748
rect 5508 2746 5532 2748
rect 5588 2746 5612 2748
rect 5668 2746 5674 2748
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3436 2553 3464 2586
rect 3422 2544 3478 2553
rect 3422 2479 3478 2488
rect 4632 2446 4660 2746
rect 5428 2694 5430 2746
rect 5610 2694 5612 2746
rect 5366 2692 5372 2694
rect 5428 2692 5452 2694
rect 5508 2692 5532 2694
rect 5588 2692 5612 2694
rect 5668 2692 5674 2694
rect 5366 2683 5674 2692
rect 6104 2446 6132 2790
rect 6748 2650 6776 7754
rect 6838 7644 7146 7653
rect 6838 7642 6844 7644
rect 6900 7642 6924 7644
rect 6980 7642 7004 7644
rect 7060 7642 7084 7644
rect 7140 7642 7146 7644
rect 6900 7590 6902 7642
rect 7082 7590 7084 7642
rect 6838 7588 6844 7590
rect 6900 7588 6924 7590
rect 6980 7588 7004 7590
rect 7060 7588 7084 7590
rect 7140 7588 7146 7590
rect 6838 7579 7146 7588
rect 7208 7562 7236 10950
rect 8310 10364 8618 10373
rect 8310 10362 8316 10364
rect 8372 10362 8396 10364
rect 8452 10362 8476 10364
rect 8532 10362 8556 10364
rect 8612 10362 8618 10364
rect 8372 10310 8374 10362
rect 8554 10310 8556 10362
rect 8310 10308 8316 10310
rect 8372 10308 8396 10310
rect 8452 10308 8476 10310
rect 8532 10308 8556 10310
rect 8612 10308 8618 10310
rect 8310 10299 8618 10308
rect 8310 9276 8618 9285
rect 8310 9274 8316 9276
rect 8372 9274 8396 9276
rect 8452 9274 8476 9276
rect 8532 9274 8556 9276
rect 8612 9274 8618 9276
rect 8372 9222 8374 9274
rect 8554 9222 8556 9274
rect 8310 9220 8316 9222
rect 8372 9220 8396 9222
rect 8452 9220 8476 9222
rect 8532 9220 8556 9222
rect 8612 9220 8618 9222
rect 8310 9211 8618 9220
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7208 7534 7328 7562
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7208 7002 7236 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 6838 6556 7146 6565
rect 6838 6554 6844 6556
rect 6900 6554 6924 6556
rect 6980 6554 7004 6556
rect 7060 6554 7084 6556
rect 7140 6554 7146 6556
rect 6900 6502 6902 6554
rect 7082 6502 7084 6554
rect 6838 6500 6844 6502
rect 6900 6500 6924 6502
rect 6980 6500 7004 6502
rect 7060 6500 7084 6502
rect 7140 6500 7146 6502
rect 6838 6491 7146 6500
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5642 7236 6190
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6838 5468 7146 5477
rect 6838 5466 6844 5468
rect 6900 5466 6924 5468
rect 6980 5466 7004 5468
rect 7060 5466 7084 5468
rect 7140 5466 7146 5468
rect 6900 5414 6902 5466
rect 7082 5414 7084 5466
rect 6838 5412 6844 5414
rect 6900 5412 6924 5414
rect 6980 5412 7004 5414
rect 7060 5412 7084 5414
rect 7140 5412 7146 5414
rect 6838 5403 7146 5412
rect 6838 4380 7146 4389
rect 6838 4378 6844 4380
rect 6900 4378 6924 4380
rect 6980 4378 7004 4380
rect 7060 4378 7084 4380
rect 7140 4378 7146 4380
rect 6900 4326 6902 4378
rect 7082 4326 7084 4378
rect 6838 4324 6844 4326
rect 6900 4324 6924 4326
rect 6980 4324 7004 4326
rect 7060 4324 7084 4326
rect 7140 4324 7146 4326
rect 6838 4315 7146 4324
rect 6838 3292 7146 3301
rect 6838 3290 6844 3292
rect 6900 3290 6924 3292
rect 6980 3290 7004 3292
rect 7060 3290 7084 3292
rect 7140 3290 7146 3292
rect 6900 3238 6902 3290
rect 7082 3238 7084 3290
rect 6838 3236 6844 3238
rect 6900 3236 6924 3238
rect 6980 3236 7004 3238
rect 7060 3236 7084 3238
rect 7140 3236 7146 3238
rect 6838 3227 7146 3236
rect 7300 2774 7328 7534
rect 7668 7410 7696 7686
rect 7852 7546 7880 8910
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8566 8524 8774
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8310 8188 8618 8197
rect 8310 8186 8316 8188
rect 8372 8186 8396 8188
rect 8452 8186 8476 8188
rect 8532 8186 8556 8188
rect 8612 8186 8618 8188
rect 8372 8134 8374 8186
rect 8554 8134 8556 8186
rect 8310 8132 8316 8134
rect 8372 8132 8396 8134
rect 8452 8132 8476 8134
rect 8532 8132 8556 8134
rect 8612 8132 8618 8134
rect 8310 8123 8618 8132
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 5778 7696 7346
rect 7852 6798 7880 7482
rect 8310 7100 8618 7109
rect 8310 7098 8316 7100
rect 8372 7098 8396 7100
rect 8452 7098 8476 7100
rect 8532 7098 8556 7100
rect 8612 7098 8618 7100
rect 8372 7046 8374 7098
rect 8554 7046 8556 7098
rect 8310 7044 8316 7046
rect 8372 7044 8396 7046
rect 8452 7044 8476 7046
rect 8532 7044 8556 7046
rect 8612 7044 8618 7046
rect 8310 7035 8618 7044
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8310 6012 8618 6021
rect 8310 6010 8316 6012
rect 8372 6010 8396 6012
rect 8452 6010 8476 6012
rect 8532 6010 8556 6012
rect 8612 6010 8618 6012
rect 8372 5958 8374 6010
rect 8554 5958 8556 6010
rect 8310 5956 8316 5958
rect 8372 5956 8396 5958
rect 8452 5956 8476 5958
rect 8532 5956 8556 5958
rect 8612 5956 8618 5958
rect 8310 5947 8618 5956
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7392 5370 7420 5578
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7852 5098 7880 5578
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7852 3534 7880 5034
rect 8310 4924 8618 4933
rect 8310 4922 8316 4924
rect 8372 4922 8396 4924
rect 8452 4922 8476 4924
rect 8532 4922 8556 4924
rect 8612 4922 8618 4924
rect 8372 4870 8374 4922
rect 8554 4870 8556 4922
rect 8310 4868 8316 4870
rect 8372 4868 8396 4870
rect 8452 4868 8476 4870
rect 8532 4868 8556 4870
rect 8612 4868 8618 4870
rect 8310 4859 8618 4868
rect 8310 3836 8618 3845
rect 8310 3834 8316 3836
rect 8372 3834 8396 3836
rect 8452 3834 8476 3836
rect 8532 3834 8556 3836
rect 8612 3834 8618 3836
rect 8372 3782 8374 3834
rect 8554 3782 8556 3834
rect 8310 3780 8316 3782
rect 8372 3780 8396 3782
rect 8452 3780 8476 3782
rect 8532 3780 8556 3782
rect 8612 3780 8618 3782
rect 8310 3771 8618 3780
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7208 2746 7328 2774
rect 8310 2748 8618 2757
rect 8310 2746 8316 2748
rect 8372 2746 8396 2748
rect 8452 2746 8476 2748
rect 8532 2746 8556 2748
rect 8612 2746 8618 2748
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7208 2446 7236 2746
rect 8372 2694 8374 2746
rect 8554 2694 8556 2746
rect 8310 2692 8316 2694
rect 8372 2692 8396 2694
rect 8452 2692 8476 2694
rect 8532 2692 8556 2694
rect 8612 2692 8618 2694
rect 8310 2683 8618 2692
rect 8680 2632 8708 11222
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9324 11098 9352 13200
rect 10520 12434 10548 13200
rect 10520 12406 10640 12434
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 9404 11144 9456 11150
rect 9324 11092 9404 11098
rect 9324 11086 9456 11092
rect 10152 11098 10180 11222
rect 10612 11150 10640 12406
rect 10600 11144 10652 11150
rect 9140 10810 9168 11086
rect 9324 11070 9444 11086
rect 10152 11070 10272 11098
rect 10600 11086 10652 11092
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9600 10810 9628 10950
rect 9782 10908 10090 10917
rect 9782 10906 9788 10908
rect 9844 10906 9868 10908
rect 9924 10906 9948 10908
rect 10004 10906 10028 10908
rect 10084 10906 10090 10908
rect 9844 10854 9846 10906
rect 10026 10854 10028 10906
rect 9782 10852 9788 10854
rect 9844 10852 9868 10854
rect 9924 10852 9948 10854
rect 10004 10852 10028 10854
rect 10084 10852 10090 10854
rect 9782 10843 10090 10852
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10266 9076 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9140 9518 9168 10610
rect 10152 10606 10180 10950
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9968 10266 9996 10542
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9782 9820 10090 9829
rect 9782 9818 9788 9820
rect 9844 9818 9868 9820
rect 9924 9818 9948 9820
rect 10004 9818 10028 9820
rect 10084 9818 10090 9820
rect 9844 9766 9846 9818
rect 10026 9766 10028 9818
rect 9782 9764 9788 9766
rect 9844 9764 9868 9766
rect 9924 9764 9948 9766
rect 10004 9764 10028 9766
rect 10084 9764 10090 9766
rect 9782 9755 10090 9764
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8430 9076 8910
rect 9140 8498 9168 9454
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 8974 9812 9318
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9782 8732 10090 8741
rect 9782 8730 9788 8732
rect 9844 8730 9868 8732
rect 9924 8730 9948 8732
rect 10004 8730 10028 8732
rect 10084 8730 10090 8732
rect 9844 8678 9846 8730
rect 10026 8678 10028 8730
rect 9782 8676 9788 8678
rect 9844 8676 9868 8678
rect 9924 8676 9948 8678
rect 10004 8676 10028 8678
rect 10084 8676 10090 8678
rect 9782 8667 10090 8676
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8956 7274 8984 7754
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 6934 8892 7142
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8496 2604 8708 2632
rect 8496 2446 8524 2604
rect 8956 2514 8984 7210
rect 9048 7206 9076 8366
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 7886 10180 8230
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6866 9076 7142
rect 9232 7002 9260 7754
rect 9600 7546 9628 7754
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9692 6798 9720 7686
rect 9782 7644 10090 7653
rect 9782 7642 9788 7644
rect 9844 7642 9868 7644
rect 9924 7642 9948 7644
rect 10004 7642 10028 7644
rect 10084 7642 10090 7644
rect 9844 7590 9846 7642
rect 10026 7590 10028 7642
rect 9782 7588 9788 7590
rect 9844 7588 9868 7590
rect 9924 7588 9948 7590
rect 10004 7588 10028 7590
rect 10084 7588 10090 7590
rect 9782 7579 10090 7588
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 6866 10088 7414
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9782 6556 10090 6565
rect 9782 6554 9788 6556
rect 9844 6554 9868 6556
rect 9924 6554 9948 6556
rect 10004 6554 10028 6556
rect 10084 6554 10090 6556
rect 9844 6502 9846 6554
rect 10026 6502 10028 6554
rect 9782 6500 9788 6502
rect 9844 6500 9868 6502
rect 9924 6500 9948 6502
rect 10004 6500 10028 6502
rect 10084 6500 10090 6502
rect 9782 6491 10090 6500
rect 10152 6322 10180 7822
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 5914 9352 6054
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 5370 9720 5646
rect 9782 5468 10090 5477
rect 9782 5466 9788 5468
rect 9844 5466 9868 5468
rect 9924 5466 9948 5468
rect 10004 5466 10028 5468
rect 10084 5466 10090 5468
rect 9844 5414 9846 5466
rect 10026 5414 10028 5466
rect 9782 5412 9788 5414
rect 9844 5412 9868 5414
rect 9924 5412 9948 5414
rect 10004 5412 10028 5414
rect 10084 5412 10090 5414
rect 9782 5403 10090 5412
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9782 4380 10090 4389
rect 9782 4378 9788 4380
rect 9844 4378 9868 4380
rect 9924 4378 9948 4380
rect 10004 4378 10028 4380
rect 10084 4378 10090 4380
rect 9844 4326 9846 4378
rect 10026 4326 10028 4378
rect 9782 4324 9788 4326
rect 9844 4324 9868 4326
rect 9924 4324 9948 4326
rect 10004 4324 10028 4326
rect 10084 4324 10090 4326
rect 9782 4315 10090 4324
rect 9782 3292 10090 3301
rect 9782 3290 9788 3292
rect 9844 3290 9868 3292
rect 9924 3290 9948 3292
rect 10004 3290 10028 3292
rect 10084 3290 10090 3292
rect 9844 3238 9846 3290
rect 10026 3238 10028 3290
rect 9782 3236 9788 3238
rect 9844 3236 9868 3238
rect 9924 3236 9948 3238
rect 10004 3236 10028 3238
rect 10084 3236 10090 3238
rect 9782 3227 10090 3236
rect 10244 2774 10272 11070
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 8566 10548 10406
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9042 10732 9454
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8634 10640 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6458 10456 6598
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5914 10364 6190
rect 10428 5914 10456 6394
rect 10612 6322 10640 7686
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 5914 10732 6190
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10244 2746 10364 2774
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 10336 2446 10364 2746
rect 10796 2446 10824 10950
rect 10980 10810 11008 13359
rect 11702 13200 11758 14000
rect 12898 13200 12954 14000
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11150 11192 11562
rect 11254 11452 11562 11461
rect 11254 11450 11260 11452
rect 11316 11450 11340 11452
rect 11396 11450 11420 11452
rect 11476 11450 11500 11452
rect 11556 11450 11562 11452
rect 11316 11398 11318 11450
rect 11498 11398 11500 11450
rect 11254 11396 11260 11398
rect 11316 11396 11340 11398
rect 11396 11396 11420 11398
rect 11476 11396 11500 11398
rect 11556 11396 11562 11398
rect 11254 11387 11562 11396
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10980 9058 11008 10542
rect 11072 10470 11100 11018
rect 11348 10742 11376 11018
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11164 9178 11192 10542
rect 11254 10364 11562 10373
rect 11254 10362 11260 10364
rect 11316 10362 11340 10364
rect 11396 10362 11420 10364
rect 11476 10362 11500 10364
rect 11556 10362 11562 10364
rect 11316 10310 11318 10362
rect 11498 10310 11500 10362
rect 11254 10308 11260 10310
rect 11316 10308 11340 10310
rect 11396 10308 11420 10310
rect 11476 10308 11500 10310
rect 11556 10308 11562 10310
rect 11254 10299 11562 10308
rect 11254 9276 11562 9285
rect 11254 9274 11260 9276
rect 11316 9274 11340 9276
rect 11396 9274 11420 9276
rect 11476 9274 11500 9276
rect 11556 9274 11562 9276
rect 11316 9222 11318 9274
rect 11498 9222 11500 9274
rect 11254 9220 11260 9222
rect 11316 9220 11340 9222
rect 11396 9220 11420 9222
rect 11476 9220 11500 9222
rect 11556 9220 11562 9222
rect 11254 9211 11562 9220
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10888 9042 11008 9058
rect 10888 9036 11020 9042
rect 10888 9030 10968 9036
rect 10888 2582 10916 9030
rect 10968 8978 11020 8984
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8634 11008 8842
rect 11624 8634 11652 11222
rect 11716 11150 11744 13200
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 11354 12480 12271
rect 12912 11626 12940 13200
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12162 11248 12218 11257
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8634 11744 8774
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7886 11192 8230
rect 11254 8188 11562 8197
rect 11254 8186 11260 8188
rect 11316 8186 11340 8188
rect 11396 8186 11420 8188
rect 11476 8186 11500 8188
rect 11556 8186 11562 8188
rect 11316 8134 11318 8186
rect 11498 8134 11500 8186
rect 11254 8132 11260 8134
rect 11316 8132 11340 8134
rect 11396 8132 11420 8134
rect 11476 8132 11500 8134
rect 11556 8132 11562 8134
rect 11254 8123 11562 8132
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7342 11652 7686
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6798 11100 7142
rect 11254 7100 11562 7109
rect 11254 7098 11260 7100
rect 11316 7098 11340 7100
rect 11396 7098 11420 7100
rect 11476 7098 11500 7100
rect 11556 7098 11562 7100
rect 11316 7046 11318 7098
rect 11498 7046 11500 7098
rect 11254 7044 11260 7046
rect 11316 7044 11340 7046
rect 11396 7044 11420 7046
rect 11476 7044 11500 7046
rect 11556 7044 11562 7046
rect 11254 7035 11562 7044
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 5914 11192 6258
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11254 6012 11562 6021
rect 11254 6010 11260 6012
rect 11316 6010 11340 6012
rect 11396 6010 11420 6012
rect 11476 6010 11500 6012
rect 11556 6010 11562 6012
rect 11316 5958 11318 6010
rect 11498 5958 11500 6010
rect 11254 5956 11260 5958
rect 11316 5956 11340 5958
rect 11396 5956 11420 5958
rect 11476 5956 11500 5958
rect 11556 5956 11562 5958
rect 11254 5947 11562 5956
rect 11624 5914 11652 6190
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 4146 11100 5510
rect 11716 5234 11744 8298
rect 11808 7886 11836 10950
rect 12084 9586 12112 11222
rect 12162 11183 12218 11192
rect 12176 10674 12204 11183
rect 12726 10908 13034 10917
rect 12726 10906 12732 10908
rect 12788 10906 12812 10908
rect 12868 10906 12892 10908
rect 12948 10906 12972 10908
rect 13028 10906 13034 10908
rect 12788 10854 12790 10906
rect 12970 10854 12972 10906
rect 12726 10852 12732 10854
rect 12788 10852 12812 10854
rect 12868 10852 12892 10854
rect 12948 10852 12972 10854
rect 13028 10852 13034 10854
rect 12726 10843 13034 10852
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 9722 12296 10610
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10169 12480 10406
rect 12438 10160 12494 10169
rect 12438 10095 12494 10104
rect 12726 9820 13034 9829
rect 12726 9818 12732 9820
rect 12788 9818 12812 9820
rect 12868 9818 12892 9820
rect 12948 9818 12972 9820
rect 13028 9818 13034 9820
rect 12788 9766 12790 9818
rect 12970 9766 12972 9818
rect 12726 9764 12732 9766
rect 12788 9764 12812 9766
rect 12868 9764 12892 9766
rect 12948 9764 12972 9766
rect 13028 9764 13034 9766
rect 12726 9755 13034 9764
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11900 6882 11928 9522
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 11808 6854 11928 6882
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11254 4924 11562 4933
rect 11254 4922 11260 4924
rect 11316 4922 11340 4924
rect 11396 4922 11420 4924
rect 11476 4922 11500 4924
rect 11556 4922 11562 4924
rect 11316 4870 11318 4922
rect 11498 4870 11500 4922
rect 11254 4868 11260 4870
rect 11316 4868 11340 4870
rect 11396 4868 11420 4870
rect 11476 4868 11500 4870
rect 11556 4868 11562 4870
rect 11254 4859 11562 4868
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11808 3942 11836 6854
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11254 3836 11562 3845
rect 11254 3834 11260 3836
rect 11316 3834 11340 3836
rect 11396 3834 11420 3836
rect 11476 3834 11500 3836
rect 11556 3834 11562 3836
rect 11316 3782 11318 3834
rect 11498 3782 11500 3834
rect 11254 3780 11260 3782
rect 11316 3780 11340 3782
rect 11396 3780 11420 3782
rect 11476 3780 11500 3782
rect 11556 3780 11562 3782
rect 11254 3771 11562 3780
rect 11900 3194 11928 6734
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5914 12020 6054
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12176 5710 12204 9318
rect 12452 9081 12480 9318
rect 12438 9072 12494 9081
rect 12438 9007 12494 9016
rect 12726 8732 13034 8741
rect 12726 8730 12732 8732
rect 12788 8730 12812 8732
rect 12868 8730 12892 8732
rect 12948 8730 12972 8732
rect 13028 8730 13034 8732
rect 12788 8678 12790 8730
rect 12970 8678 12972 8730
rect 12726 8676 12732 8678
rect 12788 8676 12812 8678
rect 12868 8676 12892 8678
rect 12948 8676 12972 8678
rect 13028 8676 13034 8678
rect 12726 8667 13034 8676
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12360 7993 12388 8298
rect 12346 7984 12402 7993
rect 12346 7919 12402 7928
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 6905 12296 7686
rect 12726 7644 13034 7653
rect 12726 7642 12732 7644
rect 12788 7642 12812 7644
rect 12868 7642 12892 7644
rect 12948 7642 12972 7644
rect 13028 7642 13034 7644
rect 12788 7590 12790 7642
rect 12970 7590 12972 7642
rect 12726 7588 12732 7590
rect 12788 7588 12812 7590
rect 12868 7588 12892 7590
rect 12948 7588 12972 7590
rect 13028 7588 13034 7590
rect 12726 7579 13034 7588
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12452 7002 12480 7414
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12726 6556 13034 6565
rect 12726 6554 12732 6556
rect 12788 6554 12812 6556
rect 12868 6554 12892 6556
rect 12948 6554 12972 6556
rect 13028 6554 13034 6556
rect 12788 6502 12790 6554
rect 12970 6502 12972 6554
rect 12726 6500 12732 6502
rect 12788 6500 12812 6502
rect 12868 6500 12892 6502
rect 12948 6500 12972 6502
rect 13028 6500 13034 6502
rect 12726 6491 13034 6500
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 5914 12296 6258
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12452 5817 12480 6054
rect 12438 5808 12494 5817
rect 12438 5743 12494 5752
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11254 2748 11562 2757
rect 11254 2746 11260 2748
rect 11316 2746 11340 2748
rect 11396 2746 11420 2748
rect 11476 2746 11500 2748
rect 11556 2746 11562 2748
rect 11316 2694 11318 2746
rect 11498 2694 11500 2746
rect 11254 2692 11260 2694
rect 11316 2692 11340 2694
rect 11396 2692 11420 2694
rect 11476 2692 11500 2694
rect 11556 2692 11562 2694
rect 11254 2683 11562 2692
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10784 2440 10836 2446
rect 11992 2394 12020 5510
rect 12726 5468 13034 5477
rect 12726 5466 12732 5468
rect 12788 5466 12812 5468
rect 12868 5466 12892 5468
rect 12948 5466 12972 5468
rect 13028 5466 13034 5468
rect 12788 5414 12790 5466
rect 12970 5414 12972 5466
rect 12726 5412 12732 5414
rect 12788 5412 12812 5414
rect 12868 5412 12892 5414
rect 12948 5412 12972 5414
rect 13028 5412 13034 5414
rect 12726 5403 13034 5412
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4729 12480 4966
rect 12438 4720 12494 4729
rect 12438 4655 12494 4664
rect 12726 4380 13034 4389
rect 12726 4378 12732 4380
rect 12788 4378 12812 4380
rect 12868 4378 12892 4380
rect 12948 4378 12972 4380
rect 13028 4378 13034 4380
rect 12788 4326 12790 4378
rect 12970 4326 12972 4378
rect 12726 4324 12732 4326
rect 12788 4324 12812 4326
rect 12868 4324 12892 4326
rect 12948 4324 12972 4326
rect 13028 4324 13034 4326
rect 12726 4315 13034 4324
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3641 12480 3878
rect 12438 3632 12494 3641
rect 12438 3567 12494 3576
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12084 3194 12112 3334
rect 12360 3194 12388 3334
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12360 2553 12388 2790
rect 12346 2544 12402 2553
rect 12346 2479 12402 2488
rect 10784 2382 10836 2388
rect 11900 2378 12020 2394
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 756 2372 808 2378
rect 756 2314 808 2320
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 11888 2372 12020 2378
rect 11940 2366 12020 2372
rect 11888 2314 11940 2320
rect 768 800 796 2314
rect 2240 1170 2268 2314
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 2148 1142 2268 1170
rect 2148 800 2176 1142
rect 3528 870 3648 898
rect 3528 800 3556 870
rect 754 0 810 800
rect 2134 0 2190 800
rect 3514 0 3570 800
rect 3620 762 3648 870
rect 3804 762 3832 2246
rect 3894 2204 4202 2213
rect 3894 2202 3900 2204
rect 3956 2202 3980 2204
rect 4036 2202 4060 2204
rect 4116 2202 4140 2204
rect 4196 2202 4202 2204
rect 3956 2150 3958 2202
rect 4138 2150 4140 2202
rect 3894 2148 3900 2150
rect 3956 2148 3980 2150
rect 4036 2148 4060 2150
rect 4116 2148 4140 2150
rect 4196 2148 4202 2150
rect 3894 2139 4202 2148
rect 4908 870 5028 898
rect 4908 800 4936 870
rect 3620 734 3832 762
rect 4894 0 4950 800
rect 5000 762 5028 870
rect 5184 762 5212 2246
rect 6288 800 6316 2246
rect 6838 2204 7146 2213
rect 6838 2202 6844 2204
rect 6900 2202 6924 2204
rect 6980 2202 7004 2204
rect 7060 2202 7084 2204
rect 7140 2202 7146 2204
rect 6900 2150 6902 2202
rect 7082 2150 7084 2202
rect 6838 2148 6844 2150
rect 6900 2148 6924 2150
rect 6980 2148 7004 2150
rect 7060 2148 7084 2150
rect 7140 2148 7146 2150
rect 6838 2139 7146 2148
rect 7668 800 7696 2246
rect 9048 800 9076 2246
rect 9782 2204 10090 2213
rect 9782 2202 9788 2204
rect 9844 2202 9868 2204
rect 9924 2202 9948 2204
rect 10004 2202 10028 2204
rect 10084 2202 10090 2204
rect 9844 2150 9846 2202
rect 10026 2150 10028 2202
rect 9782 2148 9788 2150
rect 9844 2148 9868 2150
rect 9924 2148 9948 2150
rect 10004 2148 10028 2150
rect 10084 2148 10090 2150
rect 9782 2139 10090 2148
rect 10428 870 10548 898
rect 10428 800 10456 870
rect 5000 734 5212 762
rect 6274 0 6330 800
rect 7654 0 7710 800
rect 9034 0 9090 800
rect 10414 0 10470 800
rect 10520 762 10548 870
rect 10704 762 10732 2246
rect 11808 870 11928 898
rect 11808 800 11836 870
rect 10520 734 10732 762
rect 11794 0 11850 800
rect 11900 762 11928 870
rect 12084 762 12112 2246
rect 12452 1465 12480 2382
rect 12438 1456 12494 1465
rect 12438 1391 12494 1400
rect 11900 734 12112 762
rect 12636 377 12664 3334
rect 12726 3292 13034 3301
rect 12726 3290 12732 3292
rect 12788 3290 12812 3292
rect 12868 3290 12892 3292
rect 12948 3290 12972 3292
rect 13028 3290 13034 3292
rect 12788 3238 12790 3290
rect 12970 3238 12972 3290
rect 12726 3236 12732 3238
rect 12788 3236 12812 3238
rect 12868 3236 12892 3238
rect 12948 3236 12972 3238
rect 13028 3236 13034 3238
rect 12726 3227 13034 3236
rect 12726 2204 13034 2213
rect 12726 2202 12732 2204
rect 12788 2202 12812 2204
rect 12868 2202 12892 2204
rect 12948 2202 12972 2204
rect 13028 2202 13034 2204
rect 12788 2150 12790 2202
rect 12970 2150 12972 2202
rect 12726 2148 12732 2150
rect 12788 2148 12812 2150
rect 12868 2148 12892 2150
rect 12948 2148 12972 2150
rect 13028 2148 13034 2150
rect 12726 2139 13034 2148
rect 12622 368 12678 377
rect 12622 303 12678 312
<< via2 >>
rect 938 12280 994 12336
rect 10966 13368 11022 13424
rect 2428 11450 2484 11452
rect 2508 11450 2564 11452
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2428 11398 2474 11450
rect 2474 11398 2484 11450
rect 2508 11398 2538 11450
rect 2538 11398 2550 11450
rect 2550 11398 2564 11450
rect 2588 11398 2602 11450
rect 2602 11398 2614 11450
rect 2614 11398 2644 11450
rect 2668 11398 2678 11450
rect 2678 11398 2724 11450
rect 2428 11396 2484 11398
rect 2508 11396 2564 11398
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 938 10104 994 10160
rect 938 9016 994 9072
rect 1398 8200 1454 8256
rect 1858 11056 1914 11112
rect 2428 10362 2484 10364
rect 2508 10362 2564 10364
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2428 10310 2474 10362
rect 2474 10310 2484 10362
rect 2508 10310 2538 10362
rect 2538 10310 2550 10362
rect 2550 10310 2564 10362
rect 2588 10310 2602 10362
rect 2602 10310 2614 10362
rect 2614 10310 2644 10362
rect 2668 10310 2678 10362
rect 2678 10310 2724 10362
rect 2428 10308 2484 10310
rect 2508 10308 2564 10310
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2428 9274 2484 9276
rect 2508 9274 2564 9276
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2428 9222 2474 9274
rect 2474 9222 2484 9274
rect 2508 9222 2538 9274
rect 2538 9222 2550 9274
rect 2550 9222 2564 9274
rect 2588 9222 2602 9274
rect 2602 9222 2614 9274
rect 2614 9222 2644 9274
rect 2668 9222 2678 9274
rect 2678 9222 2724 9274
rect 2428 9220 2484 9222
rect 2508 9220 2564 9222
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2428 8186 2484 8188
rect 2508 8186 2564 8188
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2428 8134 2474 8186
rect 2474 8134 2484 8186
rect 2508 8134 2538 8186
rect 2538 8134 2550 8186
rect 2550 8134 2564 8186
rect 2588 8134 2602 8186
rect 2602 8134 2614 8186
rect 2614 8134 2644 8186
rect 2668 8134 2678 8186
rect 2678 8134 2724 8186
rect 2428 8132 2484 8134
rect 2508 8132 2564 8134
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 1766 6840 1822 6896
rect 2428 7098 2484 7100
rect 2508 7098 2564 7100
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2428 7046 2474 7098
rect 2474 7046 2484 7098
rect 2508 7046 2538 7098
rect 2538 7046 2550 7098
rect 2550 7046 2564 7098
rect 2588 7046 2602 7098
rect 2602 7046 2614 7098
rect 2614 7046 2644 7098
rect 2668 7046 2678 7098
rect 2678 7046 2724 7098
rect 2428 7044 2484 7046
rect 2508 7044 2564 7046
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2428 6010 2484 6012
rect 2508 6010 2564 6012
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2428 5958 2474 6010
rect 2474 5958 2484 6010
rect 2508 5958 2538 6010
rect 2538 5958 2550 6010
rect 2550 5958 2564 6010
rect 2588 5958 2602 6010
rect 2602 5958 2614 6010
rect 2614 5958 2644 6010
rect 2668 5958 2678 6010
rect 2678 5958 2724 6010
rect 2428 5956 2484 5958
rect 2508 5956 2564 5958
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 1030 5752 1086 5808
rect 2428 4922 2484 4924
rect 2508 4922 2564 4924
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2428 4870 2474 4922
rect 2474 4870 2484 4922
rect 2508 4870 2538 4922
rect 2538 4870 2550 4922
rect 2550 4870 2564 4922
rect 2588 4870 2602 4922
rect 2602 4870 2614 4922
rect 2614 4870 2644 4922
rect 2668 4870 2678 4922
rect 2678 4870 2724 4922
rect 2428 4868 2484 4870
rect 2508 4868 2564 4870
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 938 4664 994 4720
rect 2428 3834 2484 3836
rect 2508 3834 2564 3836
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2428 3782 2474 3834
rect 2474 3782 2484 3834
rect 2508 3782 2538 3834
rect 2538 3782 2550 3834
rect 2550 3782 2564 3834
rect 2588 3782 2602 3834
rect 2602 3782 2614 3834
rect 2614 3782 2644 3834
rect 2668 3782 2678 3834
rect 2678 3782 2724 3834
rect 2428 3780 2484 3782
rect 2508 3780 2564 3782
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 938 3576 994 3632
rect 2428 2746 2484 2748
rect 2508 2746 2564 2748
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2428 2694 2474 2746
rect 2474 2694 2484 2746
rect 2508 2694 2538 2746
rect 2538 2694 2550 2746
rect 2550 2694 2564 2746
rect 2588 2694 2602 2746
rect 2602 2694 2614 2746
rect 2614 2694 2644 2746
rect 2668 2694 2678 2746
rect 2678 2694 2724 2746
rect 2428 2692 2484 2694
rect 2508 2692 2564 2694
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 5372 11450 5428 11452
rect 5452 11450 5508 11452
rect 5532 11450 5588 11452
rect 5612 11450 5668 11452
rect 5372 11398 5418 11450
rect 5418 11398 5428 11450
rect 5452 11398 5482 11450
rect 5482 11398 5494 11450
rect 5494 11398 5508 11450
rect 5532 11398 5546 11450
rect 5546 11398 5558 11450
rect 5558 11398 5588 11450
rect 5612 11398 5622 11450
rect 5622 11398 5668 11450
rect 5372 11396 5428 11398
rect 5452 11396 5508 11398
rect 5532 11396 5588 11398
rect 5612 11396 5668 11398
rect 8316 11450 8372 11452
rect 8396 11450 8452 11452
rect 8476 11450 8532 11452
rect 8556 11450 8612 11452
rect 8316 11398 8362 11450
rect 8362 11398 8372 11450
rect 8396 11398 8426 11450
rect 8426 11398 8438 11450
rect 8438 11398 8452 11450
rect 8476 11398 8490 11450
rect 8490 11398 8502 11450
rect 8502 11398 8532 11450
rect 8556 11398 8566 11450
rect 8566 11398 8612 11450
rect 8316 11396 8372 11398
rect 8396 11396 8452 11398
rect 8476 11396 8532 11398
rect 8556 11396 8612 11398
rect 3900 10906 3956 10908
rect 3980 10906 4036 10908
rect 4060 10906 4116 10908
rect 4140 10906 4196 10908
rect 3900 10854 3946 10906
rect 3946 10854 3956 10906
rect 3980 10854 4010 10906
rect 4010 10854 4022 10906
rect 4022 10854 4036 10906
rect 4060 10854 4074 10906
rect 4074 10854 4086 10906
rect 4086 10854 4116 10906
rect 4140 10854 4150 10906
rect 4150 10854 4196 10906
rect 3900 10852 3956 10854
rect 3980 10852 4036 10854
rect 4060 10852 4116 10854
rect 4140 10852 4196 10854
rect 3900 9818 3956 9820
rect 3980 9818 4036 9820
rect 4060 9818 4116 9820
rect 4140 9818 4196 9820
rect 3900 9766 3946 9818
rect 3946 9766 3956 9818
rect 3980 9766 4010 9818
rect 4010 9766 4022 9818
rect 4022 9766 4036 9818
rect 4060 9766 4074 9818
rect 4074 9766 4086 9818
rect 4086 9766 4116 9818
rect 4140 9766 4150 9818
rect 4150 9766 4196 9818
rect 3900 9764 3956 9766
rect 3980 9764 4036 9766
rect 4060 9764 4116 9766
rect 4140 9764 4196 9766
rect 3900 8730 3956 8732
rect 3980 8730 4036 8732
rect 4060 8730 4116 8732
rect 4140 8730 4196 8732
rect 3900 8678 3946 8730
rect 3946 8678 3956 8730
rect 3980 8678 4010 8730
rect 4010 8678 4022 8730
rect 4022 8678 4036 8730
rect 4060 8678 4074 8730
rect 4074 8678 4086 8730
rect 4086 8678 4116 8730
rect 4140 8678 4150 8730
rect 4150 8678 4196 8730
rect 3900 8676 3956 8678
rect 3980 8676 4036 8678
rect 4060 8676 4116 8678
rect 4140 8676 4196 8678
rect 3900 7642 3956 7644
rect 3980 7642 4036 7644
rect 4060 7642 4116 7644
rect 4140 7642 4196 7644
rect 3900 7590 3946 7642
rect 3946 7590 3956 7642
rect 3980 7590 4010 7642
rect 4010 7590 4022 7642
rect 4022 7590 4036 7642
rect 4060 7590 4074 7642
rect 4074 7590 4086 7642
rect 4086 7590 4116 7642
rect 4140 7590 4150 7642
rect 4150 7590 4196 7642
rect 3900 7588 3956 7590
rect 3980 7588 4036 7590
rect 4060 7588 4116 7590
rect 4140 7588 4196 7590
rect 3900 6554 3956 6556
rect 3980 6554 4036 6556
rect 4060 6554 4116 6556
rect 4140 6554 4196 6556
rect 3900 6502 3946 6554
rect 3946 6502 3956 6554
rect 3980 6502 4010 6554
rect 4010 6502 4022 6554
rect 4022 6502 4036 6554
rect 4060 6502 4074 6554
rect 4074 6502 4086 6554
rect 4086 6502 4116 6554
rect 4140 6502 4150 6554
rect 4150 6502 4196 6554
rect 3900 6500 3956 6502
rect 3980 6500 4036 6502
rect 4060 6500 4116 6502
rect 4140 6500 4196 6502
rect 3900 5466 3956 5468
rect 3980 5466 4036 5468
rect 4060 5466 4116 5468
rect 4140 5466 4196 5468
rect 3900 5414 3946 5466
rect 3946 5414 3956 5466
rect 3980 5414 4010 5466
rect 4010 5414 4022 5466
rect 4022 5414 4036 5466
rect 4060 5414 4074 5466
rect 4074 5414 4086 5466
rect 4086 5414 4116 5466
rect 4140 5414 4150 5466
rect 4150 5414 4196 5466
rect 3900 5412 3956 5414
rect 3980 5412 4036 5414
rect 4060 5412 4116 5414
rect 4140 5412 4196 5414
rect 3900 4378 3956 4380
rect 3980 4378 4036 4380
rect 4060 4378 4116 4380
rect 4140 4378 4196 4380
rect 3900 4326 3946 4378
rect 3946 4326 3956 4378
rect 3980 4326 4010 4378
rect 4010 4326 4022 4378
rect 4022 4326 4036 4378
rect 4060 4326 4074 4378
rect 4074 4326 4086 4378
rect 4086 4326 4116 4378
rect 4140 4326 4150 4378
rect 4150 4326 4196 4378
rect 3900 4324 3956 4326
rect 3980 4324 4036 4326
rect 4060 4324 4116 4326
rect 4140 4324 4196 4326
rect 3900 3290 3956 3292
rect 3980 3290 4036 3292
rect 4060 3290 4116 3292
rect 4140 3290 4196 3292
rect 3900 3238 3946 3290
rect 3946 3238 3956 3290
rect 3980 3238 4010 3290
rect 4010 3238 4022 3290
rect 4022 3238 4036 3290
rect 4060 3238 4074 3290
rect 4074 3238 4086 3290
rect 4086 3238 4116 3290
rect 4140 3238 4150 3290
rect 4150 3238 4196 3290
rect 3900 3236 3956 3238
rect 3980 3236 4036 3238
rect 4060 3236 4116 3238
rect 4140 3236 4196 3238
rect 5372 10362 5428 10364
rect 5452 10362 5508 10364
rect 5532 10362 5588 10364
rect 5612 10362 5668 10364
rect 5372 10310 5418 10362
rect 5418 10310 5428 10362
rect 5452 10310 5482 10362
rect 5482 10310 5494 10362
rect 5494 10310 5508 10362
rect 5532 10310 5546 10362
rect 5546 10310 5558 10362
rect 5558 10310 5588 10362
rect 5612 10310 5622 10362
rect 5622 10310 5668 10362
rect 5372 10308 5428 10310
rect 5452 10308 5508 10310
rect 5532 10308 5588 10310
rect 5612 10308 5668 10310
rect 5372 9274 5428 9276
rect 5452 9274 5508 9276
rect 5532 9274 5588 9276
rect 5612 9274 5668 9276
rect 5372 9222 5418 9274
rect 5418 9222 5428 9274
rect 5452 9222 5482 9274
rect 5482 9222 5494 9274
rect 5494 9222 5508 9274
rect 5532 9222 5546 9274
rect 5546 9222 5558 9274
rect 5558 9222 5588 9274
rect 5612 9222 5622 9274
rect 5622 9222 5668 9274
rect 5372 9220 5428 9222
rect 5452 9220 5508 9222
rect 5532 9220 5588 9222
rect 5612 9220 5668 9222
rect 5372 8186 5428 8188
rect 5452 8186 5508 8188
rect 5532 8186 5588 8188
rect 5612 8186 5668 8188
rect 5372 8134 5418 8186
rect 5418 8134 5428 8186
rect 5452 8134 5482 8186
rect 5482 8134 5494 8186
rect 5494 8134 5508 8186
rect 5532 8134 5546 8186
rect 5546 8134 5558 8186
rect 5558 8134 5588 8186
rect 5612 8134 5622 8186
rect 5622 8134 5668 8186
rect 5372 8132 5428 8134
rect 5452 8132 5508 8134
rect 5532 8132 5588 8134
rect 5612 8132 5668 8134
rect 5372 7098 5428 7100
rect 5452 7098 5508 7100
rect 5532 7098 5588 7100
rect 5612 7098 5668 7100
rect 5372 7046 5418 7098
rect 5418 7046 5428 7098
rect 5452 7046 5482 7098
rect 5482 7046 5494 7098
rect 5494 7046 5508 7098
rect 5532 7046 5546 7098
rect 5546 7046 5558 7098
rect 5558 7046 5588 7098
rect 5612 7046 5622 7098
rect 5622 7046 5668 7098
rect 5372 7044 5428 7046
rect 5452 7044 5508 7046
rect 5532 7044 5588 7046
rect 5612 7044 5668 7046
rect 5372 6010 5428 6012
rect 5452 6010 5508 6012
rect 5532 6010 5588 6012
rect 5612 6010 5668 6012
rect 5372 5958 5418 6010
rect 5418 5958 5428 6010
rect 5452 5958 5482 6010
rect 5482 5958 5494 6010
rect 5494 5958 5508 6010
rect 5532 5958 5546 6010
rect 5546 5958 5558 6010
rect 5558 5958 5588 6010
rect 5612 5958 5622 6010
rect 5622 5958 5668 6010
rect 5372 5956 5428 5958
rect 5452 5956 5508 5958
rect 5532 5956 5588 5958
rect 5612 5956 5668 5958
rect 5372 4922 5428 4924
rect 5452 4922 5508 4924
rect 5532 4922 5588 4924
rect 5612 4922 5668 4924
rect 5372 4870 5418 4922
rect 5418 4870 5428 4922
rect 5452 4870 5482 4922
rect 5482 4870 5494 4922
rect 5494 4870 5508 4922
rect 5532 4870 5546 4922
rect 5546 4870 5558 4922
rect 5558 4870 5588 4922
rect 5612 4870 5622 4922
rect 5622 4870 5668 4922
rect 5372 4868 5428 4870
rect 5452 4868 5508 4870
rect 5532 4868 5588 4870
rect 5612 4868 5668 4870
rect 5372 3834 5428 3836
rect 5452 3834 5508 3836
rect 5532 3834 5588 3836
rect 5612 3834 5668 3836
rect 5372 3782 5418 3834
rect 5418 3782 5428 3834
rect 5452 3782 5482 3834
rect 5482 3782 5494 3834
rect 5494 3782 5508 3834
rect 5532 3782 5546 3834
rect 5546 3782 5558 3834
rect 5558 3782 5588 3834
rect 5612 3782 5622 3834
rect 5622 3782 5668 3834
rect 5372 3780 5428 3782
rect 5452 3780 5508 3782
rect 5532 3780 5588 3782
rect 5612 3780 5668 3782
rect 6844 10906 6900 10908
rect 6924 10906 6980 10908
rect 7004 10906 7060 10908
rect 7084 10906 7140 10908
rect 6844 10854 6890 10906
rect 6890 10854 6900 10906
rect 6924 10854 6954 10906
rect 6954 10854 6966 10906
rect 6966 10854 6980 10906
rect 7004 10854 7018 10906
rect 7018 10854 7030 10906
rect 7030 10854 7060 10906
rect 7084 10854 7094 10906
rect 7094 10854 7140 10906
rect 6844 10852 6900 10854
rect 6924 10852 6980 10854
rect 7004 10852 7060 10854
rect 7084 10852 7140 10854
rect 6844 9818 6900 9820
rect 6924 9818 6980 9820
rect 7004 9818 7060 9820
rect 7084 9818 7140 9820
rect 6844 9766 6890 9818
rect 6890 9766 6900 9818
rect 6924 9766 6954 9818
rect 6954 9766 6966 9818
rect 6966 9766 6980 9818
rect 7004 9766 7018 9818
rect 7018 9766 7030 9818
rect 7030 9766 7060 9818
rect 7084 9766 7094 9818
rect 7094 9766 7140 9818
rect 6844 9764 6900 9766
rect 6924 9764 6980 9766
rect 7004 9764 7060 9766
rect 7084 9764 7140 9766
rect 6844 8730 6900 8732
rect 6924 8730 6980 8732
rect 7004 8730 7060 8732
rect 7084 8730 7140 8732
rect 6844 8678 6890 8730
rect 6890 8678 6900 8730
rect 6924 8678 6954 8730
rect 6954 8678 6966 8730
rect 6966 8678 6980 8730
rect 7004 8678 7018 8730
rect 7018 8678 7030 8730
rect 7030 8678 7060 8730
rect 7084 8678 7094 8730
rect 7094 8678 7140 8730
rect 6844 8676 6900 8678
rect 6924 8676 6980 8678
rect 7004 8676 7060 8678
rect 7084 8676 7140 8678
rect 5372 2746 5428 2748
rect 5452 2746 5508 2748
rect 5532 2746 5588 2748
rect 5612 2746 5668 2748
rect 3422 2488 3478 2544
rect 5372 2694 5418 2746
rect 5418 2694 5428 2746
rect 5452 2694 5482 2746
rect 5482 2694 5494 2746
rect 5494 2694 5508 2746
rect 5532 2694 5546 2746
rect 5546 2694 5558 2746
rect 5558 2694 5588 2746
rect 5612 2694 5622 2746
rect 5622 2694 5668 2746
rect 5372 2692 5428 2694
rect 5452 2692 5508 2694
rect 5532 2692 5588 2694
rect 5612 2692 5668 2694
rect 6844 7642 6900 7644
rect 6924 7642 6980 7644
rect 7004 7642 7060 7644
rect 7084 7642 7140 7644
rect 6844 7590 6890 7642
rect 6890 7590 6900 7642
rect 6924 7590 6954 7642
rect 6954 7590 6966 7642
rect 6966 7590 6980 7642
rect 7004 7590 7018 7642
rect 7018 7590 7030 7642
rect 7030 7590 7060 7642
rect 7084 7590 7094 7642
rect 7094 7590 7140 7642
rect 6844 7588 6900 7590
rect 6924 7588 6980 7590
rect 7004 7588 7060 7590
rect 7084 7588 7140 7590
rect 8316 10362 8372 10364
rect 8396 10362 8452 10364
rect 8476 10362 8532 10364
rect 8556 10362 8612 10364
rect 8316 10310 8362 10362
rect 8362 10310 8372 10362
rect 8396 10310 8426 10362
rect 8426 10310 8438 10362
rect 8438 10310 8452 10362
rect 8476 10310 8490 10362
rect 8490 10310 8502 10362
rect 8502 10310 8532 10362
rect 8556 10310 8566 10362
rect 8566 10310 8612 10362
rect 8316 10308 8372 10310
rect 8396 10308 8452 10310
rect 8476 10308 8532 10310
rect 8556 10308 8612 10310
rect 8316 9274 8372 9276
rect 8396 9274 8452 9276
rect 8476 9274 8532 9276
rect 8556 9274 8612 9276
rect 8316 9222 8362 9274
rect 8362 9222 8372 9274
rect 8396 9222 8426 9274
rect 8426 9222 8438 9274
rect 8438 9222 8452 9274
rect 8476 9222 8490 9274
rect 8490 9222 8502 9274
rect 8502 9222 8532 9274
rect 8556 9222 8566 9274
rect 8566 9222 8612 9274
rect 8316 9220 8372 9222
rect 8396 9220 8452 9222
rect 8476 9220 8532 9222
rect 8556 9220 8612 9222
rect 6844 6554 6900 6556
rect 6924 6554 6980 6556
rect 7004 6554 7060 6556
rect 7084 6554 7140 6556
rect 6844 6502 6890 6554
rect 6890 6502 6900 6554
rect 6924 6502 6954 6554
rect 6954 6502 6966 6554
rect 6966 6502 6980 6554
rect 7004 6502 7018 6554
rect 7018 6502 7030 6554
rect 7030 6502 7060 6554
rect 7084 6502 7094 6554
rect 7094 6502 7140 6554
rect 6844 6500 6900 6502
rect 6924 6500 6980 6502
rect 7004 6500 7060 6502
rect 7084 6500 7140 6502
rect 6844 5466 6900 5468
rect 6924 5466 6980 5468
rect 7004 5466 7060 5468
rect 7084 5466 7140 5468
rect 6844 5414 6890 5466
rect 6890 5414 6900 5466
rect 6924 5414 6954 5466
rect 6954 5414 6966 5466
rect 6966 5414 6980 5466
rect 7004 5414 7018 5466
rect 7018 5414 7030 5466
rect 7030 5414 7060 5466
rect 7084 5414 7094 5466
rect 7094 5414 7140 5466
rect 6844 5412 6900 5414
rect 6924 5412 6980 5414
rect 7004 5412 7060 5414
rect 7084 5412 7140 5414
rect 6844 4378 6900 4380
rect 6924 4378 6980 4380
rect 7004 4378 7060 4380
rect 7084 4378 7140 4380
rect 6844 4326 6890 4378
rect 6890 4326 6900 4378
rect 6924 4326 6954 4378
rect 6954 4326 6966 4378
rect 6966 4326 6980 4378
rect 7004 4326 7018 4378
rect 7018 4326 7030 4378
rect 7030 4326 7060 4378
rect 7084 4326 7094 4378
rect 7094 4326 7140 4378
rect 6844 4324 6900 4326
rect 6924 4324 6980 4326
rect 7004 4324 7060 4326
rect 7084 4324 7140 4326
rect 6844 3290 6900 3292
rect 6924 3290 6980 3292
rect 7004 3290 7060 3292
rect 7084 3290 7140 3292
rect 6844 3238 6890 3290
rect 6890 3238 6900 3290
rect 6924 3238 6954 3290
rect 6954 3238 6966 3290
rect 6966 3238 6980 3290
rect 7004 3238 7018 3290
rect 7018 3238 7030 3290
rect 7030 3238 7060 3290
rect 7084 3238 7094 3290
rect 7094 3238 7140 3290
rect 6844 3236 6900 3238
rect 6924 3236 6980 3238
rect 7004 3236 7060 3238
rect 7084 3236 7140 3238
rect 8316 8186 8372 8188
rect 8396 8186 8452 8188
rect 8476 8186 8532 8188
rect 8556 8186 8612 8188
rect 8316 8134 8362 8186
rect 8362 8134 8372 8186
rect 8396 8134 8426 8186
rect 8426 8134 8438 8186
rect 8438 8134 8452 8186
rect 8476 8134 8490 8186
rect 8490 8134 8502 8186
rect 8502 8134 8532 8186
rect 8556 8134 8566 8186
rect 8566 8134 8612 8186
rect 8316 8132 8372 8134
rect 8396 8132 8452 8134
rect 8476 8132 8532 8134
rect 8556 8132 8612 8134
rect 8316 7098 8372 7100
rect 8396 7098 8452 7100
rect 8476 7098 8532 7100
rect 8556 7098 8612 7100
rect 8316 7046 8362 7098
rect 8362 7046 8372 7098
rect 8396 7046 8426 7098
rect 8426 7046 8438 7098
rect 8438 7046 8452 7098
rect 8476 7046 8490 7098
rect 8490 7046 8502 7098
rect 8502 7046 8532 7098
rect 8556 7046 8566 7098
rect 8566 7046 8612 7098
rect 8316 7044 8372 7046
rect 8396 7044 8452 7046
rect 8476 7044 8532 7046
rect 8556 7044 8612 7046
rect 8316 6010 8372 6012
rect 8396 6010 8452 6012
rect 8476 6010 8532 6012
rect 8556 6010 8612 6012
rect 8316 5958 8362 6010
rect 8362 5958 8372 6010
rect 8396 5958 8426 6010
rect 8426 5958 8438 6010
rect 8438 5958 8452 6010
rect 8476 5958 8490 6010
rect 8490 5958 8502 6010
rect 8502 5958 8532 6010
rect 8556 5958 8566 6010
rect 8566 5958 8612 6010
rect 8316 5956 8372 5958
rect 8396 5956 8452 5958
rect 8476 5956 8532 5958
rect 8556 5956 8612 5958
rect 8316 4922 8372 4924
rect 8396 4922 8452 4924
rect 8476 4922 8532 4924
rect 8556 4922 8612 4924
rect 8316 4870 8362 4922
rect 8362 4870 8372 4922
rect 8396 4870 8426 4922
rect 8426 4870 8438 4922
rect 8438 4870 8452 4922
rect 8476 4870 8490 4922
rect 8490 4870 8502 4922
rect 8502 4870 8532 4922
rect 8556 4870 8566 4922
rect 8566 4870 8612 4922
rect 8316 4868 8372 4870
rect 8396 4868 8452 4870
rect 8476 4868 8532 4870
rect 8556 4868 8612 4870
rect 8316 3834 8372 3836
rect 8396 3834 8452 3836
rect 8476 3834 8532 3836
rect 8556 3834 8612 3836
rect 8316 3782 8362 3834
rect 8362 3782 8372 3834
rect 8396 3782 8426 3834
rect 8426 3782 8438 3834
rect 8438 3782 8452 3834
rect 8476 3782 8490 3834
rect 8490 3782 8502 3834
rect 8502 3782 8532 3834
rect 8556 3782 8566 3834
rect 8566 3782 8612 3834
rect 8316 3780 8372 3782
rect 8396 3780 8452 3782
rect 8476 3780 8532 3782
rect 8556 3780 8612 3782
rect 8316 2746 8372 2748
rect 8396 2746 8452 2748
rect 8476 2746 8532 2748
rect 8556 2746 8612 2748
rect 8316 2694 8362 2746
rect 8362 2694 8372 2746
rect 8396 2694 8426 2746
rect 8426 2694 8438 2746
rect 8438 2694 8452 2746
rect 8476 2694 8490 2746
rect 8490 2694 8502 2746
rect 8502 2694 8532 2746
rect 8556 2694 8566 2746
rect 8566 2694 8612 2746
rect 8316 2692 8372 2694
rect 8396 2692 8452 2694
rect 8476 2692 8532 2694
rect 8556 2692 8612 2694
rect 9788 10906 9844 10908
rect 9868 10906 9924 10908
rect 9948 10906 10004 10908
rect 10028 10906 10084 10908
rect 9788 10854 9834 10906
rect 9834 10854 9844 10906
rect 9868 10854 9898 10906
rect 9898 10854 9910 10906
rect 9910 10854 9924 10906
rect 9948 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 10004 10906
rect 10028 10854 10038 10906
rect 10038 10854 10084 10906
rect 9788 10852 9844 10854
rect 9868 10852 9924 10854
rect 9948 10852 10004 10854
rect 10028 10852 10084 10854
rect 9788 9818 9844 9820
rect 9868 9818 9924 9820
rect 9948 9818 10004 9820
rect 10028 9818 10084 9820
rect 9788 9766 9834 9818
rect 9834 9766 9844 9818
rect 9868 9766 9898 9818
rect 9898 9766 9910 9818
rect 9910 9766 9924 9818
rect 9948 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 10004 9818
rect 10028 9766 10038 9818
rect 10038 9766 10084 9818
rect 9788 9764 9844 9766
rect 9868 9764 9924 9766
rect 9948 9764 10004 9766
rect 10028 9764 10084 9766
rect 9788 8730 9844 8732
rect 9868 8730 9924 8732
rect 9948 8730 10004 8732
rect 10028 8730 10084 8732
rect 9788 8678 9834 8730
rect 9834 8678 9844 8730
rect 9868 8678 9898 8730
rect 9898 8678 9910 8730
rect 9910 8678 9924 8730
rect 9948 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 10004 8730
rect 10028 8678 10038 8730
rect 10038 8678 10084 8730
rect 9788 8676 9844 8678
rect 9868 8676 9924 8678
rect 9948 8676 10004 8678
rect 10028 8676 10084 8678
rect 9788 7642 9844 7644
rect 9868 7642 9924 7644
rect 9948 7642 10004 7644
rect 10028 7642 10084 7644
rect 9788 7590 9834 7642
rect 9834 7590 9844 7642
rect 9868 7590 9898 7642
rect 9898 7590 9910 7642
rect 9910 7590 9924 7642
rect 9948 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 10004 7642
rect 10028 7590 10038 7642
rect 10038 7590 10084 7642
rect 9788 7588 9844 7590
rect 9868 7588 9924 7590
rect 9948 7588 10004 7590
rect 10028 7588 10084 7590
rect 9788 6554 9844 6556
rect 9868 6554 9924 6556
rect 9948 6554 10004 6556
rect 10028 6554 10084 6556
rect 9788 6502 9834 6554
rect 9834 6502 9844 6554
rect 9868 6502 9898 6554
rect 9898 6502 9910 6554
rect 9910 6502 9924 6554
rect 9948 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 10004 6554
rect 10028 6502 10038 6554
rect 10038 6502 10084 6554
rect 9788 6500 9844 6502
rect 9868 6500 9924 6502
rect 9948 6500 10004 6502
rect 10028 6500 10084 6502
rect 9788 5466 9844 5468
rect 9868 5466 9924 5468
rect 9948 5466 10004 5468
rect 10028 5466 10084 5468
rect 9788 5414 9834 5466
rect 9834 5414 9844 5466
rect 9868 5414 9898 5466
rect 9898 5414 9910 5466
rect 9910 5414 9924 5466
rect 9948 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 10004 5466
rect 10028 5414 10038 5466
rect 10038 5414 10084 5466
rect 9788 5412 9844 5414
rect 9868 5412 9924 5414
rect 9948 5412 10004 5414
rect 10028 5412 10084 5414
rect 9788 4378 9844 4380
rect 9868 4378 9924 4380
rect 9948 4378 10004 4380
rect 10028 4378 10084 4380
rect 9788 4326 9834 4378
rect 9834 4326 9844 4378
rect 9868 4326 9898 4378
rect 9898 4326 9910 4378
rect 9910 4326 9924 4378
rect 9948 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 10004 4378
rect 10028 4326 10038 4378
rect 10038 4326 10084 4378
rect 9788 4324 9844 4326
rect 9868 4324 9924 4326
rect 9948 4324 10004 4326
rect 10028 4324 10084 4326
rect 9788 3290 9844 3292
rect 9868 3290 9924 3292
rect 9948 3290 10004 3292
rect 10028 3290 10084 3292
rect 9788 3238 9834 3290
rect 9834 3238 9844 3290
rect 9868 3238 9898 3290
rect 9898 3238 9910 3290
rect 9910 3238 9924 3290
rect 9948 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 10004 3290
rect 10028 3238 10038 3290
rect 10038 3238 10084 3290
rect 9788 3236 9844 3238
rect 9868 3236 9924 3238
rect 9948 3236 10004 3238
rect 10028 3236 10084 3238
rect 11260 11450 11316 11452
rect 11340 11450 11396 11452
rect 11420 11450 11476 11452
rect 11500 11450 11556 11452
rect 11260 11398 11306 11450
rect 11306 11398 11316 11450
rect 11340 11398 11370 11450
rect 11370 11398 11382 11450
rect 11382 11398 11396 11450
rect 11420 11398 11434 11450
rect 11434 11398 11446 11450
rect 11446 11398 11476 11450
rect 11500 11398 11510 11450
rect 11510 11398 11556 11450
rect 11260 11396 11316 11398
rect 11340 11396 11396 11398
rect 11420 11396 11476 11398
rect 11500 11396 11556 11398
rect 11260 10362 11316 10364
rect 11340 10362 11396 10364
rect 11420 10362 11476 10364
rect 11500 10362 11556 10364
rect 11260 10310 11306 10362
rect 11306 10310 11316 10362
rect 11340 10310 11370 10362
rect 11370 10310 11382 10362
rect 11382 10310 11396 10362
rect 11420 10310 11434 10362
rect 11434 10310 11446 10362
rect 11446 10310 11476 10362
rect 11500 10310 11510 10362
rect 11510 10310 11556 10362
rect 11260 10308 11316 10310
rect 11340 10308 11396 10310
rect 11420 10308 11476 10310
rect 11500 10308 11556 10310
rect 11260 9274 11316 9276
rect 11340 9274 11396 9276
rect 11420 9274 11476 9276
rect 11500 9274 11556 9276
rect 11260 9222 11306 9274
rect 11306 9222 11316 9274
rect 11340 9222 11370 9274
rect 11370 9222 11382 9274
rect 11382 9222 11396 9274
rect 11420 9222 11434 9274
rect 11434 9222 11446 9274
rect 11446 9222 11476 9274
rect 11500 9222 11510 9274
rect 11510 9222 11556 9274
rect 11260 9220 11316 9222
rect 11340 9220 11396 9222
rect 11420 9220 11476 9222
rect 11500 9220 11556 9222
rect 12438 12280 12494 12336
rect 11260 8186 11316 8188
rect 11340 8186 11396 8188
rect 11420 8186 11476 8188
rect 11500 8186 11556 8188
rect 11260 8134 11306 8186
rect 11306 8134 11316 8186
rect 11340 8134 11370 8186
rect 11370 8134 11382 8186
rect 11382 8134 11396 8186
rect 11420 8134 11434 8186
rect 11434 8134 11446 8186
rect 11446 8134 11476 8186
rect 11500 8134 11510 8186
rect 11510 8134 11556 8186
rect 11260 8132 11316 8134
rect 11340 8132 11396 8134
rect 11420 8132 11476 8134
rect 11500 8132 11556 8134
rect 11260 7098 11316 7100
rect 11340 7098 11396 7100
rect 11420 7098 11476 7100
rect 11500 7098 11556 7100
rect 11260 7046 11306 7098
rect 11306 7046 11316 7098
rect 11340 7046 11370 7098
rect 11370 7046 11382 7098
rect 11382 7046 11396 7098
rect 11420 7046 11434 7098
rect 11434 7046 11446 7098
rect 11446 7046 11476 7098
rect 11500 7046 11510 7098
rect 11510 7046 11556 7098
rect 11260 7044 11316 7046
rect 11340 7044 11396 7046
rect 11420 7044 11476 7046
rect 11500 7044 11556 7046
rect 11260 6010 11316 6012
rect 11340 6010 11396 6012
rect 11420 6010 11476 6012
rect 11500 6010 11556 6012
rect 11260 5958 11306 6010
rect 11306 5958 11316 6010
rect 11340 5958 11370 6010
rect 11370 5958 11382 6010
rect 11382 5958 11396 6010
rect 11420 5958 11434 6010
rect 11434 5958 11446 6010
rect 11446 5958 11476 6010
rect 11500 5958 11510 6010
rect 11510 5958 11556 6010
rect 11260 5956 11316 5958
rect 11340 5956 11396 5958
rect 11420 5956 11476 5958
rect 11500 5956 11556 5958
rect 12162 11192 12218 11248
rect 12732 10906 12788 10908
rect 12812 10906 12868 10908
rect 12892 10906 12948 10908
rect 12972 10906 13028 10908
rect 12732 10854 12778 10906
rect 12778 10854 12788 10906
rect 12812 10854 12842 10906
rect 12842 10854 12854 10906
rect 12854 10854 12868 10906
rect 12892 10854 12906 10906
rect 12906 10854 12918 10906
rect 12918 10854 12948 10906
rect 12972 10854 12982 10906
rect 12982 10854 13028 10906
rect 12732 10852 12788 10854
rect 12812 10852 12868 10854
rect 12892 10852 12948 10854
rect 12972 10852 13028 10854
rect 12438 10104 12494 10160
rect 12732 9818 12788 9820
rect 12812 9818 12868 9820
rect 12892 9818 12948 9820
rect 12972 9818 13028 9820
rect 12732 9766 12778 9818
rect 12778 9766 12788 9818
rect 12812 9766 12842 9818
rect 12842 9766 12854 9818
rect 12854 9766 12868 9818
rect 12892 9766 12906 9818
rect 12906 9766 12918 9818
rect 12918 9766 12948 9818
rect 12972 9766 12982 9818
rect 12982 9766 13028 9818
rect 12732 9764 12788 9766
rect 12812 9764 12868 9766
rect 12892 9764 12948 9766
rect 12972 9764 13028 9766
rect 11260 4922 11316 4924
rect 11340 4922 11396 4924
rect 11420 4922 11476 4924
rect 11500 4922 11556 4924
rect 11260 4870 11306 4922
rect 11306 4870 11316 4922
rect 11340 4870 11370 4922
rect 11370 4870 11382 4922
rect 11382 4870 11396 4922
rect 11420 4870 11434 4922
rect 11434 4870 11446 4922
rect 11446 4870 11476 4922
rect 11500 4870 11510 4922
rect 11510 4870 11556 4922
rect 11260 4868 11316 4870
rect 11340 4868 11396 4870
rect 11420 4868 11476 4870
rect 11500 4868 11556 4870
rect 11260 3834 11316 3836
rect 11340 3834 11396 3836
rect 11420 3834 11476 3836
rect 11500 3834 11556 3836
rect 11260 3782 11306 3834
rect 11306 3782 11316 3834
rect 11340 3782 11370 3834
rect 11370 3782 11382 3834
rect 11382 3782 11396 3834
rect 11420 3782 11434 3834
rect 11434 3782 11446 3834
rect 11446 3782 11476 3834
rect 11500 3782 11510 3834
rect 11510 3782 11556 3834
rect 11260 3780 11316 3782
rect 11340 3780 11396 3782
rect 11420 3780 11476 3782
rect 11500 3780 11556 3782
rect 12438 9016 12494 9072
rect 12732 8730 12788 8732
rect 12812 8730 12868 8732
rect 12892 8730 12948 8732
rect 12972 8730 13028 8732
rect 12732 8678 12778 8730
rect 12778 8678 12788 8730
rect 12812 8678 12842 8730
rect 12842 8678 12854 8730
rect 12854 8678 12868 8730
rect 12892 8678 12906 8730
rect 12906 8678 12918 8730
rect 12918 8678 12948 8730
rect 12972 8678 12982 8730
rect 12982 8678 13028 8730
rect 12732 8676 12788 8678
rect 12812 8676 12868 8678
rect 12892 8676 12948 8678
rect 12972 8676 13028 8678
rect 12346 7928 12402 7984
rect 12732 7642 12788 7644
rect 12812 7642 12868 7644
rect 12892 7642 12948 7644
rect 12972 7642 13028 7644
rect 12732 7590 12778 7642
rect 12778 7590 12788 7642
rect 12812 7590 12842 7642
rect 12842 7590 12854 7642
rect 12854 7590 12868 7642
rect 12892 7590 12906 7642
rect 12906 7590 12918 7642
rect 12918 7590 12948 7642
rect 12972 7590 12982 7642
rect 12982 7590 13028 7642
rect 12732 7588 12788 7590
rect 12812 7588 12868 7590
rect 12892 7588 12948 7590
rect 12972 7588 13028 7590
rect 12254 6840 12310 6896
rect 12732 6554 12788 6556
rect 12812 6554 12868 6556
rect 12892 6554 12948 6556
rect 12972 6554 13028 6556
rect 12732 6502 12778 6554
rect 12778 6502 12788 6554
rect 12812 6502 12842 6554
rect 12842 6502 12854 6554
rect 12854 6502 12868 6554
rect 12892 6502 12906 6554
rect 12906 6502 12918 6554
rect 12918 6502 12948 6554
rect 12972 6502 12982 6554
rect 12982 6502 13028 6554
rect 12732 6500 12788 6502
rect 12812 6500 12868 6502
rect 12892 6500 12948 6502
rect 12972 6500 13028 6502
rect 12438 5752 12494 5808
rect 11260 2746 11316 2748
rect 11340 2746 11396 2748
rect 11420 2746 11476 2748
rect 11500 2746 11556 2748
rect 11260 2694 11306 2746
rect 11306 2694 11316 2746
rect 11340 2694 11370 2746
rect 11370 2694 11382 2746
rect 11382 2694 11396 2746
rect 11420 2694 11434 2746
rect 11434 2694 11446 2746
rect 11446 2694 11476 2746
rect 11500 2694 11510 2746
rect 11510 2694 11556 2746
rect 11260 2692 11316 2694
rect 11340 2692 11396 2694
rect 11420 2692 11476 2694
rect 11500 2692 11556 2694
rect 12732 5466 12788 5468
rect 12812 5466 12868 5468
rect 12892 5466 12948 5468
rect 12972 5466 13028 5468
rect 12732 5414 12778 5466
rect 12778 5414 12788 5466
rect 12812 5414 12842 5466
rect 12842 5414 12854 5466
rect 12854 5414 12868 5466
rect 12892 5414 12906 5466
rect 12906 5414 12918 5466
rect 12918 5414 12948 5466
rect 12972 5414 12982 5466
rect 12982 5414 13028 5466
rect 12732 5412 12788 5414
rect 12812 5412 12868 5414
rect 12892 5412 12948 5414
rect 12972 5412 13028 5414
rect 12438 4664 12494 4720
rect 12732 4378 12788 4380
rect 12812 4378 12868 4380
rect 12892 4378 12948 4380
rect 12972 4378 13028 4380
rect 12732 4326 12778 4378
rect 12778 4326 12788 4378
rect 12812 4326 12842 4378
rect 12842 4326 12854 4378
rect 12854 4326 12868 4378
rect 12892 4326 12906 4378
rect 12906 4326 12918 4378
rect 12918 4326 12948 4378
rect 12972 4326 12982 4378
rect 12982 4326 13028 4378
rect 12732 4324 12788 4326
rect 12812 4324 12868 4326
rect 12892 4324 12948 4326
rect 12972 4324 13028 4326
rect 12438 3576 12494 3632
rect 12346 2488 12402 2544
rect 3900 2202 3956 2204
rect 3980 2202 4036 2204
rect 4060 2202 4116 2204
rect 4140 2202 4196 2204
rect 3900 2150 3946 2202
rect 3946 2150 3956 2202
rect 3980 2150 4010 2202
rect 4010 2150 4022 2202
rect 4022 2150 4036 2202
rect 4060 2150 4074 2202
rect 4074 2150 4086 2202
rect 4086 2150 4116 2202
rect 4140 2150 4150 2202
rect 4150 2150 4196 2202
rect 3900 2148 3956 2150
rect 3980 2148 4036 2150
rect 4060 2148 4116 2150
rect 4140 2148 4196 2150
rect 6844 2202 6900 2204
rect 6924 2202 6980 2204
rect 7004 2202 7060 2204
rect 7084 2202 7140 2204
rect 6844 2150 6890 2202
rect 6890 2150 6900 2202
rect 6924 2150 6954 2202
rect 6954 2150 6966 2202
rect 6966 2150 6980 2202
rect 7004 2150 7018 2202
rect 7018 2150 7030 2202
rect 7030 2150 7060 2202
rect 7084 2150 7094 2202
rect 7094 2150 7140 2202
rect 6844 2148 6900 2150
rect 6924 2148 6980 2150
rect 7004 2148 7060 2150
rect 7084 2148 7140 2150
rect 9788 2202 9844 2204
rect 9868 2202 9924 2204
rect 9948 2202 10004 2204
rect 10028 2202 10084 2204
rect 9788 2150 9834 2202
rect 9834 2150 9844 2202
rect 9868 2150 9898 2202
rect 9898 2150 9910 2202
rect 9910 2150 9924 2202
rect 9948 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 10004 2202
rect 10028 2150 10038 2202
rect 10038 2150 10084 2202
rect 9788 2148 9844 2150
rect 9868 2148 9924 2150
rect 9948 2148 10004 2150
rect 10028 2148 10084 2150
rect 12438 1400 12494 1456
rect 12732 3290 12788 3292
rect 12812 3290 12868 3292
rect 12892 3290 12948 3292
rect 12972 3290 13028 3292
rect 12732 3238 12778 3290
rect 12778 3238 12788 3290
rect 12812 3238 12842 3290
rect 12842 3238 12854 3290
rect 12854 3238 12868 3290
rect 12892 3238 12906 3290
rect 12906 3238 12918 3290
rect 12918 3238 12948 3290
rect 12972 3238 12982 3290
rect 12982 3238 13028 3290
rect 12732 3236 12788 3238
rect 12812 3236 12868 3238
rect 12892 3236 12948 3238
rect 12972 3236 13028 3238
rect 12732 2202 12788 2204
rect 12812 2202 12868 2204
rect 12892 2202 12948 2204
rect 12972 2202 13028 2204
rect 12732 2150 12778 2202
rect 12778 2150 12788 2202
rect 12812 2150 12842 2202
rect 12842 2150 12854 2202
rect 12854 2150 12868 2202
rect 12892 2150 12906 2202
rect 12906 2150 12918 2202
rect 12918 2150 12948 2202
rect 12972 2150 12982 2202
rect 12982 2150 13028 2202
rect 12732 2148 12788 2150
rect 12812 2148 12868 2150
rect 12892 2148 12948 2150
rect 12972 2148 13028 2150
rect 12622 312 12678 368
<< metal3 >>
rect 10961 13426 11027 13429
rect 13200 13426 14000 13456
rect 10961 13424 14000 13426
rect 10961 13368 10966 13424
rect 11022 13368 14000 13424
rect 10961 13366 14000 13368
rect 10961 13363 11027 13366
rect 13200 13336 14000 13366
rect 0 12338 800 12368
rect 933 12338 999 12341
rect 0 12336 999 12338
rect 0 12280 938 12336
rect 994 12280 999 12336
rect 0 12278 999 12280
rect 0 12248 800 12278
rect 933 12275 999 12278
rect 12433 12338 12499 12341
rect 13200 12338 14000 12368
rect 12433 12336 14000 12338
rect 12433 12280 12438 12336
rect 12494 12280 14000 12336
rect 12433 12278 14000 12280
rect 12433 12275 12499 12278
rect 13200 12248 14000 12278
rect 2418 11456 2734 11457
rect 2418 11392 2424 11456
rect 2488 11392 2504 11456
rect 2568 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2734 11456
rect 2418 11391 2734 11392
rect 5362 11456 5678 11457
rect 5362 11392 5368 11456
rect 5432 11392 5448 11456
rect 5512 11392 5528 11456
rect 5592 11392 5608 11456
rect 5672 11392 5678 11456
rect 5362 11391 5678 11392
rect 8306 11456 8622 11457
rect 8306 11392 8312 11456
rect 8376 11392 8392 11456
rect 8456 11392 8472 11456
rect 8536 11392 8552 11456
rect 8616 11392 8622 11456
rect 8306 11391 8622 11392
rect 11250 11456 11566 11457
rect 11250 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11566 11456
rect 11250 11391 11566 11392
rect 0 11250 800 11280
rect 12157 11250 12223 11253
rect 13200 11250 14000 11280
rect 0 11190 1042 11250
rect 0 11160 800 11190
rect 982 11114 1042 11190
rect 12157 11248 14000 11250
rect 12157 11192 12162 11248
rect 12218 11192 14000 11248
rect 12157 11190 14000 11192
rect 12157 11187 12223 11190
rect 13200 11160 14000 11190
rect 1853 11114 1919 11117
rect 982 11112 1919 11114
rect 982 11056 1858 11112
rect 1914 11056 1919 11112
rect 982 11054 1919 11056
rect 1853 11051 1919 11054
rect 3890 10912 4206 10913
rect 3890 10848 3896 10912
rect 3960 10848 3976 10912
rect 4040 10848 4056 10912
rect 4120 10848 4136 10912
rect 4200 10848 4206 10912
rect 3890 10847 4206 10848
rect 6834 10912 7150 10913
rect 6834 10848 6840 10912
rect 6904 10848 6920 10912
rect 6984 10848 7000 10912
rect 7064 10848 7080 10912
rect 7144 10848 7150 10912
rect 6834 10847 7150 10848
rect 9778 10912 10094 10913
rect 9778 10848 9784 10912
rect 9848 10848 9864 10912
rect 9928 10848 9944 10912
rect 10008 10848 10024 10912
rect 10088 10848 10094 10912
rect 9778 10847 10094 10848
rect 12722 10912 13038 10913
rect 12722 10848 12728 10912
rect 12792 10848 12808 10912
rect 12872 10848 12888 10912
rect 12952 10848 12968 10912
rect 13032 10848 13038 10912
rect 12722 10847 13038 10848
rect 2418 10368 2734 10369
rect 2418 10304 2424 10368
rect 2488 10304 2504 10368
rect 2568 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2734 10368
rect 2418 10303 2734 10304
rect 5362 10368 5678 10369
rect 5362 10304 5368 10368
rect 5432 10304 5448 10368
rect 5512 10304 5528 10368
rect 5592 10304 5608 10368
rect 5672 10304 5678 10368
rect 5362 10303 5678 10304
rect 8306 10368 8622 10369
rect 8306 10304 8312 10368
rect 8376 10304 8392 10368
rect 8456 10304 8472 10368
rect 8536 10304 8552 10368
rect 8616 10304 8622 10368
rect 8306 10303 8622 10304
rect 11250 10368 11566 10369
rect 11250 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11566 10368
rect 11250 10303 11566 10304
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 12433 10162 12499 10165
rect 13200 10162 14000 10192
rect 12433 10160 14000 10162
rect 12433 10104 12438 10160
rect 12494 10104 14000 10160
rect 12433 10102 14000 10104
rect 12433 10099 12499 10102
rect 13200 10072 14000 10102
rect 3890 9824 4206 9825
rect 3890 9760 3896 9824
rect 3960 9760 3976 9824
rect 4040 9760 4056 9824
rect 4120 9760 4136 9824
rect 4200 9760 4206 9824
rect 3890 9759 4206 9760
rect 6834 9824 7150 9825
rect 6834 9760 6840 9824
rect 6904 9760 6920 9824
rect 6984 9760 7000 9824
rect 7064 9760 7080 9824
rect 7144 9760 7150 9824
rect 6834 9759 7150 9760
rect 9778 9824 10094 9825
rect 9778 9760 9784 9824
rect 9848 9760 9864 9824
rect 9928 9760 9944 9824
rect 10008 9760 10024 9824
rect 10088 9760 10094 9824
rect 9778 9759 10094 9760
rect 12722 9824 13038 9825
rect 12722 9760 12728 9824
rect 12792 9760 12808 9824
rect 12872 9760 12888 9824
rect 12952 9760 12968 9824
rect 13032 9760 13038 9824
rect 12722 9759 13038 9760
rect 2418 9280 2734 9281
rect 2418 9216 2424 9280
rect 2488 9216 2504 9280
rect 2568 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2734 9280
rect 2418 9215 2734 9216
rect 5362 9280 5678 9281
rect 5362 9216 5368 9280
rect 5432 9216 5448 9280
rect 5512 9216 5528 9280
rect 5592 9216 5608 9280
rect 5672 9216 5678 9280
rect 5362 9215 5678 9216
rect 8306 9280 8622 9281
rect 8306 9216 8312 9280
rect 8376 9216 8392 9280
rect 8456 9216 8472 9280
rect 8536 9216 8552 9280
rect 8616 9216 8622 9280
rect 8306 9215 8622 9216
rect 11250 9280 11566 9281
rect 11250 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11566 9280
rect 11250 9215 11566 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 12433 9074 12499 9077
rect 13200 9074 14000 9104
rect 12433 9072 14000 9074
rect 12433 9016 12438 9072
rect 12494 9016 14000 9072
rect 12433 9014 14000 9016
rect 12433 9011 12499 9014
rect 13200 8984 14000 9014
rect 3890 8736 4206 8737
rect 3890 8672 3896 8736
rect 3960 8672 3976 8736
rect 4040 8672 4056 8736
rect 4120 8672 4136 8736
rect 4200 8672 4206 8736
rect 3890 8671 4206 8672
rect 6834 8736 7150 8737
rect 6834 8672 6840 8736
rect 6904 8672 6920 8736
rect 6984 8672 7000 8736
rect 7064 8672 7080 8736
rect 7144 8672 7150 8736
rect 6834 8671 7150 8672
rect 9778 8736 10094 8737
rect 9778 8672 9784 8736
rect 9848 8672 9864 8736
rect 9928 8672 9944 8736
rect 10008 8672 10024 8736
rect 10088 8672 10094 8736
rect 9778 8671 10094 8672
rect 12722 8736 13038 8737
rect 12722 8672 12728 8736
rect 12792 8672 12808 8736
rect 12872 8672 12888 8736
rect 12952 8672 12968 8736
rect 13032 8672 13038 8736
rect 12722 8671 13038 8672
rect 1393 8258 1459 8261
rect 798 8256 1459 8258
rect 798 8200 1398 8256
rect 1454 8200 1459 8256
rect 798 8198 1459 8200
rect 798 8016 858 8198
rect 1393 8195 1459 8198
rect 2418 8192 2734 8193
rect 2418 8128 2424 8192
rect 2488 8128 2504 8192
rect 2568 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2734 8192
rect 2418 8127 2734 8128
rect 5362 8192 5678 8193
rect 5362 8128 5368 8192
rect 5432 8128 5448 8192
rect 5512 8128 5528 8192
rect 5592 8128 5608 8192
rect 5672 8128 5678 8192
rect 5362 8127 5678 8128
rect 8306 8192 8622 8193
rect 8306 8128 8312 8192
rect 8376 8128 8392 8192
rect 8456 8128 8472 8192
rect 8536 8128 8552 8192
rect 8616 8128 8622 8192
rect 8306 8127 8622 8128
rect 11250 8192 11566 8193
rect 11250 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11566 8192
rect 11250 8127 11566 8128
rect 0 7926 858 8016
rect 12341 7986 12407 7989
rect 13200 7986 14000 8016
rect 12341 7984 14000 7986
rect 12341 7928 12346 7984
rect 12402 7928 14000 7984
rect 12341 7926 14000 7928
rect 0 7896 800 7926
rect 12341 7923 12407 7926
rect 13200 7896 14000 7926
rect 3890 7648 4206 7649
rect 3890 7584 3896 7648
rect 3960 7584 3976 7648
rect 4040 7584 4056 7648
rect 4120 7584 4136 7648
rect 4200 7584 4206 7648
rect 3890 7583 4206 7584
rect 6834 7648 7150 7649
rect 6834 7584 6840 7648
rect 6904 7584 6920 7648
rect 6984 7584 7000 7648
rect 7064 7584 7080 7648
rect 7144 7584 7150 7648
rect 6834 7583 7150 7584
rect 9778 7648 10094 7649
rect 9778 7584 9784 7648
rect 9848 7584 9864 7648
rect 9928 7584 9944 7648
rect 10008 7584 10024 7648
rect 10088 7584 10094 7648
rect 9778 7583 10094 7584
rect 12722 7648 13038 7649
rect 12722 7584 12728 7648
rect 12792 7584 12808 7648
rect 12872 7584 12888 7648
rect 12952 7584 12968 7648
rect 13032 7584 13038 7648
rect 12722 7583 13038 7584
rect 2418 7104 2734 7105
rect 2418 7040 2424 7104
rect 2488 7040 2504 7104
rect 2568 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2734 7104
rect 2418 7039 2734 7040
rect 5362 7104 5678 7105
rect 5362 7040 5368 7104
rect 5432 7040 5448 7104
rect 5512 7040 5528 7104
rect 5592 7040 5608 7104
rect 5672 7040 5678 7104
rect 5362 7039 5678 7040
rect 8306 7104 8622 7105
rect 8306 7040 8312 7104
rect 8376 7040 8392 7104
rect 8456 7040 8472 7104
rect 8536 7040 8552 7104
rect 8616 7040 8622 7104
rect 8306 7039 8622 7040
rect 11250 7104 11566 7105
rect 11250 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11566 7104
rect 11250 7039 11566 7040
rect 0 6898 800 6928
rect 1761 6898 1827 6901
rect 0 6896 1827 6898
rect 0 6840 1766 6896
rect 1822 6840 1827 6896
rect 0 6838 1827 6840
rect 0 6808 800 6838
rect 1761 6835 1827 6838
rect 12249 6898 12315 6901
rect 13200 6898 14000 6928
rect 12249 6896 14000 6898
rect 12249 6840 12254 6896
rect 12310 6840 14000 6896
rect 12249 6838 14000 6840
rect 12249 6835 12315 6838
rect 13200 6808 14000 6838
rect 3890 6560 4206 6561
rect 3890 6496 3896 6560
rect 3960 6496 3976 6560
rect 4040 6496 4056 6560
rect 4120 6496 4136 6560
rect 4200 6496 4206 6560
rect 3890 6495 4206 6496
rect 6834 6560 7150 6561
rect 6834 6496 6840 6560
rect 6904 6496 6920 6560
rect 6984 6496 7000 6560
rect 7064 6496 7080 6560
rect 7144 6496 7150 6560
rect 6834 6495 7150 6496
rect 9778 6560 10094 6561
rect 9778 6496 9784 6560
rect 9848 6496 9864 6560
rect 9928 6496 9944 6560
rect 10008 6496 10024 6560
rect 10088 6496 10094 6560
rect 9778 6495 10094 6496
rect 12722 6560 13038 6561
rect 12722 6496 12728 6560
rect 12792 6496 12808 6560
rect 12872 6496 12888 6560
rect 12952 6496 12968 6560
rect 13032 6496 13038 6560
rect 12722 6495 13038 6496
rect 2418 6016 2734 6017
rect 2418 5952 2424 6016
rect 2488 5952 2504 6016
rect 2568 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2734 6016
rect 2418 5951 2734 5952
rect 5362 6016 5678 6017
rect 5362 5952 5368 6016
rect 5432 5952 5448 6016
rect 5512 5952 5528 6016
rect 5592 5952 5608 6016
rect 5672 5952 5678 6016
rect 5362 5951 5678 5952
rect 8306 6016 8622 6017
rect 8306 5952 8312 6016
rect 8376 5952 8392 6016
rect 8456 5952 8472 6016
rect 8536 5952 8552 6016
rect 8616 5952 8622 6016
rect 8306 5951 8622 5952
rect 11250 6016 11566 6017
rect 11250 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11566 6016
rect 11250 5951 11566 5952
rect 0 5810 800 5840
rect 1025 5810 1091 5813
rect 0 5808 1091 5810
rect 0 5752 1030 5808
rect 1086 5752 1091 5808
rect 0 5750 1091 5752
rect 0 5720 800 5750
rect 1025 5747 1091 5750
rect 12433 5810 12499 5813
rect 13200 5810 14000 5840
rect 12433 5808 14000 5810
rect 12433 5752 12438 5808
rect 12494 5752 14000 5808
rect 12433 5750 14000 5752
rect 12433 5747 12499 5750
rect 13200 5720 14000 5750
rect 3890 5472 4206 5473
rect 3890 5408 3896 5472
rect 3960 5408 3976 5472
rect 4040 5408 4056 5472
rect 4120 5408 4136 5472
rect 4200 5408 4206 5472
rect 3890 5407 4206 5408
rect 6834 5472 7150 5473
rect 6834 5408 6840 5472
rect 6904 5408 6920 5472
rect 6984 5408 7000 5472
rect 7064 5408 7080 5472
rect 7144 5408 7150 5472
rect 6834 5407 7150 5408
rect 9778 5472 10094 5473
rect 9778 5408 9784 5472
rect 9848 5408 9864 5472
rect 9928 5408 9944 5472
rect 10008 5408 10024 5472
rect 10088 5408 10094 5472
rect 9778 5407 10094 5408
rect 12722 5472 13038 5473
rect 12722 5408 12728 5472
rect 12792 5408 12808 5472
rect 12872 5408 12888 5472
rect 12952 5408 12968 5472
rect 13032 5408 13038 5472
rect 12722 5407 13038 5408
rect 2418 4928 2734 4929
rect 2418 4864 2424 4928
rect 2488 4864 2504 4928
rect 2568 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2734 4928
rect 2418 4863 2734 4864
rect 5362 4928 5678 4929
rect 5362 4864 5368 4928
rect 5432 4864 5448 4928
rect 5512 4864 5528 4928
rect 5592 4864 5608 4928
rect 5672 4864 5678 4928
rect 5362 4863 5678 4864
rect 8306 4928 8622 4929
rect 8306 4864 8312 4928
rect 8376 4864 8392 4928
rect 8456 4864 8472 4928
rect 8536 4864 8552 4928
rect 8616 4864 8622 4928
rect 8306 4863 8622 4864
rect 11250 4928 11566 4929
rect 11250 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11566 4928
rect 11250 4863 11566 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 12433 4722 12499 4725
rect 13200 4722 14000 4752
rect 12433 4720 14000 4722
rect 12433 4664 12438 4720
rect 12494 4664 14000 4720
rect 12433 4662 14000 4664
rect 12433 4659 12499 4662
rect 13200 4632 14000 4662
rect 3890 4384 4206 4385
rect 3890 4320 3896 4384
rect 3960 4320 3976 4384
rect 4040 4320 4056 4384
rect 4120 4320 4136 4384
rect 4200 4320 4206 4384
rect 3890 4319 4206 4320
rect 6834 4384 7150 4385
rect 6834 4320 6840 4384
rect 6904 4320 6920 4384
rect 6984 4320 7000 4384
rect 7064 4320 7080 4384
rect 7144 4320 7150 4384
rect 6834 4319 7150 4320
rect 9778 4384 10094 4385
rect 9778 4320 9784 4384
rect 9848 4320 9864 4384
rect 9928 4320 9944 4384
rect 10008 4320 10024 4384
rect 10088 4320 10094 4384
rect 9778 4319 10094 4320
rect 12722 4384 13038 4385
rect 12722 4320 12728 4384
rect 12792 4320 12808 4384
rect 12872 4320 12888 4384
rect 12952 4320 12968 4384
rect 13032 4320 13038 4384
rect 12722 4319 13038 4320
rect 2418 3840 2734 3841
rect 2418 3776 2424 3840
rect 2488 3776 2504 3840
rect 2568 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2734 3840
rect 2418 3775 2734 3776
rect 5362 3840 5678 3841
rect 5362 3776 5368 3840
rect 5432 3776 5448 3840
rect 5512 3776 5528 3840
rect 5592 3776 5608 3840
rect 5672 3776 5678 3840
rect 5362 3775 5678 3776
rect 8306 3840 8622 3841
rect 8306 3776 8312 3840
rect 8376 3776 8392 3840
rect 8456 3776 8472 3840
rect 8536 3776 8552 3840
rect 8616 3776 8622 3840
rect 8306 3775 8622 3776
rect 11250 3840 11566 3841
rect 11250 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11566 3840
rect 11250 3775 11566 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 12433 3634 12499 3637
rect 13200 3634 14000 3664
rect 12433 3632 14000 3634
rect 12433 3576 12438 3632
rect 12494 3576 14000 3632
rect 12433 3574 14000 3576
rect 12433 3571 12499 3574
rect 13200 3544 14000 3574
rect 3890 3296 4206 3297
rect 3890 3232 3896 3296
rect 3960 3232 3976 3296
rect 4040 3232 4056 3296
rect 4120 3232 4136 3296
rect 4200 3232 4206 3296
rect 3890 3231 4206 3232
rect 6834 3296 7150 3297
rect 6834 3232 6840 3296
rect 6904 3232 6920 3296
rect 6984 3232 7000 3296
rect 7064 3232 7080 3296
rect 7144 3232 7150 3296
rect 6834 3231 7150 3232
rect 9778 3296 10094 3297
rect 9778 3232 9784 3296
rect 9848 3232 9864 3296
rect 9928 3232 9944 3296
rect 10008 3232 10024 3296
rect 10088 3232 10094 3296
rect 9778 3231 10094 3232
rect 12722 3296 13038 3297
rect 12722 3232 12728 3296
rect 12792 3232 12808 3296
rect 12872 3232 12888 3296
rect 12952 3232 12968 3296
rect 13032 3232 13038 3296
rect 12722 3231 13038 3232
rect 2418 2752 2734 2753
rect 2418 2688 2424 2752
rect 2488 2688 2504 2752
rect 2568 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2734 2752
rect 2418 2687 2734 2688
rect 5362 2752 5678 2753
rect 5362 2688 5368 2752
rect 5432 2688 5448 2752
rect 5512 2688 5528 2752
rect 5592 2688 5608 2752
rect 5672 2688 5678 2752
rect 5362 2687 5678 2688
rect 8306 2752 8622 2753
rect 8306 2688 8312 2752
rect 8376 2688 8392 2752
rect 8456 2688 8472 2752
rect 8536 2688 8552 2752
rect 8616 2688 8622 2752
rect 8306 2687 8622 2688
rect 11250 2752 11566 2753
rect 11250 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11566 2752
rect 11250 2687 11566 2688
rect 0 2546 800 2576
rect 3417 2546 3483 2549
rect 0 2544 3483 2546
rect 0 2488 3422 2544
rect 3478 2488 3483 2544
rect 0 2486 3483 2488
rect 0 2456 800 2486
rect 3417 2483 3483 2486
rect 12341 2546 12407 2549
rect 13200 2546 14000 2576
rect 12341 2544 14000 2546
rect 12341 2488 12346 2544
rect 12402 2488 14000 2544
rect 12341 2486 14000 2488
rect 12341 2483 12407 2486
rect 13200 2456 14000 2486
rect 3890 2208 4206 2209
rect 3890 2144 3896 2208
rect 3960 2144 3976 2208
rect 4040 2144 4056 2208
rect 4120 2144 4136 2208
rect 4200 2144 4206 2208
rect 3890 2143 4206 2144
rect 6834 2208 7150 2209
rect 6834 2144 6840 2208
rect 6904 2144 6920 2208
rect 6984 2144 7000 2208
rect 7064 2144 7080 2208
rect 7144 2144 7150 2208
rect 6834 2143 7150 2144
rect 9778 2208 10094 2209
rect 9778 2144 9784 2208
rect 9848 2144 9864 2208
rect 9928 2144 9944 2208
rect 10008 2144 10024 2208
rect 10088 2144 10094 2208
rect 9778 2143 10094 2144
rect 12722 2208 13038 2209
rect 12722 2144 12728 2208
rect 12792 2144 12808 2208
rect 12872 2144 12888 2208
rect 12952 2144 12968 2208
rect 13032 2144 13038 2208
rect 12722 2143 13038 2144
rect 12433 1458 12499 1461
rect 13200 1458 14000 1488
rect 12433 1456 14000 1458
rect 12433 1400 12438 1456
rect 12494 1400 14000 1456
rect 12433 1398 14000 1400
rect 12433 1395 12499 1398
rect 13200 1368 14000 1398
rect 12617 370 12683 373
rect 13200 370 14000 400
rect 12617 368 14000 370
rect 12617 312 12622 368
rect 12678 312 14000 368
rect 12617 310 14000 312
rect 12617 307 12683 310
rect 13200 280 14000 310
<< via3 >>
rect 2424 11452 2488 11456
rect 2424 11396 2428 11452
rect 2428 11396 2484 11452
rect 2484 11396 2488 11452
rect 2424 11392 2488 11396
rect 2504 11452 2568 11456
rect 2504 11396 2508 11452
rect 2508 11396 2564 11452
rect 2564 11396 2568 11452
rect 2504 11392 2568 11396
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 5368 11452 5432 11456
rect 5368 11396 5372 11452
rect 5372 11396 5428 11452
rect 5428 11396 5432 11452
rect 5368 11392 5432 11396
rect 5448 11452 5512 11456
rect 5448 11396 5452 11452
rect 5452 11396 5508 11452
rect 5508 11396 5512 11452
rect 5448 11392 5512 11396
rect 5528 11452 5592 11456
rect 5528 11396 5532 11452
rect 5532 11396 5588 11452
rect 5588 11396 5592 11452
rect 5528 11392 5592 11396
rect 5608 11452 5672 11456
rect 5608 11396 5612 11452
rect 5612 11396 5668 11452
rect 5668 11396 5672 11452
rect 5608 11392 5672 11396
rect 8312 11452 8376 11456
rect 8312 11396 8316 11452
rect 8316 11396 8372 11452
rect 8372 11396 8376 11452
rect 8312 11392 8376 11396
rect 8392 11452 8456 11456
rect 8392 11396 8396 11452
rect 8396 11396 8452 11452
rect 8452 11396 8456 11452
rect 8392 11392 8456 11396
rect 8472 11452 8536 11456
rect 8472 11396 8476 11452
rect 8476 11396 8532 11452
rect 8532 11396 8536 11452
rect 8472 11392 8536 11396
rect 8552 11452 8616 11456
rect 8552 11396 8556 11452
rect 8556 11396 8612 11452
rect 8612 11396 8616 11452
rect 8552 11392 8616 11396
rect 11256 11452 11320 11456
rect 11256 11396 11260 11452
rect 11260 11396 11316 11452
rect 11316 11396 11320 11452
rect 11256 11392 11320 11396
rect 11336 11452 11400 11456
rect 11336 11396 11340 11452
rect 11340 11396 11396 11452
rect 11396 11396 11400 11452
rect 11336 11392 11400 11396
rect 11416 11452 11480 11456
rect 11416 11396 11420 11452
rect 11420 11396 11476 11452
rect 11476 11396 11480 11452
rect 11416 11392 11480 11396
rect 11496 11452 11560 11456
rect 11496 11396 11500 11452
rect 11500 11396 11556 11452
rect 11556 11396 11560 11452
rect 11496 11392 11560 11396
rect 3896 10908 3960 10912
rect 3896 10852 3900 10908
rect 3900 10852 3956 10908
rect 3956 10852 3960 10908
rect 3896 10848 3960 10852
rect 3976 10908 4040 10912
rect 3976 10852 3980 10908
rect 3980 10852 4036 10908
rect 4036 10852 4040 10908
rect 3976 10848 4040 10852
rect 4056 10908 4120 10912
rect 4056 10852 4060 10908
rect 4060 10852 4116 10908
rect 4116 10852 4120 10908
rect 4056 10848 4120 10852
rect 4136 10908 4200 10912
rect 4136 10852 4140 10908
rect 4140 10852 4196 10908
rect 4196 10852 4200 10908
rect 4136 10848 4200 10852
rect 6840 10908 6904 10912
rect 6840 10852 6844 10908
rect 6844 10852 6900 10908
rect 6900 10852 6904 10908
rect 6840 10848 6904 10852
rect 6920 10908 6984 10912
rect 6920 10852 6924 10908
rect 6924 10852 6980 10908
rect 6980 10852 6984 10908
rect 6920 10848 6984 10852
rect 7000 10908 7064 10912
rect 7000 10852 7004 10908
rect 7004 10852 7060 10908
rect 7060 10852 7064 10908
rect 7000 10848 7064 10852
rect 7080 10908 7144 10912
rect 7080 10852 7084 10908
rect 7084 10852 7140 10908
rect 7140 10852 7144 10908
rect 7080 10848 7144 10852
rect 9784 10908 9848 10912
rect 9784 10852 9788 10908
rect 9788 10852 9844 10908
rect 9844 10852 9848 10908
rect 9784 10848 9848 10852
rect 9864 10908 9928 10912
rect 9864 10852 9868 10908
rect 9868 10852 9924 10908
rect 9924 10852 9928 10908
rect 9864 10848 9928 10852
rect 9944 10908 10008 10912
rect 9944 10852 9948 10908
rect 9948 10852 10004 10908
rect 10004 10852 10008 10908
rect 9944 10848 10008 10852
rect 10024 10908 10088 10912
rect 10024 10852 10028 10908
rect 10028 10852 10084 10908
rect 10084 10852 10088 10908
rect 10024 10848 10088 10852
rect 12728 10908 12792 10912
rect 12728 10852 12732 10908
rect 12732 10852 12788 10908
rect 12788 10852 12792 10908
rect 12728 10848 12792 10852
rect 12808 10908 12872 10912
rect 12808 10852 12812 10908
rect 12812 10852 12868 10908
rect 12868 10852 12872 10908
rect 12808 10848 12872 10852
rect 12888 10908 12952 10912
rect 12888 10852 12892 10908
rect 12892 10852 12948 10908
rect 12948 10852 12952 10908
rect 12888 10848 12952 10852
rect 12968 10908 13032 10912
rect 12968 10852 12972 10908
rect 12972 10852 13028 10908
rect 13028 10852 13032 10908
rect 12968 10848 13032 10852
rect 2424 10364 2488 10368
rect 2424 10308 2428 10364
rect 2428 10308 2484 10364
rect 2484 10308 2488 10364
rect 2424 10304 2488 10308
rect 2504 10364 2568 10368
rect 2504 10308 2508 10364
rect 2508 10308 2564 10364
rect 2564 10308 2568 10364
rect 2504 10304 2568 10308
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 5368 10364 5432 10368
rect 5368 10308 5372 10364
rect 5372 10308 5428 10364
rect 5428 10308 5432 10364
rect 5368 10304 5432 10308
rect 5448 10364 5512 10368
rect 5448 10308 5452 10364
rect 5452 10308 5508 10364
rect 5508 10308 5512 10364
rect 5448 10304 5512 10308
rect 5528 10364 5592 10368
rect 5528 10308 5532 10364
rect 5532 10308 5588 10364
rect 5588 10308 5592 10364
rect 5528 10304 5592 10308
rect 5608 10364 5672 10368
rect 5608 10308 5612 10364
rect 5612 10308 5668 10364
rect 5668 10308 5672 10364
rect 5608 10304 5672 10308
rect 8312 10364 8376 10368
rect 8312 10308 8316 10364
rect 8316 10308 8372 10364
rect 8372 10308 8376 10364
rect 8312 10304 8376 10308
rect 8392 10364 8456 10368
rect 8392 10308 8396 10364
rect 8396 10308 8452 10364
rect 8452 10308 8456 10364
rect 8392 10304 8456 10308
rect 8472 10364 8536 10368
rect 8472 10308 8476 10364
rect 8476 10308 8532 10364
rect 8532 10308 8536 10364
rect 8472 10304 8536 10308
rect 8552 10364 8616 10368
rect 8552 10308 8556 10364
rect 8556 10308 8612 10364
rect 8612 10308 8616 10364
rect 8552 10304 8616 10308
rect 11256 10364 11320 10368
rect 11256 10308 11260 10364
rect 11260 10308 11316 10364
rect 11316 10308 11320 10364
rect 11256 10304 11320 10308
rect 11336 10364 11400 10368
rect 11336 10308 11340 10364
rect 11340 10308 11396 10364
rect 11396 10308 11400 10364
rect 11336 10304 11400 10308
rect 11416 10364 11480 10368
rect 11416 10308 11420 10364
rect 11420 10308 11476 10364
rect 11476 10308 11480 10364
rect 11416 10304 11480 10308
rect 11496 10364 11560 10368
rect 11496 10308 11500 10364
rect 11500 10308 11556 10364
rect 11556 10308 11560 10364
rect 11496 10304 11560 10308
rect 3896 9820 3960 9824
rect 3896 9764 3900 9820
rect 3900 9764 3956 9820
rect 3956 9764 3960 9820
rect 3896 9760 3960 9764
rect 3976 9820 4040 9824
rect 3976 9764 3980 9820
rect 3980 9764 4036 9820
rect 4036 9764 4040 9820
rect 3976 9760 4040 9764
rect 4056 9820 4120 9824
rect 4056 9764 4060 9820
rect 4060 9764 4116 9820
rect 4116 9764 4120 9820
rect 4056 9760 4120 9764
rect 4136 9820 4200 9824
rect 4136 9764 4140 9820
rect 4140 9764 4196 9820
rect 4196 9764 4200 9820
rect 4136 9760 4200 9764
rect 6840 9820 6904 9824
rect 6840 9764 6844 9820
rect 6844 9764 6900 9820
rect 6900 9764 6904 9820
rect 6840 9760 6904 9764
rect 6920 9820 6984 9824
rect 6920 9764 6924 9820
rect 6924 9764 6980 9820
rect 6980 9764 6984 9820
rect 6920 9760 6984 9764
rect 7000 9820 7064 9824
rect 7000 9764 7004 9820
rect 7004 9764 7060 9820
rect 7060 9764 7064 9820
rect 7000 9760 7064 9764
rect 7080 9820 7144 9824
rect 7080 9764 7084 9820
rect 7084 9764 7140 9820
rect 7140 9764 7144 9820
rect 7080 9760 7144 9764
rect 9784 9820 9848 9824
rect 9784 9764 9788 9820
rect 9788 9764 9844 9820
rect 9844 9764 9848 9820
rect 9784 9760 9848 9764
rect 9864 9820 9928 9824
rect 9864 9764 9868 9820
rect 9868 9764 9924 9820
rect 9924 9764 9928 9820
rect 9864 9760 9928 9764
rect 9944 9820 10008 9824
rect 9944 9764 9948 9820
rect 9948 9764 10004 9820
rect 10004 9764 10008 9820
rect 9944 9760 10008 9764
rect 10024 9820 10088 9824
rect 10024 9764 10028 9820
rect 10028 9764 10084 9820
rect 10084 9764 10088 9820
rect 10024 9760 10088 9764
rect 12728 9820 12792 9824
rect 12728 9764 12732 9820
rect 12732 9764 12788 9820
rect 12788 9764 12792 9820
rect 12728 9760 12792 9764
rect 12808 9820 12872 9824
rect 12808 9764 12812 9820
rect 12812 9764 12868 9820
rect 12868 9764 12872 9820
rect 12808 9760 12872 9764
rect 12888 9820 12952 9824
rect 12888 9764 12892 9820
rect 12892 9764 12948 9820
rect 12948 9764 12952 9820
rect 12888 9760 12952 9764
rect 12968 9820 13032 9824
rect 12968 9764 12972 9820
rect 12972 9764 13028 9820
rect 13028 9764 13032 9820
rect 12968 9760 13032 9764
rect 2424 9276 2488 9280
rect 2424 9220 2428 9276
rect 2428 9220 2484 9276
rect 2484 9220 2488 9276
rect 2424 9216 2488 9220
rect 2504 9276 2568 9280
rect 2504 9220 2508 9276
rect 2508 9220 2564 9276
rect 2564 9220 2568 9276
rect 2504 9216 2568 9220
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 5368 9276 5432 9280
rect 5368 9220 5372 9276
rect 5372 9220 5428 9276
rect 5428 9220 5432 9276
rect 5368 9216 5432 9220
rect 5448 9276 5512 9280
rect 5448 9220 5452 9276
rect 5452 9220 5508 9276
rect 5508 9220 5512 9276
rect 5448 9216 5512 9220
rect 5528 9276 5592 9280
rect 5528 9220 5532 9276
rect 5532 9220 5588 9276
rect 5588 9220 5592 9276
rect 5528 9216 5592 9220
rect 5608 9276 5672 9280
rect 5608 9220 5612 9276
rect 5612 9220 5668 9276
rect 5668 9220 5672 9276
rect 5608 9216 5672 9220
rect 8312 9276 8376 9280
rect 8312 9220 8316 9276
rect 8316 9220 8372 9276
rect 8372 9220 8376 9276
rect 8312 9216 8376 9220
rect 8392 9276 8456 9280
rect 8392 9220 8396 9276
rect 8396 9220 8452 9276
rect 8452 9220 8456 9276
rect 8392 9216 8456 9220
rect 8472 9276 8536 9280
rect 8472 9220 8476 9276
rect 8476 9220 8532 9276
rect 8532 9220 8536 9276
rect 8472 9216 8536 9220
rect 8552 9276 8616 9280
rect 8552 9220 8556 9276
rect 8556 9220 8612 9276
rect 8612 9220 8616 9276
rect 8552 9216 8616 9220
rect 11256 9276 11320 9280
rect 11256 9220 11260 9276
rect 11260 9220 11316 9276
rect 11316 9220 11320 9276
rect 11256 9216 11320 9220
rect 11336 9276 11400 9280
rect 11336 9220 11340 9276
rect 11340 9220 11396 9276
rect 11396 9220 11400 9276
rect 11336 9216 11400 9220
rect 11416 9276 11480 9280
rect 11416 9220 11420 9276
rect 11420 9220 11476 9276
rect 11476 9220 11480 9276
rect 11416 9216 11480 9220
rect 11496 9276 11560 9280
rect 11496 9220 11500 9276
rect 11500 9220 11556 9276
rect 11556 9220 11560 9276
rect 11496 9216 11560 9220
rect 3896 8732 3960 8736
rect 3896 8676 3900 8732
rect 3900 8676 3956 8732
rect 3956 8676 3960 8732
rect 3896 8672 3960 8676
rect 3976 8732 4040 8736
rect 3976 8676 3980 8732
rect 3980 8676 4036 8732
rect 4036 8676 4040 8732
rect 3976 8672 4040 8676
rect 4056 8732 4120 8736
rect 4056 8676 4060 8732
rect 4060 8676 4116 8732
rect 4116 8676 4120 8732
rect 4056 8672 4120 8676
rect 4136 8732 4200 8736
rect 4136 8676 4140 8732
rect 4140 8676 4196 8732
rect 4196 8676 4200 8732
rect 4136 8672 4200 8676
rect 6840 8732 6904 8736
rect 6840 8676 6844 8732
rect 6844 8676 6900 8732
rect 6900 8676 6904 8732
rect 6840 8672 6904 8676
rect 6920 8732 6984 8736
rect 6920 8676 6924 8732
rect 6924 8676 6980 8732
rect 6980 8676 6984 8732
rect 6920 8672 6984 8676
rect 7000 8732 7064 8736
rect 7000 8676 7004 8732
rect 7004 8676 7060 8732
rect 7060 8676 7064 8732
rect 7000 8672 7064 8676
rect 7080 8732 7144 8736
rect 7080 8676 7084 8732
rect 7084 8676 7140 8732
rect 7140 8676 7144 8732
rect 7080 8672 7144 8676
rect 9784 8732 9848 8736
rect 9784 8676 9788 8732
rect 9788 8676 9844 8732
rect 9844 8676 9848 8732
rect 9784 8672 9848 8676
rect 9864 8732 9928 8736
rect 9864 8676 9868 8732
rect 9868 8676 9924 8732
rect 9924 8676 9928 8732
rect 9864 8672 9928 8676
rect 9944 8732 10008 8736
rect 9944 8676 9948 8732
rect 9948 8676 10004 8732
rect 10004 8676 10008 8732
rect 9944 8672 10008 8676
rect 10024 8732 10088 8736
rect 10024 8676 10028 8732
rect 10028 8676 10084 8732
rect 10084 8676 10088 8732
rect 10024 8672 10088 8676
rect 12728 8732 12792 8736
rect 12728 8676 12732 8732
rect 12732 8676 12788 8732
rect 12788 8676 12792 8732
rect 12728 8672 12792 8676
rect 12808 8732 12872 8736
rect 12808 8676 12812 8732
rect 12812 8676 12868 8732
rect 12868 8676 12872 8732
rect 12808 8672 12872 8676
rect 12888 8732 12952 8736
rect 12888 8676 12892 8732
rect 12892 8676 12948 8732
rect 12948 8676 12952 8732
rect 12888 8672 12952 8676
rect 12968 8732 13032 8736
rect 12968 8676 12972 8732
rect 12972 8676 13028 8732
rect 13028 8676 13032 8732
rect 12968 8672 13032 8676
rect 2424 8188 2488 8192
rect 2424 8132 2428 8188
rect 2428 8132 2484 8188
rect 2484 8132 2488 8188
rect 2424 8128 2488 8132
rect 2504 8188 2568 8192
rect 2504 8132 2508 8188
rect 2508 8132 2564 8188
rect 2564 8132 2568 8188
rect 2504 8128 2568 8132
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 5368 8188 5432 8192
rect 5368 8132 5372 8188
rect 5372 8132 5428 8188
rect 5428 8132 5432 8188
rect 5368 8128 5432 8132
rect 5448 8188 5512 8192
rect 5448 8132 5452 8188
rect 5452 8132 5508 8188
rect 5508 8132 5512 8188
rect 5448 8128 5512 8132
rect 5528 8188 5592 8192
rect 5528 8132 5532 8188
rect 5532 8132 5588 8188
rect 5588 8132 5592 8188
rect 5528 8128 5592 8132
rect 5608 8188 5672 8192
rect 5608 8132 5612 8188
rect 5612 8132 5668 8188
rect 5668 8132 5672 8188
rect 5608 8128 5672 8132
rect 8312 8188 8376 8192
rect 8312 8132 8316 8188
rect 8316 8132 8372 8188
rect 8372 8132 8376 8188
rect 8312 8128 8376 8132
rect 8392 8188 8456 8192
rect 8392 8132 8396 8188
rect 8396 8132 8452 8188
rect 8452 8132 8456 8188
rect 8392 8128 8456 8132
rect 8472 8188 8536 8192
rect 8472 8132 8476 8188
rect 8476 8132 8532 8188
rect 8532 8132 8536 8188
rect 8472 8128 8536 8132
rect 8552 8188 8616 8192
rect 8552 8132 8556 8188
rect 8556 8132 8612 8188
rect 8612 8132 8616 8188
rect 8552 8128 8616 8132
rect 11256 8188 11320 8192
rect 11256 8132 11260 8188
rect 11260 8132 11316 8188
rect 11316 8132 11320 8188
rect 11256 8128 11320 8132
rect 11336 8188 11400 8192
rect 11336 8132 11340 8188
rect 11340 8132 11396 8188
rect 11396 8132 11400 8188
rect 11336 8128 11400 8132
rect 11416 8188 11480 8192
rect 11416 8132 11420 8188
rect 11420 8132 11476 8188
rect 11476 8132 11480 8188
rect 11416 8128 11480 8132
rect 11496 8188 11560 8192
rect 11496 8132 11500 8188
rect 11500 8132 11556 8188
rect 11556 8132 11560 8188
rect 11496 8128 11560 8132
rect 3896 7644 3960 7648
rect 3896 7588 3900 7644
rect 3900 7588 3956 7644
rect 3956 7588 3960 7644
rect 3896 7584 3960 7588
rect 3976 7644 4040 7648
rect 3976 7588 3980 7644
rect 3980 7588 4036 7644
rect 4036 7588 4040 7644
rect 3976 7584 4040 7588
rect 4056 7644 4120 7648
rect 4056 7588 4060 7644
rect 4060 7588 4116 7644
rect 4116 7588 4120 7644
rect 4056 7584 4120 7588
rect 4136 7644 4200 7648
rect 4136 7588 4140 7644
rect 4140 7588 4196 7644
rect 4196 7588 4200 7644
rect 4136 7584 4200 7588
rect 6840 7644 6904 7648
rect 6840 7588 6844 7644
rect 6844 7588 6900 7644
rect 6900 7588 6904 7644
rect 6840 7584 6904 7588
rect 6920 7644 6984 7648
rect 6920 7588 6924 7644
rect 6924 7588 6980 7644
rect 6980 7588 6984 7644
rect 6920 7584 6984 7588
rect 7000 7644 7064 7648
rect 7000 7588 7004 7644
rect 7004 7588 7060 7644
rect 7060 7588 7064 7644
rect 7000 7584 7064 7588
rect 7080 7644 7144 7648
rect 7080 7588 7084 7644
rect 7084 7588 7140 7644
rect 7140 7588 7144 7644
rect 7080 7584 7144 7588
rect 9784 7644 9848 7648
rect 9784 7588 9788 7644
rect 9788 7588 9844 7644
rect 9844 7588 9848 7644
rect 9784 7584 9848 7588
rect 9864 7644 9928 7648
rect 9864 7588 9868 7644
rect 9868 7588 9924 7644
rect 9924 7588 9928 7644
rect 9864 7584 9928 7588
rect 9944 7644 10008 7648
rect 9944 7588 9948 7644
rect 9948 7588 10004 7644
rect 10004 7588 10008 7644
rect 9944 7584 10008 7588
rect 10024 7644 10088 7648
rect 10024 7588 10028 7644
rect 10028 7588 10084 7644
rect 10084 7588 10088 7644
rect 10024 7584 10088 7588
rect 12728 7644 12792 7648
rect 12728 7588 12732 7644
rect 12732 7588 12788 7644
rect 12788 7588 12792 7644
rect 12728 7584 12792 7588
rect 12808 7644 12872 7648
rect 12808 7588 12812 7644
rect 12812 7588 12868 7644
rect 12868 7588 12872 7644
rect 12808 7584 12872 7588
rect 12888 7644 12952 7648
rect 12888 7588 12892 7644
rect 12892 7588 12948 7644
rect 12948 7588 12952 7644
rect 12888 7584 12952 7588
rect 12968 7644 13032 7648
rect 12968 7588 12972 7644
rect 12972 7588 13028 7644
rect 13028 7588 13032 7644
rect 12968 7584 13032 7588
rect 2424 7100 2488 7104
rect 2424 7044 2428 7100
rect 2428 7044 2484 7100
rect 2484 7044 2488 7100
rect 2424 7040 2488 7044
rect 2504 7100 2568 7104
rect 2504 7044 2508 7100
rect 2508 7044 2564 7100
rect 2564 7044 2568 7100
rect 2504 7040 2568 7044
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 5368 7100 5432 7104
rect 5368 7044 5372 7100
rect 5372 7044 5428 7100
rect 5428 7044 5432 7100
rect 5368 7040 5432 7044
rect 5448 7100 5512 7104
rect 5448 7044 5452 7100
rect 5452 7044 5508 7100
rect 5508 7044 5512 7100
rect 5448 7040 5512 7044
rect 5528 7100 5592 7104
rect 5528 7044 5532 7100
rect 5532 7044 5588 7100
rect 5588 7044 5592 7100
rect 5528 7040 5592 7044
rect 5608 7100 5672 7104
rect 5608 7044 5612 7100
rect 5612 7044 5668 7100
rect 5668 7044 5672 7100
rect 5608 7040 5672 7044
rect 8312 7100 8376 7104
rect 8312 7044 8316 7100
rect 8316 7044 8372 7100
rect 8372 7044 8376 7100
rect 8312 7040 8376 7044
rect 8392 7100 8456 7104
rect 8392 7044 8396 7100
rect 8396 7044 8452 7100
rect 8452 7044 8456 7100
rect 8392 7040 8456 7044
rect 8472 7100 8536 7104
rect 8472 7044 8476 7100
rect 8476 7044 8532 7100
rect 8532 7044 8536 7100
rect 8472 7040 8536 7044
rect 8552 7100 8616 7104
rect 8552 7044 8556 7100
rect 8556 7044 8612 7100
rect 8612 7044 8616 7100
rect 8552 7040 8616 7044
rect 11256 7100 11320 7104
rect 11256 7044 11260 7100
rect 11260 7044 11316 7100
rect 11316 7044 11320 7100
rect 11256 7040 11320 7044
rect 11336 7100 11400 7104
rect 11336 7044 11340 7100
rect 11340 7044 11396 7100
rect 11396 7044 11400 7100
rect 11336 7040 11400 7044
rect 11416 7100 11480 7104
rect 11416 7044 11420 7100
rect 11420 7044 11476 7100
rect 11476 7044 11480 7100
rect 11416 7040 11480 7044
rect 11496 7100 11560 7104
rect 11496 7044 11500 7100
rect 11500 7044 11556 7100
rect 11556 7044 11560 7100
rect 11496 7040 11560 7044
rect 3896 6556 3960 6560
rect 3896 6500 3900 6556
rect 3900 6500 3956 6556
rect 3956 6500 3960 6556
rect 3896 6496 3960 6500
rect 3976 6556 4040 6560
rect 3976 6500 3980 6556
rect 3980 6500 4036 6556
rect 4036 6500 4040 6556
rect 3976 6496 4040 6500
rect 4056 6556 4120 6560
rect 4056 6500 4060 6556
rect 4060 6500 4116 6556
rect 4116 6500 4120 6556
rect 4056 6496 4120 6500
rect 4136 6556 4200 6560
rect 4136 6500 4140 6556
rect 4140 6500 4196 6556
rect 4196 6500 4200 6556
rect 4136 6496 4200 6500
rect 6840 6556 6904 6560
rect 6840 6500 6844 6556
rect 6844 6500 6900 6556
rect 6900 6500 6904 6556
rect 6840 6496 6904 6500
rect 6920 6556 6984 6560
rect 6920 6500 6924 6556
rect 6924 6500 6980 6556
rect 6980 6500 6984 6556
rect 6920 6496 6984 6500
rect 7000 6556 7064 6560
rect 7000 6500 7004 6556
rect 7004 6500 7060 6556
rect 7060 6500 7064 6556
rect 7000 6496 7064 6500
rect 7080 6556 7144 6560
rect 7080 6500 7084 6556
rect 7084 6500 7140 6556
rect 7140 6500 7144 6556
rect 7080 6496 7144 6500
rect 9784 6556 9848 6560
rect 9784 6500 9788 6556
rect 9788 6500 9844 6556
rect 9844 6500 9848 6556
rect 9784 6496 9848 6500
rect 9864 6556 9928 6560
rect 9864 6500 9868 6556
rect 9868 6500 9924 6556
rect 9924 6500 9928 6556
rect 9864 6496 9928 6500
rect 9944 6556 10008 6560
rect 9944 6500 9948 6556
rect 9948 6500 10004 6556
rect 10004 6500 10008 6556
rect 9944 6496 10008 6500
rect 10024 6556 10088 6560
rect 10024 6500 10028 6556
rect 10028 6500 10084 6556
rect 10084 6500 10088 6556
rect 10024 6496 10088 6500
rect 12728 6556 12792 6560
rect 12728 6500 12732 6556
rect 12732 6500 12788 6556
rect 12788 6500 12792 6556
rect 12728 6496 12792 6500
rect 12808 6556 12872 6560
rect 12808 6500 12812 6556
rect 12812 6500 12868 6556
rect 12868 6500 12872 6556
rect 12808 6496 12872 6500
rect 12888 6556 12952 6560
rect 12888 6500 12892 6556
rect 12892 6500 12948 6556
rect 12948 6500 12952 6556
rect 12888 6496 12952 6500
rect 12968 6556 13032 6560
rect 12968 6500 12972 6556
rect 12972 6500 13028 6556
rect 13028 6500 13032 6556
rect 12968 6496 13032 6500
rect 2424 6012 2488 6016
rect 2424 5956 2428 6012
rect 2428 5956 2484 6012
rect 2484 5956 2488 6012
rect 2424 5952 2488 5956
rect 2504 6012 2568 6016
rect 2504 5956 2508 6012
rect 2508 5956 2564 6012
rect 2564 5956 2568 6012
rect 2504 5952 2568 5956
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 5368 6012 5432 6016
rect 5368 5956 5372 6012
rect 5372 5956 5428 6012
rect 5428 5956 5432 6012
rect 5368 5952 5432 5956
rect 5448 6012 5512 6016
rect 5448 5956 5452 6012
rect 5452 5956 5508 6012
rect 5508 5956 5512 6012
rect 5448 5952 5512 5956
rect 5528 6012 5592 6016
rect 5528 5956 5532 6012
rect 5532 5956 5588 6012
rect 5588 5956 5592 6012
rect 5528 5952 5592 5956
rect 5608 6012 5672 6016
rect 5608 5956 5612 6012
rect 5612 5956 5668 6012
rect 5668 5956 5672 6012
rect 5608 5952 5672 5956
rect 8312 6012 8376 6016
rect 8312 5956 8316 6012
rect 8316 5956 8372 6012
rect 8372 5956 8376 6012
rect 8312 5952 8376 5956
rect 8392 6012 8456 6016
rect 8392 5956 8396 6012
rect 8396 5956 8452 6012
rect 8452 5956 8456 6012
rect 8392 5952 8456 5956
rect 8472 6012 8536 6016
rect 8472 5956 8476 6012
rect 8476 5956 8532 6012
rect 8532 5956 8536 6012
rect 8472 5952 8536 5956
rect 8552 6012 8616 6016
rect 8552 5956 8556 6012
rect 8556 5956 8612 6012
rect 8612 5956 8616 6012
rect 8552 5952 8616 5956
rect 11256 6012 11320 6016
rect 11256 5956 11260 6012
rect 11260 5956 11316 6012
rect 11316 5956 11320 6012
rect 11256 5952 11320 5956
rect 11336 6012 11400 6016
rect 11336 5956 11340 6012
rect 11340 5956 11396 6012
rect 11396 5956 11400 6012
rect 11336 5952 11400 5956
rect 11416 6012 11480 6016
rect 11416 5956 11420 6012
rect 11420 5956 11476 6012
rect 11476 5956 11480 6012
rect 11416 5952 11480 5956
rect 11496 6012 11560 6016
rect 11496 5956 11500 6012
rect 11500 5956 11556 6012
rect 11556 5956 11560 6012
rect 11496 5952 11560 5956
rect 3896 5468 3960 5472
rect 3896 5412 3900 5468
rect 3900 5412 3956 5468
rect 3956 5412 3960 5468
rect 3896 5408 3960 5412
rect 3976 5468 4040 5472
rect 3976 5412 3980 5468
rect 3980 5412 4036 5468
rect 4036 5412 4040 5468
rect 3976 5408 4040 5412
rect 4056 5468 4120 5472
rect 4056 5412 4060 5468
rect 4060 5412 4116 5468
rect 4116 5412 4120 5468
rect 4056 5408 4120 5412
rect 4136 5468 4200 5472
rect 4136 5412 4140 5468
rect 4140 5412 4196 5468
rect 4196 5412 4200 5468
rect 4136 5408 4200 5412
rect 6840 5468 6904 5472
rect 6840 5412 6844 5468
rect 6844 5412 6900 5468
rect 6900 5412 6904 5468
rect 6840 5408 6904 5412
rect 6920 5468 6984 5472
rect 6920 5412 6924 5468
rect 6924 5412 6980 5468
rect 6980 5412 6984 5468
rect 6920 5408 6984 5412
rect 7000 5468 7064 5472
rect 7000 5412 7004 5468
rect 7004 5412 7060 5468
rect 7060 5412 7064 5468
rect 7000 5408 7064 5412
rect 7080 5468 7144 5472
rect 7080 5412 7084 5468
rect 7084 5412 7140 5468
rect 7140 5412 7144 5468
rect 7080 5408 7144 5412
rect 9784 5468 9848 5472
rect 9784 5412 9788 5468
rect 9788 5412 9844 5468
rect 9844 5412 9848 5468
rect 9784 5408 9848 5412
rect 9864 5468 9928 5472
rect 9864 5412 9868 5468
rect 9868 5412 9924 5468
rect 9924 5412 9928 5468
rect 9864 5408 9928 5412
rect 9944 5468 10008 5472
rect 9944 5412 9948 5468
rect 9948 5412 10004 5468
rect 10004 5412 10008 5468
rect 9944 5408 10008 5412
rect 10024 5468 10088 5472
rect 10024 5412 10028 5468
rect 10028 5412 10084 5468
rect 10084 5412 10088 5468
rect 10024 5408 10088 5412
rect 12728 5468 12792 5472
rect 12728 5412 12732 5468
rect 12732 5412 12788 5468
rect 12788 5412 12792 5468
rect 12728 5408 12792 5412
rect 12808 5468 12872 5472
rect 12808 5412 12812 5468
rect 12812 5412 12868 5468
rect 12868 5412 12872 5468
rect 12808 5408 12872 5412
rect 12888 5468 12952 5472
rect 12888 5412 12892 5468
rect 12892 5412 12948 5468
rect 12948 5412 12952 5468
rect 12888 5408 12952 5412
rect 12968 5468 13032 5472
rect 12968 5412 12972 5468
rect 12972 5412 13028 5468
rect 13028 5412 13032 5468
rect 12968 5408 13032 5412
rect 2424 4924 2488 4928
rect 2424 4868 2428 4924
rect 2428 4868 2484 4924
rect 2484 4868 2488 4924
rect 2424 4864 2488 4868
rect 2504 4924 2568 4928
rect 2504 4868 2508 4924
rect 2508 4868 2564 4924
rect 2564 4868 2568 4924
rect 2504 4864 2568 4868
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 5368 4924 5432 4928
rect 5368 4868 5372 4924
rect 5372 4868 5428 4924
rect 5428 4868 5432 4924
rect 5368 4864 5432 4868
rect 5448 4924 5512 4928
rect 5448 4868 5452 4924
rect 5452 4868 5508 4924
rect 5508 4868 5512 4924
rect 5448 4864 5512 4868
rect 5528 4924 5592 4928
rect 5528 4868 5532 4924
rect 5532 4868 5588 4924
rect 5588 4868 5592 4924
rect 5528 4864 5592 4868
rect 5608 4924 5672 4928
rect 5608 4868 5612 4924
rect 5612 4868 5668 4924
rect 5668 4868 5672 4924
rect 5608 4864 5672 4868
rect 8312 4924 8376 4928
rect 8312 4868 8316 4924
rect 8316 4868 8372 4924
rect 8372 4868 8376 4924
rect 8312 4864 8376 4868
rect 8392 4924 8456 4928
rect 8392 4868 8396 4924
rect 8396 4868 8452 4924
rect 8452 4868 8456 4924
rect 8392 4864 8456 4868
rect 8472 4924 8536 4928
rect 8472 4868 8476 4924
rect 8476 4868 8532 4924
rect 8532 4868 8536 4924
rect 8472 4864 8536 4868
rect 8552 4924 8616 4928
rect 8552 4868 8556 4924
rect 8556 4868 8612 4924
rect 8612 4868 8616 4924
rect 8552 4864 8616 4868
rect 11256 4924 11320 4928
rect 11256 4868 11260 4924
rect 11260 4868 11316 4924
rect 11316 4868 11320 4924
rect 11256 4864 11320 4868
rect 11336 4924 11400 4928
rect 11336 4868 11340 4924
rect 11340 4868 11396 4924
rect 11396 4868 11400 4924
rect 11336 4864 11400 4868
rect 11416 4924 11480 4928
rect 11416 4868 11420 4924
rect 11420 4868 11476 4924
rect 11476 4868 11480 4924
rect 11416 4864 11480 4868
rect 11496 4924 11560 4928
rect 11496 4868 11500 4924
rect 11500 4868 11556 4924
rect 11556 4868 11560 4924
rect 11496 4864 11560 4868
rect 3896 4380 3960 4384
rect 3896 4324 3900 4380
rect 3900 4324 3956 4380
rect 3956 4324 3960 4380
rect 3896 4320 3960 4324
rect 3976 4380 4040 4384
rect 3976 4324 3980 4380
rect 3980 4324 4036 4380
rect 4036 4324 4040 4380
rect 3976 4320 4040 4324
rect 4056 4380 4120 4384
rect 4056 4324 4060 4380
rect 4060 4324 4116 4380
rect 4116 4324 4120 4380
rect 4056 4320 4120 4324
rect 4136 4380 4200 4384
rect 4136 4324 4140 4380
rect 4140 4324 4196 4380
rect 4196 4324 4200 4380
rect 4136 4320 4200 4324
rect 6840 4380 6904 4384
rect 6840 4324 6844 4380
rect 6844 4324 6900 4380
rect 6900 4324 6904 4380
rect 6840 4320 6904 4324
rect 6920 4380 6984 4384
rect 6920 4324 6924 4380
rect 6924 4324 6980 4380
rect 6980 4324 6984 4380
rect 6920 4320 6984 4324
rect 7000 4380 7064 4384
rect 7000 4324 7004 4380
rect 7004 4324 7060 4380
rect 7060 4324 7064 4380
rect 7000 4320 7064 4324
rect 7080 4380 7144 4384
rect 7080 4324 7084 4380
rect 7084 4324 7140 4380
rect 7140 4324 7144 4380
rect 7080 4320 7144 4324
rect 9784 4380 9848 4384
rect 9784 4324 9788 4380
rect 9788 4324 9844 4380
rect 9844 4324 9848 4380
rect 9784 4320 9848 4324
rect 9864 4380 9928 4384
rect 9864 4324 9868 4380
rect 9868 4324 9924 4380
rect 9924 4324 9928 4380
rect 9864 4320 9928 4324
rect 9944 4380 10008 4384
rect 9944 4324 9948 4380
rect 9948 4324 10004 4380
rect 10004 4324 10008 4380
rect 9944 4320 10008 4324
rect 10024 4380 10088 4384
rect 10024 4324 10028 4380
rect 10028 4324 10084 4380
rect 10084 4324 10088 4380
rect 10024 4320 10088 4324
rect 12728 4380 12792 4384
rect 12728 4324 12732 4380
rect 12732 4324 12788 4380
rect 12788 4324 12792 4380
rect 12728 4320 12792 4324
rect 12808 4380 12872 4384
rect 12808 4324 12812 4380
rect 12812 4324 12868 4380
rect 12868 4324 12872 4380
rect 12808 4320 12872 4324
rect 12888 4380 12952 4384
rect 12888 4324 12892 4380
rect 12892 4324 12948 4380
rect 12948 4324 12952 4380
rect 12888 4320 12952 4324
rect 12968 4380 13032 4384
rect 12968 4324 12972 4380
rect 12972 4324 13028 4380
rect 13028 4324 13032 4380
rect 12968 4320 13032 4324
rect 2424 3836 2488 3840
rect 2424 3780 2428 3836
rect 2428 3780 2484 3836
rect 2484 3780 2488 3836
rect 2424 3776 2488 3780
rect 2504 3836 2568 3840
rect 2504 3780 2508 3836
rect 2508 3780 2564 3836
rect 2564 3780 2568 3836
rect 2504 3776 2568 3780
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 5368 3836 5432 3840
rect 5368 3780 5372 3836
rect 5372 3780 5428 3836
rect 5428 3780 5432 3836
rect 5368 3776 5432 3780
rect 5448 3836 5512 3840
rect 5448 3780 5452 3836
rect 5452 3780 5508 3836
rect 5508 3780 5512 3836
rect 5448 3776 5512 3780
rect 5528 3836 5592 3840
rect 5528 3780 5532 3836
rect 5532 3780 5588 3836
rect 5588 3780 5592 3836
rect 5528 3776 5592 3780
rect 5608 3836 5672 3840
rect 5608 3780 5612 3836
rect 5612 3780 5668 3836
rect 5668 3780 5672 3836
rect 5608 3776 5672 3780
rect 8312 3836 8376 3840
rect 8312 3780 8316 3836
rect 8316 3780 8372 3836
rect 8372 3780 8376 3836
rect 8312 3776 8376 3780
rect 8392 3836 8456 3840
rect 8392 3780 8396 3836
rect 8396 3780 8452 3836
rect 8452 3780 8456 3836
rect 8392 3776 8456 3780
rect 8472 3836 8536 3840
rect 8472 3780 8476 3836
rect 8476 3780 8532 3836
rect 8532 3780 8536 3836
rect 8472 3776 8536 3780
rect 8552 3836 8616 3840
rect 8552 3780 8556 3836
rect 8556 3780 8612 3836
rect 8612 3780 8616 3836
rect 8552 3776 8616 3780
rect 11256 3836 11320 3840
rect 11256 3780 11260 3836
rect 11260 3780 11316 3836
rect 11316 3780 11320 3836
rect 11256 3776 11320 3780
rect 11336 3836 11400 3840
rect 11336 3780 11340 3836
rect 11340 3780 11396 3836
rect 11396 3780 11400 3836
rect 11336 3776 11400 3780
rect 11416 3836 11480 3840
rect 11416 3780 11420 3836
rect 11420 3780 11476 3836
rect 11476 3780 11480 3836
rect 11416 3776 11480 3780
rect 11496 3836 11560 3840
rect 11496 3780 11500 3836
rect 11500 3780 11556 3836
rect 11556 3780 11560 3836
rect 11496 3776 11560 3780
rect 3896 3292 3960 3296
rect 3896 3236 3900 3292
rect 3900 3236 3956 3292
rect 3956 3236 3960 3292
rect 3896 3232 3960 3236
rect 3976 3292 4040 3296
rect 3976 3236 3980 3292
rect 3980 3236 4036 3292
rect 4036 3236 4040 3292
rect 3976 3232 4040 3236
rect 4056 3292 4120 3296
rect 4056 3236 4060 3292
rect 4060 3236 4116 3292
rect 4116 3236 4120 3292
rect 4056 3232 4120 3236
rect 4136 3292 4200 3296
rect 4136 3236 4140 3292
rect 4140 3236 4196 3292
rect 4196 3236 4200 3292
rect 4136 3232 4200 3236
rect 6840 3292 6904 3296
rect 6840 3236 6844 3292
rect 6844 3236 6900 3292
rect 6900 3236 6904 3292
rect 6840 3232 6904 3236
rect 6920 3292 6984 3296
rect 6920 3236 6924 3292
rect 6924 3236 6980 3292
rect 6980 3236 6984 3292
rect 6920 3232 6984 3236
rect 7000 3292 7064 3296
rect 7000 3236 7004 3292
rect 7004 3236 7060 3292
rect 7060 3236 7064 3292
rect 7000 3232 7064 3236
rect 7080 3292 7144 3296
rect 7080 3236 7084 3292
rect 7084 3236 7140 3292
rect 7140 3236 7144 3292
rect 7080 3232 7144 3236
rect 9784 3292 9848 3296
rect 9784 3236 9788 3292
rect 9788 3236 9844 3292
rect 9844 3236 9848 3292
rect 9784 3232 9848 3236
rect 9864 3292 9928 3296
rect 9864 3236 9868 3292
rect 9868 3236 9924 3292
rect 9924 3236 9928 3292
rect 9864 3232 9928 3236
rect 9944 3292 10008 3296
rect 9944 3236 9948 3292
rect 9948 3236 10004 3292
rect 10004 3236 10008 3292
rect 9944 3232 10008 3236
rect 10024 3292 10088 3296
rect 10024 3236 10028 3292
rect 10028 3236 10084 3292
rect 10084 3236 10088 3292
rect 10024 3232 10088 3236
rect 12728 3292 12792 3296
rect 12728 3236 12732 3292
rect 12732 3236 12788 3292
rect 12788 3236 12792 3292
rect 12728 3232 12792 3236
rect 12808 3292 12872 3296
rect 12808 3236 12812 3292
rect 12812 3236 12868 3292
rect 12868 3236 12872 3292
rect 12808 3232 12872 3236
rect 12888 3292 12952 3296
rect 12888 3236 12892 3292
rect 12892 3236 12948 3292
rect 12948 3236 12952 3292
rect 12888 3232 12952 3236
rect 12968 3292 13032 3296
rect 12968 3236 12972 3292
rect 12972 3236 13028 3292
rect 13028 3236 13032 3292
rect 12968 3232 13032 3236
rect 2424 2748 2488 2752
rect 2424 2692 2428 2748
rect 2428 2692 2484 2748
rect 2484 2692 2488 2748
rect 2424 2688 2488 2692
rect 2504 2748 2568 2752
rect 2504 2692 2508 2748
rect 2508 2692 2564 2748
rect 2564 2692 2568 2748
rect 2504 2688 2568 2692
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 5368 2748 5432 2752
rect 5368 2692 5372 2748
rect 5372 2692 5428 2748
rect 5428 2692 5432 2748
rect 5368 2688 5432 2692
rect 5448 2748 5512 2752
rect 5448 2692 5452 2748
rect 5452 2692 5508 2748
rect 5508 2692 5512 2748
rect 5448 2688 5512 2692
rect 5528 2748 5592 2752
rect 5528 2692 5532 2748
rect 5532 2692 5588 2748
rect 5588 2692 5592 2748
rect 5528 2688 5592 2692
rect 5608 2748 5672 2752
rect 5608 2692 5612 2748
rect 5612 2692 5668 2748
rect 5668 2692 5672 2748
rect 5608 2688 5672 2692
rect 8312 2748 8376 2752
rect 8312 2692 8316 2748
rect 8316 2692 8372 2748
rect 8372 2692 8376 2748
rect 8312 2688 8376 2692
rect 8392 2748 8456 2752
rect 8392 2692 8396 2748
rect 8396 2692 8452 2748
rect 8452 2692 8456 2748
rect 8392 2688 8456 2692
rect 8472 2748 8536 2752
rect 8472 2692 8476 2748
rect 8476 2692 8532 2748
rect 8532 2692 8536 2748
rect 8472 2688 8536 2692
rect 8552 2748 8616 2752
rect 8552 2692 8556 2748
rect 8556 2692 8612 2748
rect 8612 2692 8616 2748
rect 8552 2688 8616 2692
rect 11256 2748 11320 2752
rect 11256 2692 11260 2748
rect 11260 2692 11316 2748
rect 11316 2692 11320 2748
rect 11256 2688 11320 2692
rect 11336 2748 11400 2752
rect 11336 2692 11340 2748
rect 11340 2692 11396 2748
rect 11396 2692 11400 2748
rect 11336 2688 11400 2692
rect 11416 2748 11480 2752
rect 11416 2692 11420 2748
rect 11420 2692 11476 2748
rect 11476 2692 11480 2748
rect 11416 2688 11480 2692
rect 11496 2748 11560 2752
rect 11496 2692 11500 2748
rect 11500 2692 11556 2748
rect 11556 2692 11560 2748
rect 11496 2688 11560 2692
rect 3896 2204 3960 2208
rect 3896 2148 3900 2204
rect 3900 2148 3956 2204
rect 3956 2148 3960 2204
rect 3896 2144 3960 2148
rect 3976 2204 4040 2208
rect 3976 2148 3980 2204
rect 3980 2148 4036 2204
rect 4036 2148 4040 2204
rect 3976 2144 4040 2148
rect 4056 2204 4120 2208
rect 4056 2148 4060 2204
rect 4060 2148 4116 2204
rect 4116 2148 4120 2204
rect 4056 2144 4120 2148
rect 4136 2204 4200 2208
rect 4136 2148 4140 2204
rect 4140 2148 4196 2204
rect 4196 2148 4200 2204
rect 4136 2144 4200 2148
rect 6840 2204 6904 2208
rect 6840 2148 6844 2204
rect 6844 2148 6900 2204
rect 6900 2148 6904 2204
rect 6840 2144 6904 2148
rect 6920 2204 6984 2208
rect 6920 2148 6924 2204
rect 6924 2148 6980 2204
rect 6980 2148 6984 2204
rect 6920 2144 6984 2148
rect 7000 2204 7064 2208
rect 7000 2148 7004 2204
rect 7004 2148 7060 2204
rect 7060 2148 7064 2204
rect 7000 2144 7064 2148
rect 7080 2204 7144 2208
rect 7080 2148 7084 2204
rect 7084 2148 7140 2204
rect 7140 2148 7144 2204
rect 7080 2144 7144 2148
rect 9784 2204 9848 2208
rect 9784 2148 9788 2204
rect 9788 2148 9844 2204
rect 9844 2148 9848 2204
rect 9784 2144 9848 2148
rect 9864 2204 9928 2208
rect 9864 2148 9868 2204
rect 9868 2148 9924 2204
rect 9924 2148 9928 2204
rect 9864 2144 9928 2148
rect 9944 2204 10008 2208
rect 9944 2148 9948 2204
rect 9948 2148 10004 2204
rect 10004 2148 10008 2204
rect 9944 2144 10008 2148
rect 10024 2204 10088 2208
rect 10024 2148 10028 2204
rect 10028 2148 10084 2204
rect 10084 2148 10088 2204
rect 10024 2144 10088 2148
rect 12728 2204 12792 2208
rect 12728 2148 12732 2204
rect 12732 2148 12788 2204
rect 12788 2148 12792 2204
rect 12728 2144 12792 2148
rect 12808 2204 12872 2208
rect 12808 2148 12812 2204
rect 12812 2148 12868 2204
rect 12868 2148 12872 2204
rect 12808 2144 12872 2148
rect 12888 2204 12952 2208
rect 12888 2148 12892 2204
rect 12892 2148 12948 2204
rect 12948 2148 12952 2204
rect 12888 2144 12952 2148
rect 12968 2204 13032 2208
rect 12968 2148 12972 2204
rect 12972 2148 13028 2204
rect 13028 2148 13032 2204
rect 12968 2144 13032 2148
<< metal4 >>
rect 2416 11456 2736 11472
rect 2416 11392 2424 11456
rect 2488 11392 2504 11456
rect 2568 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2736 11456
rect 2416 10368 2736 11392
rect 2416 10304 2424 10368
rect 2488 10304 2504 10368
rect 2568 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2736 10368
rect 2416 9280 2736 10304
rect 2416 9216 2424 9280
rect 2488 9216 2504 9280
rect 2568 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2736 9280
rect 2416 8192 2736 9216
rect 2416 8128 2424 8192
rect 2488 8128 2504 8192
rect 2568 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2736 8192
rect 2416 7104 2736 8128
rect 2416 7040 2424 7104
rect 2488 7040 2504 7104
rect 2568 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2736 7104
rect 2416 6016 2736 7040
rect 2416 5952 2424 6016
rect 2488 5952 2504 6016
rect 2568 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2736 6016
rect 2416 4928 2736 5952
rect 2416 4864 2424 4928
rect 2488 4864 2504 4928
rect 2568 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2736 4928
rect 2416 3840 2736 4864
rect 2416 3776 2424 3840
rect 2488 3776 2504 3840
rect 2568 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2736 3840
rect 2416 2752 2736 3776
rect 2416 2688 2424 2752
rect 2488 2688 2504 2752
rect 2568 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2736 2752
rect 2416 2128 2736 2688
rect 3888 10912 4208 11472
rect 3888 10848 3896 10912
rect 3960 10848 3976 10912
rect 4040 10848 4056 10912
rect 4120 10848 4136 10912
rect 4200 10848 4208 10912
rect 3888 9824 4208 10848
rect 3888 9760 3896 9824
rect 3960 9760 3976 9824
rect 4040 9760 4056 9824
rect 4120 9760 4136 9824
rect 4200 9760 4208 9824
rect 3888 8736 4208 9760
rect 3888 8672 3896 8736
rect 3960 8672 3976 8736
rect 4040 8672 4056 8736
rect 4120 8672 4136 8736
rect 4200 8672 4208 8736
rect 3888 7648 4208 8672
rect 3888 7584 3896 7648
rect 3960 7584 3976 7648
rect 4040 7584 4056 7648
rect 4120 7584 4136 7648
rect 4200 7584 4208 7648
rect 3888 6560 4208 7584
rect 3888 6496 3896 6560
rect 3960 6496 3976 6560
rect 4040 6496 4056 6560
rect 4120 6496 4136 6560
rect 4200 6496 4208 6560
rect 3888 5472 4208 6496
rect 3888 5408 3896 5472
rect 3960 5408 3976 5472
rect 4040 5408 4056 5472
rect 4120 5408 4136 5472
rect 4200 5408 4208 5472
rect 3888 4384 4208 5408
rect 3888 4320 3896 4384
rect 3960 4320 3976 4384
rect 4040 4320 4056 4384
rect 4120 4320 4136 4384
rect 4200 4320 4208 4384
rect 3888 3296 4208 4320
rect 3888 3232 3896 3296
rect 3960 3232 3976 3296
rect 4040 3232 4056 3296
rect 4120 3232 4136 3296
rect 4200 3232 4208 3296
rect 3888 2208 4208 3232
rect 3888 2144 3896 2208
rect 3960 2144 3976 2208
rect 4040 2144 4056 2208
rect 4120 2144 4136 2208
rect 4200 2144 4208 2208
rect 3888 2128 4208 2144
rect 5360 11456 5680 11472
rect 5360 11392 5368 11456
rect 5432 11392 5448 11456
rect 5512 11392 5528 11456
rect 5592 11392 5608 11456
rect 5672 11392 5680 11456
rect 5360 10368 5680 11392
rect 5360 10304 5368 10368
rect 5432 10304 5448 10368
rect 5512 10304 5528 10368
rect 5592 10304 5608 10368
rect 5672 10304 5680 10368
rect 5360 9280 5680 10304
rect 5360 9216 5368 9280
rect 5432 9216 5448 9280
rect 5512 9216 5528 9280
rect 5592 9216 5608 9280
rect 5672 9216 5680 9280
rect 5360 8192 5680 9216
rect 5360 8128 5368 8192
rect 5432 8128 5448 8192
rect 5512 8128 5528 8192
rect 5592 8128 5608 8192
rect 5672 8128 5680 8192
rect 5360 7104 5680 8128
rect 5360 7040 5368 7104
rect 5432 7040 5448 7104
rect 5512 7040 5528 7104
rect 5592 7040 5608 7104
rect 5672 7040 5680 7104
rect 5360 6016 5680 7040
rect 5360 5952 5368 6016
rect 5432 5952 5448 6016
rect 5512 5952 5528 6016
rect 5592 5952 5608 6016
rect 5672 5952 5680 6016
rect 5360 4928 5680 5952
rect 5360 4864 5368 4928
rect 5432 4864 5448 4928
rect 5512 4864 5528 4928
rect 5592 4864 5608 4928
rect 5672 4864 5680 4928
rect 5360 3840 5680 4864
rect 5360 3776 5368 3840
rect 5432 3776 5448 3840
rect 5512 3776 5528 3840
rect 5592 3776 5608 3840
rect 5672 3776 5680 3840
rect 5360 2752 5680 3776
rect 5360 2688 5368 2752
rect 5432 2688 5448 2752
rect 5512 2688 5528 2752
rect 5592 2688 5608 2752
rect 5672 2688 5680 2752
rect 5360 2128 5680 2688
rect 6832 10912 7152 11472
rect 6832 10848 6840 10912
rect 6904 10848 6920 10912
rect 6984 10848 7000 10912
rect 7064 10848 7080 10912
rect 7144 10848 7152 10912
rect 6832 9824 7152 10848
rect 6832 9760 6840 9824
rect 6904 9760 6920 9824
rect 6984 9760 7000 9824
rect 7064 9760 7080 9824
rect 7144 9760 7152 9824
rect 6832 8736 7152 9760
rect 6832 8672 6840 8736
rect 6904 8672 6920 8736
rect 6984 8672 7000 8736
rect 7064 8672 7080 8736
rect 7144 8672 7152 8736
rect 6832 7648 7152 8672
rect 6832 7584 6840 7648
rect 6904 7584 6920 7648
rect 6984 7584 7000 7648
rect 7064 7584 7080 7648
rect 7144 7584 7152 7648
rect 6832 6560 7152 7584
rect 6832 6496 6840 6560
rect 6904 6496 6920 6560
rect 6984 6496 7000 6560
rect 7064 6496 7080 6560
rect 7144 6496 7152 6560
rect 6832 5472 7152 6496
rect 6832 5408 6840 5472
rect 6904 5408 6920 5472
rect 6984 5408 7000 5472
rect 7064 5408 7080 5472
rect 7144 5408 7152 5472
rect 6832 4384 7152 5408
rect 6832 4320 6840 4384
rect 6904 4320 6920 4384
rect 6984 4320 7000 4384
rect 7064 4320 7080 4384
rect 7144 4320 7152 4384
rect 6832 3296 7152 4320
rect 6832 3232 6840 3296
rect 6904 3232 6920 3296
rect 6984 3232 7000 3296
rect 7064 3232 7080 3296
rect 7144 3232 7152 3296
rect 6832 2208 7152 3232
rect 6832 2144 6840 2208
rect 6904 2144 6920 2208
rect 6984 2144 7000 2208
rect 7064 2144 7080 2208
rect 7144 2144 7152 2208
rect 6832 2128 7152 2144
rect 8304 11456 8624 11472
rect 8304 11392 8312 11456
rect 8376 11392 8392 11456
rect 8456 11392 8472 11456
rect 8536 11392 8552 11456
rect 8616 11392 8624 11456
rect 8304 10368 8624 11392
rect 8304 10304 8312 10368
rect 8376 10304 8392 10368
rect 8456 10304 8472 10368
rect 8536 10304 8552 10368
rect 8616 10304 8624 10368
rect 8304 9280 8624 10304
rect 8304 9216 8312 9280
rect 8376 9216 8392 9280
rect 8456 9216 8472 9280
rect 8536 9216 8552 9280
rect 8616 9216 8624 9280
rect 8304 8192 8624 9216
rect 8304 8128 8312 8192
rect 8376 8128 8392 8192
rect 8456 8128 8472 8192
rect 8536 8128 8552 8192
rect 8616 8128 8624 8192
rect 8304 7104 8624 8128
rect 8304 7040 8312 7104
rect 8376 7040 8392 7104
rect 8456 7040 8472 7104
rect 8536 7040 8552 7104
rect 8616 7040 8624 7104
rect 8304 6016 8624 7040
rect 8304 5952 8312 6016
rect 8376 5952 8392 6016
rect 8456 5952 8472 6016
rect 8536 5952 8552 6016
rect 8616 5952 8624 6016
rect 8304 4928 8624 5952
rect 8304 4864 8312 4928
rect 8376 4864 8392 4928
rect 8456 4864 8472 4928
rect 8536 4864 8552 4928
rect 8616 4864 8624 4928
rect 8304 3840 8624 4864
rect 8304 3776 8312 3840
rect 8376 3776 8392 3840
rect 8456 3776 8472 3840
rect 8536 3776 8552 3840
rect 8616 3776 8624 3840
rect 8304 2752 8624 3776
rect 8304 2688 8312 2752
rect 8376 2688 8392 2752
rect 8456 2688 8472 2752
rect 8536 2688 8552 2752
rect 8616 2688 8624 2752
rect 8304 2128 8624 2688
rect 9776 10912 10096 11472
rect 9776 10848 9784 10912
rect 9848 10848 9864 10912
rect 9928 10848 9944 10912
rect 10008 10848 10024 10912
rect 10088 10848 10096 10912
rect 9776 9824 10096 10848
rect 9776 9760 9784 9824
rect 9848 9760 9864 9824
rect 9928 9760 9944 9824
rect 10008 9760 10024 9824
rect 10088 9760 10096 9824
rect 9776 8736 10096 9760
rect 9776 8672 9784 8736
rect 9848 8672 9864 8736
rect 9928 8672 9944 8736
rect 10008 8672 10024 8736
rect 10088 8672 10096 8736
rect 9776 7648 10096 8672
rect 9776 7584 9784 7648
rect 9848 7584 9864 7648
rect 9928 7584 9944 7648
rect 10008 7584 10024 7648
rect 10088 7584 10096 7648
rect 9776 6560 10096 7584
rect 9776 6496 9784 6560
rect 9848 6496 9864 6560
rect 9928 6496 9944 6560
rect 10008 6496 10024 6560
rect 10088 6496 10096 6560
rect 9776 5472 10096 6496
rect 9776 5408 9784 5472
rect 9848 5408 9864 5472
rect 9928 5408 9944 5472
rect 10008 5408 10024 5472
rect 10088 5408 10096 5472
rect 9776 4384 10096 5408
rect 9776 4320 9784 4384
rect 9848 4320 9864 4384
rect 9928 4320 9944 4384
rect 10008 4320 10024 4384
rect 10088 4320 10096 4384
rect 9776 3296 10096 4320
rect 9776 3232 9784 3296
rect 9848 3232 9864 3296
rect 9928 3232 9944 3296
rect 10008 3232 10024 3296
rect 10088 3232 10096 3296
rect 9776 2208 10096 3232
rect 9776 2144 9784 2208
rect 9848 2144 9864 2208
rect 9928 2144 9944 2208
rect 10008 2144 10024 2208
rect 10088 2144 10096 2208
rect 9776 2128 10096 2144
rect 11248 11456 11568 11472
rect 11248 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11568 11456
rect 11248 10368 11568 11392
rect 11248 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11568 10368
rect 11248 9280 11568 10304
rect 11248 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11568 9280
rect 11248 8192 11568 9216
rect 11248 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11568 8192
rect 11248 7104 11568 8128
rect 11248 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11568 7104
rect 11248 6016 11568 7040
rect 11248 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11568 6016
rect 11248 4928 11568 5952
rect 11248 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11568 4928
rect 11248 3840 11568 4864
rect 11248 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11568 3840
rect 11248 2752 11568 3776
rect 11248 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11568 2752
rect 11248 2128 11568 2688
rect 12720 10912 13040 11472
rect 12720 10848 12728 10912
rect 12792 10848 12808 10912
rect 12872 10848 12888 10912
rect 12952 10848 12968 10912
rect 13032 10848 13040 10912
rect 12720 9824 13040 10848
rect 12720 9760 12728 9824
rect 12792 9760 12808 9824
rect 12872 9760 12888 9824
rect 12952 9760 12968 9824
rect 13032 9760 13040 9824
rect 12720 8736 13040 9760
rect 12720 8672 12728 8736
rect 12792 8672 12808 8736
rect 12872 8672 12888 8736
rect 12952 8672 12968 8736
rect 13032 8672 13040 8736
rect 12720 7648 13040 8672
rect 12720 7584 12728 7648
rect 12792 7584 12808 7648
rect 12872 7584 12888 7648
rect 12952 7584 12968 7648
rect 13032 7584 13040 7648
rect 12720 6560 13040 7584
rect 12720 6496 12728 6560
rect 12792 6496 12808 6560
rect 12872 6496 12888 6560
rect 12952 6496 12968 6560
rect 13032 6496 13040 6560
rect 12720 5472 13040 6496
rect 12720 5408 12728 5472
rect 12792 5408 12808 5472
rect 12872 5408 12888 5472
rect 12952 5408 12968 5472
rect 13032 5408 13040 5472
rect 12720 4384 13040 5408
rect 12720 4320 12728 4384
rect 12792 4320 12808 4384
rect 12872 4320 12888 4384
rect 12952 4320 12968 4384
rect 13032 4320 13040 4384
rect 12720 3296 13040 4320
rect 12720 3232 12728 3296
rect 12792 3232 12808 3296
rect 12872 3232 12888 3296
rect 12952 3232 12968 3296
rect 13032 3232 13040 3296
rect 12720 2208 13040 3232
rect 12720 2144 12728 2208
rect 12792 2144 12808 2208
rect 12872 2144 12888 2208
rect 12952 2144 12968 2208
rect 13032 2144 13040 2208
rect 12720 2128 13040 2144
use sky130_fd_sc_hd__inv_2  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10672 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform -1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform -1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp 1688980957
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform -1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform -1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform -1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _039_
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1688980957
transform -1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform -1 0 6164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform -1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform -1 0 10672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform -1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp 1688980957
transform -1 0 12144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 1688980957
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1688980957
transform -1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1688980957
transform -1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform -1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1688980957
transform -1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1688980957
transform -1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1688980957
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform -1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _065_
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _066_
timestamp 1688980957
transform -1 0 5796 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _067_
timestamp 1688980957
transform -1 0 9016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _068_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _069_
timestamp 1688980957
transform 1 0 5704 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _070_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _071_
timestamp 1688980957
transform -1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform -1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform -1 0 11776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _085_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp 1688980957
transform 1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform -1 0 12420 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform -1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp 1688980957
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _090_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11316 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _091_
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _092_
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _093_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _093__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _094__44
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _094_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _095_
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _096_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _097_
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _098_
timestamp 1688980957
transform -1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _098__45
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _099_
timestamp 1688980957
transform 1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _100_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _101_
timestamp 1688980957
transform -1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _102_
timestamp 1688980957
transform -1 0 10212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _103__46
timestamp 1688980957
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _103_
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _104_
timestamp 1688980957
transform 1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _105_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_118
timestamp 1688980957
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_117
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_30
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_42
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 1688980957
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_42
timestamp 1688980957
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_46
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_91
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_103
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_117
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_10
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1688980957
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_74
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_89
timestamp 1688980957
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_107
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_111
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_116
timestamp 1688980957
transform 1 0 11776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_100
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_10
timestamp 1688980957
transform 1 0 2024 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_22
timestamp 1688980957
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_108
timestamp 1688980957
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_112
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_116
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_10
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_22
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_34
timestamp 1688980957
transform 1 0 4232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_46
timestamp 1688980957
transform 1 0 5336 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_94
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_117
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1688980957
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_104
timestamp 1688980957
transform 1 0 10672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_114
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_122
timestamp 1688980957
transform 1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_6
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_18
timestamp 1688980957
transform 1 0 2760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_30
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_42
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_103
timestamp 1688980957
transform 1 0 10580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_92
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_104
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_116
timestamp 1688980957
transform 1 0 11776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_124
timestamp 1688980957
transform 1 0 12512 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 1688980957
transform 1 0 9384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_13
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_20
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_24
timestamp 1688980957
transform 1 0 3312 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_49
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_54
timestamp 1688980957
transform 1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_57
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_63
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1688980957
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_96
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_106
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_119
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10304 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 4968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 10580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 11776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform -1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 2760 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform -1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 12880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 12880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 12880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 12880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 11408 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal3 s 13200 11160 14000 11280 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 13200 12248 14000 12368 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 2 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 3 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 4 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 5 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 6 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 7 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 8 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 9 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 10 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 11 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 12 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 13 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 14 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 15 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 16 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 17 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 18 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 19 nsew signal tristate
flabel metal2 s 2134 13200 2190 14000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 20 nsew signal input
flabel metal2 s 3330 13200 3386 14000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 21 nsew signal input
flabel metal2 s 4526 13200 4582 14000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 22 nsew signal input
flabel metal2 s 5722 13200 5778 14000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 23 nsew signal input
flabel metal2 s 6918 13200 6974 14000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 24 nsew signal input
flabel metal2 s 8114 13200 8170 14000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 25 nsew signal input
flabel metal2 s 9310 13200 9366 14000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 26 nsew signal input
flabel metal2 s 10506 13200 10562 14000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 27 nsew signal input
flabel metal2 s 11702 13200 11758 14000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 28 nsew signal input
flabel metal3 s 13200 1368 14000 1488 0 FreeSans 480 0 0 0 chany_top_out[0]
port 29 nsew signal tristate
flabel metal3 s 13200 2456 14000 2576 0 FreeSans 480 0 0 0 chany_top_out[1]
port 30 nsew signal tristate
flabel metal3 s 13200 3544 14000 3664 0 FreeSans 480 0 0 0 chany_top_out[2]
port 31 nsew signal tristate
flabel metal3 s 13200 4632 14000 4752 0 FreeSans 480 0 0 0 chany_top_out[3]
port 32 nsew signal tristate
flabel metal3 s 13200 5720 14000 5840 0 FreeSans 480 0 0 0 chany_top_out[4]
port 33 nsew signal tristate
flabel metal3 s 13200 6808 14000 6928 0 FreeSans 480 0 0 0 chany_top_out[5]
port 34 nsew signal tristate
flabel metal3 s 13200 7896 14000 8016 0 FreeSans 480 0 0 0 chany_top_out[6]
port 35 nsew signal tristate
flabel metal3 s 13200 8984 14000 9104 0 FreeSans 480 0 0 0 chany_top_out[7]
port 36 nsew signal tristate
flabel metal3 s 13200 10072 14000 10192 0 FreeSans 480 0 0 0 chany_top_out[8]
port 37 nsew signal tristate
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 prog_clk
port 38 nsew signal input
flabel metal3 s 13200 13336 14000 13456 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 39 nsew signal input
flabel metal3 s 13200 280 14000 400 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 40 nsew signal input
flabel metal2 s 12898 13200 12954 14000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 41 nsew signal input
flabel metal2 s 938 13200 994 14000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 42 nsew signal input
flabel metal4 s 2416 2128 2736 11472 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 5360 2128 5680 11472 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 8304 2128 8624 11472 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 11248 2128 11568 11472 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 3888 2128 4208 11472 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 6832 2128 7152 11472 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 9776 2128 10096 11472 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 12720 2128 13040 11472 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 6992 11424 6992 11424 0 vdd
rlabel via1 7072 10880 7072 10880 0 vss
rlabel metal1 10626 8534 10626 8534 0 _000_
rlabel metal1 9200 10030 9200 10030 0 _001_
rlabel metal1 11132 6766 11132 6766 0 _002_
rlabel metal1 8188 6766 8188 6766 0 _003_
rlabel metal1 1748 6290 1748 6290 0 _004_
rlabel metal1 6394 5202 6394 5202 0 _005_
rlabel metal1 11086 5712 11086 5712 0 _006_
rlabel metal1 9384 5678 9384 5678 0 _007_
rlabel metal1 11270 7922 11270 7922 0 _008_
rlabel metal1 10764 5882 10764 5882 0 _009_
rlabel metal1 9890 5780 9890 5780 0 _010_
rlabel metal1 11224 5814 11224 5814 0 _011_
rlabel metal1 7038 5338 7038 5338 0 _012_
rlabel metal1 2208 5746 2208 5746 0 _013_
rlabel metal1 2576 6222 2576 6222 0 _014_
rlabel metal1 5888 5270 5888 5270 0 _015_
rlabel metal1 8832 6970 8832 6970 0 _016_
rlabel metal1 12098 6732 12098 6732 0 _017_
rlabel metal1 11454 7378 11454 7378 0 _018_
rlabel metal1 9338 6698 9338 6698 0 _019_
rlabel metal1 9752 10234 9752 10234 0 _020_
rlabel metal1 10902 8602 10902 8602 0 _021_
rlabel metal1 10810 10710 10810 10710 0 _022_
rlabel metal1 9200 10778 9200 10778 0 _023_
rlabel metal2 12190 10931 12190 10931 0 ccff_head
rlabel metal2 12466 11815 12466 11815 0 ccff_tail
rlabel metal3 820 3604 820 3604 0 chanx_right_in[0]
rlabel metal3 820 4692 820 4692 0 chanx_right_in[1]
rlabel metal3 866 5780 866 5780 0 chanx_right_in[2]
rlabel metal3 1234 6868 1234 6868 0 chanx_right_in[3]
rlabel metal3 751 7956 751 7956 0 chanx_right_in[4]
rlabel metal3 820 9044 820 9044 0 chanx_right_in[5]
rlabel metal3 820 10132 820 10132 0 chanx_right_in[6]
rlabel metal3 843 11220 843 11220 0 chanx_right_in[7]
rlabel metal3 820 12308 820 12308 0 chanx_right_in[8]
rlabel metal2 782 1554 782 1554 0 chanx_right_out[0]
rlabel metal2 2162 959 2162 959 0 chanx_right_out[1]
rlabel metal2 3542 823 3542 823 0 chanx_right_out[2]
rlabel metal2 4922 823 4922 823 0 chanx_right_out[3]
rlabel metal2 6302 1520 6302 1520 0 chanx_right_out[4]
rlabel metal2 7682 1520 7682 1520 0 chanx_right_out[5]
rlabel metal2 9062 1520 9062 1520 0 chanx_right_out[6]
rlabel metal2 10442 823 10442 823 0 chanx_right_out[7]
rlabel metal2 11822 823 11822 823 0 chanx_right_out[8]
rlabel metal2 2714 12444 2714 12444 0 chany_top_in[0]
rlabel metal2 3358 12833 3358 12833 0 chany_top_in[1]
rlabel metal2 4554 12833 4554 12833 0 chany_top_in[2]
rlabel metal2 5750 12833 5750 12833 0 chany_top_in[3]
rlabel metal2 6946 12833 6946 12833 0 chany_top_in[4]
rlabel metal2 8142 12833 8142 12833 0 chany_top_in[5]
rlabel metal2 9384 11084 9384 11084 0 chany_top_in[6]
rlabel metal2 10534 12833 10534 12833 0 chany_top_in[7]
rlabel metal1 11868 11118 11868 11118 0 chany_top_in[8]
rlabel metal1 12006 2414 12006 2414 0 chany_top_out[0]
rlabel metal3 12842 2516 12842 2516 0 chany_top_out[1]
rlabel metal2 12466 3757 12466 3757 0 chany_top_out[2]
rlabel metal2 12466 4845 12466 4845 0 chany_top_out[3]
rlabel metal2 12466 5933 12466 5933 0 chany_top_out[4]
rlabel metal2 12282 7293 12282 7293 0 chany_top_out[5]
rlabel metal2 12374 8143 12374 8143 0 chany_top_out[6]
rlabel metal2 12466 9197 12466 9197 0 chany_top_out[7]
rlabel metal2 12466 10285 12466 10285 0 chany_top_out[8]
rlabel metal1 7774 7378 7774 7378 0 clknet_0_prog_clk
rlabel metal1 5750 6324 5750 6324 0 clknet_1_0__leaf_prog_clk
rlabel metal1 9108 7174 9108 7174 0 clknet_1_1__leaf_prog_clk
rlabel metal1 4692 6766 4692 6766 0 mem_right_track_0.DFF_0_.D
rlabel metal1 7452 6766 7452 6766 0 mem_right_track_0.DFF_0_.Q
rlabel metal1 7820 7514 7820 7514 0 mem_right_track_0.DFF_1_.Q
rlabel metal2 9154 8976 9154 8976 0 mem_right_track_2.DFF_0_.Q
rlabel metal1 10304 7854 10304 7854 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 10350 6290 10350 6290 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 1518 6256 1518 6256 0 mem_top_track_2.DFF_0_.Q
rlabel metal1 11592 7310 11592 7310 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 11868 3162 11868 3162 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 12466 7208 12466 7208 0 mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3450 2380 3450 2380 0 mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8970 11254 8970 11254 0 mux_right_track_2.INVTX1_0_.out
rlabel metal2 10166 10778 10166 10778 0 mux_right_track_2.INVTX1_1_.out
rlabel metal1 9568 10778 9568 10778 0 mux_right_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2990 2482 2990 2482 0 mux_right_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11224 7854 11224 7854 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 9522 5338 9522 5338 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 10580 6290 10580 6290 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 11546 6086 11546 6086 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 1978 6290 1978 6290 0 mux_top_track_2.INVTX1_0_.out
rlabel metal1 2254 5610 2254 5610 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 4232 5542 4232 5542 0 mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 7866 4556 7866 4556 0 mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9931 8534 9931 8534 0 net1
rlabel metal1 2346 11152 2346 11152 0 net10
rlabel metal1 2622 11047 2622 11047 0 net11
rlabel metal1 3496 11254 3496 11254 0 net12
rlabel metal2 4646 2587 4646 2587 0 net13
rlabel metal1 5980 3026 5980 3026 0 net14
rlabel metal2 7222 2587 7222 2587 0 net15
rlabel metal2 8602 2618 8602 2618 0 net16
rlabel metal1 10074 2414 10074 2414 0 net17
rlabel metal1 10948 2414 10948 2414 0 net18
rlabel metal2 11822 9418 11822 9418 0 net19
rlabel metal2 11822 5389 11822 5389 0 net2
rlabel metal1 11408 10438 11408 10438 0 net20
rlabel metal1 12144 3026 12144 3026 0 net21
rlabel metal1 11730 8466 11730 8466 0 net22
rlabel metal1 1886 11322 1886 11322 0 net23
rlabel metal1 11316 10642 11316 10642 0 net24
rlabel metal1 1932 2346 1932 2346 0 net25
rlabel metal1 2760 2346 2760 2346 0 net26
rlabel metal1 3726 2346 3726 2346 0 net27
rlabel metal1 5106 2312 5106 2312 0 net28
rlabel metal1 6302 2414 6302 2414 0 net29
rlabel metal1 2185 5338 2185 5338 0 net3
rlabel metal1 7636 2346 7636 2346 0 net30
rlabel metal1 8970 2346 8970 2346 0 net31
rlabel metal1 10626 2312 10626 2312 0 net32
rlabel metal1 12098 2346 12098 2346 0 net33
rlabel via1 11914 2363 11914 2363 0 net34
rlabel metal1 12190 3128 12190 3128 0 net35
rlabel metal2 1978 6528 1978 6528 0 net36
rlabel metal1 12236 5202 12236 5202 0 net37
rlabel metal1 12328 5882 12328 5882 0 net38
rlabel metal2 1886 7072 1886 7072 0 net39
rlabel metal1 1748 5678 1748 5678 0 net4
rlabel metal2 1794 9928 1794 9928 0 net40
rlabel metal1 12190 9554 12190 9554 0 net41
rlabel metal1 12236 9690 12236 9690 0 net42
rlabel metal1 11592 5746 11592 5746 0 net43
rlabel metal2 7222 5916 7222 5916 0 net44
rlabel metal1 10074 7514 10074 7514 0 net45
rlabel metal1 10810 9010 10810 9010 0 net46
rlabel metal1 8796 6290 8796 6290 0 net47
rlabel metal1 8606 8534 8606 8534 0 net48
rlabel metal1 5826 6698 5826 6698 0 net49
rlabel metal1 1886 6766 1886 6766 0 net5
rlabel metal1 9517 8942 9517 8942 0 net50
rlabel metal1 9517 6766 9517 6766 0 net51
rlabel metal2 7222 7174 7222 7174 0 net52
rlabel metal1 5581 6358 5581 6358 0 net53
rlabel metal1 9246 8534 9246 8534 0 net6
rlabel metal1 2185 9350 2185 9350 0 net7
rlabel metal1 1564 7378 1564 7378 0 net8
rlabel metal1 1610 10778 1610 10778 0 net9
rlabel metal3 2062 2516 2062 2516 0 prog_clk
rlabel metal3 12152 13396 12152 13396 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 12604 3502 12604 3502 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel via1 11178 11116 11178 11116 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 2254 11186 2254 11186 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
<< properties >>
string FIXED_BBOX 0 0 14000 14000
<< end >>
