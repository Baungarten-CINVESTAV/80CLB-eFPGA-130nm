* NGSPICE file created from cbx_1__10_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt cbx_1__10_ bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_ bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
+ bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ prog_clk top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_ vdd vss
XFILLER_0_13_40 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_062_ _012_ vss vss vdd vdd _040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_93 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_114_ mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net22 sky130_fd_sc_hd__inv_2
Xoutput31 net31 vss vss vdd vdd chanx_left_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 vss vss vdd vdd top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 vss vss vdd vdd bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_85 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_29 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_113_ net13 vss vss vdd vdd mux_top_ipin_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_061_ mem_top_ipin_1.DFF_1_.Q vss vss vdd vdd _012_ sky130_fd_sc_hd__clkbuf_1
Xoutput32 net32 vss vss vdd vdd chanx_left_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 vss vss vdd vdd bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_20 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_11_6 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_40 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_060_ _011_ vss vss vdd vdd _041_ sky130_fd_sc_hd__clkbuf_1
X_112_ net4 vss vss vdd vdd mux_top_ipin_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_1_52 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput22 net22 vss vss vdd vdd bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
+ sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 vss vss vdd vdd chanx_right_out[0] sky130_fd_sc_hd__clkbuf_4
X_111_ mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net21 sky130_fd_sc_hd__inv_2
Xoutput23 net23 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__clkbuf_4
Xoutput34 net34 vss vss vdd vdd chanx_right_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_66 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_13_33 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_10_56 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_110_ net16 vss vss vdd vdd mux_top_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
Xoutput24 net24 vss vss vdd vdd chanx_left_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 vss vss vdd vdd chanx_right_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_169_ mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out _035_ vss vss vdd vdd mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_13_79 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_46 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput25 net25 vss vss vdd vdd chanx_left_out[1] sky130_fd_sc_hd__clkbuf_4
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput36 net36 vss vss vdd vdd chanx_right_out[3] sky130_fd_sc_hd__clkbuf_4
X_099_ mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net42 sky130_fd_sc_hd__inv_2
X_168_ mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out _034_ vss vss vdd vdd mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
Xoutput26 net26 vss vss vdd vdd chanx_left_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput37 net37 vss vss vdd vdd chanx_right_out[4] sky130_fd_sc_hd__clkbuf_4
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_098_ _008_ vss vss vdd vdd _016_ sky130_fd_sc_hd__clkbuf_1
X_167_ mux_bottom_ipin_0.INVTX1_1_.out _033_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xoutput27 net27 vss vss vdd vdd chanx_left_out[3] sky130_fd_sc_hd__clkbuf_4
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput38 net38 vss vss vdd vdd chanx_right_out[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_097_ mem_bottom_ipin_0.DFF_1_.Q vss vss vdd vdd _008_ sky130_fd_sc_hd__clkbuf_1
X_166_ mux_top_ipin_0.INVTX1_3_.out _032_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xoutput28 net28 vss vss vdd vdd chanx_left_out[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput39 net39 vss vss vdd vdd chanx_right_out[6] sky130_fd_sc_hd__clkbuf_4
X_149_ net2 vss vss vdd vdd net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_46 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_11_82 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_165_ mux_top_ipin_0.INVTX1_5_.out _031_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_096_ _007_ vss vss vdd vdd _017_ sky130_fd_sc_hd__clkbuf_1
X_148_ net3 vss vss vdd vdd net34 sky130_fd_sc_hd__clkbuf_1
Xoutput29 net29 vss vss vdd vdd chanx_left_out[5] sky130_fd_sc_hd__clkbuf_4
X_079_ mem_top_ipin_0.DFF_1_.Q vss vss vdd vdd _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_91 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_181_ mux_top_ipin_2.INVTX1_0_.out _047_ vss vss vdd vdd mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_095_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _007_ sky130_fd_sc_hd__clkbuf_1
X_164_ mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out _030_ vss vss vdd vdd mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_078_ _001_ vss vss vdd vdd _031_ sky130_fd_sc_hd__clkbuf_1
X_147_ net4 vss vss vdd vdd net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_29 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_180_ mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out _046_ vss vss vdd vdd mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_094_ _006_ vss vss vdd vdd _020_ sky130_fd_sc_hd__clkbuf_1
X_163_ net44 _029_ vss vss vdd vdd mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_077_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _001_ sky130_fd_sc_hd__clkbuf_1
X_146_ net5 vss vss vdd vdd net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_6 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_093_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _006_ sky130_fd_sc_hd__clkbuf_1
X_162_ mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out _028_ vss vss vdd vdd mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
Xinput1 ccff_head vss vss vdd vdd net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_74 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_11_30 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_145_ net6 vss vss vdd vdd net37 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
X_076_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _037_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_28 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_059_ mem_top_ipin_1.DFF_0_.Q vss vss vdd vdd _011_ sky130_fd_sc_hd__clkbuf_1
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_71 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_42 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_161_ mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out _027_ vss vss vdd vdd mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_092_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _024_ sky130_fd_sc_hd__inv_2
Xinput2 chanx_left_in[0] vss vss vdd vdd net2 sky130_fd_sc_hd__buf_1
X_144_ net7 vss vss vdd vdd net38 sky130_fd_sc_hd__clkbuf_1
X_127_ clknet_1_1__leaf_prog_clk net51 vss vss vdd vdd mem_top_ipin_2.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_075_ mem_top_ipin_0.DFF_1_.Q vss vss vdd vdd _035_ sky130_fd_sc_hd__inv_2
X_058_ mem_top_ipin_1.DFF_0_.Q vss vss vdd vdd _043_ sky130_fd_sc_hd__inv_2
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_5_40 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_143_ net8 vss vss vdd vdd net39 sky130_fd_sc_hd__clkbuf_1
X_160_ mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out _026_ vss vss vdd vdd mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_091_ mem_bottom_ipin_0.DFF_1_.Q vss vss vdd vdd _026_ sky130_fd_sc_hd__inv_2
X_074_ _000_ vss vss vdd vdd _028_ sky130_fd_sc_hd__clkbuf_1
Xinput3 chanx_left_in[1] vss vss vdd vdd net3 sky130_fd_sc_hd__buf_1
X_126_ clknet_1_1__leaf_prog_clk net49 vss vss vdd vdd net23 sky130_fd_sc_hd__dfxtp_1
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_057_ mem_top_ipin_1.DFF_1_.Q vss vss vdd vdd _042_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_109_ net3 vss vss vdd vdd mux_top_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_0_11_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_090_ _005_ vss vss vdd vdd _018_ sky130_fd_sc_hd__clkbuf_1
Xinput4 chanx_left_in[2] vss vss vdd vdd net4 sky130_fd_sc_hd__buf_1
XFILLER_0_1_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_142_ net9 vss vss vdd vdd net40 sky130_fd_sc_hd__clkbuf_1
X_056_ _010_ vss vss vdd vdd _044_ sky130_fd_sc_hd__buf_1
X_125_ clknet_1_1__leaf_prog_clk net47 vss vss vdd vdd mem_top_ipin_1.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
X_073_ mem_top_ipin_0.DFF_2_.Q vss vss vdd vdd _000_ sky130_fd_sc_hd__clkbuf_1
X_108_ net12 vss vss vdd vdd mux_top_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_163__44 vss vss vdd vdd net44 _163__44/LO sky130_fd_sc_hd__conb_1
XTAP_50 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 chanx_left_in[3] vss vss vdd vdd net5 sky130_fd_sc_hd__buf_1
X_141_ net10 vss vss vdd vdd net41 sky130_fd_sc_hd__clkbuf_1
X_072_ _015_ vss vss vdd vdd _032_ sky130_fd_sc_hd__clkbuf_1
X_055_ net23 vss vss vdd vdd _010_ sky130_fd_sc_hd__clkbuf_1
X_124_ clknet_1_1__leaf_prog_clk net50 vss vss vdd vdd mem_top_ipin_1.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_107_ net7 vss vss vdd vdd mux_top_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_21 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_51 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 chanx_left_in[4] vss vss vdd vdd net6 sky130_fd_sc_hd__buf_1
X_071_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _015_ sky130_fd_sc_hd__clkbuf_1
XTAP_40 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_11 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_140_ net11 vss vss vdd vdd net24 sky130_fd_sc_hd__buf_1
X_054_ _009_ vss vss vdd vdd _045_ sky130_fd_sc_hd__clkbuf_1
X_123_ clknet_1_0__leaf_prog_clk net48 vss vss vdd vdd mem_top_ipin_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
X_106_ mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out vss vss vdd vdd net20 sky130_fd_sc_hd__inv_2
XFILLER_0_3_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_47 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xinput7 chanx_left_in[5] vss vss vdd vdd net7 sky130_fd_sc_hd__buf_1
XFILLER_0_10_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_41 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _038_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_77 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_11 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_30 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 chanx_left_in[8] vss vss vdd vdd net10 sky130_fd_sc_hd__buf_1
X_053_ mem_top_ipin_2.DFF_0_.Q vss vss vdd vdd _009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_56 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_122_ clknet_1_0__leaf_prog_clk net54 vss vss vdd vdd mem_top_ipin_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
X_105_ net19 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_0_8_22 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xinput8 chanx_left_in[6] vss vss vdd vdd net8 sky130_fd_sc_hd__clkbuf_1
XTAP_42 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_31 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_052_ mem_top_ipin_2.DFF_0_.Q vss vss vdd vdd _047_ sky130_fd_sc_hd__inv_2
X_104_ net11 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_121_ clknet_1_0__leaf_prog_clk net55 vss vss vdd vdd mem_top_ipin_0.DFF_2_.Q sky130_fd_sc_hd__dfxtp_1
Xinput11 chanx_right_in[0] vss vss vdd vdd net11 sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput9 chanx_left_in[7] vss vss vdd vdd net9 sky130_fd_sc_hd__clkbuf_1
XTAP_43 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_8 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_32 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_81 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput12 chanx_right_in[1] vss vss vdd vdd net12 sky130_fd_sc_hd__buf_1
X_120_ clknet_1_1__leaf_prog_clk net1 vss vss vdd vdd mem_bottom_ipin_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_103_ net2 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_12_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold1 mem_top_ipin_0.DFF_2_.Q vss vss vdd vdd net47 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_44 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_15 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_33 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ net6 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
Xinput13 chanx_right_in[2] vss vss vdd vdd net13 sky130_fd_sc_hd__buf_1
X_179_ mux_top_ipin_2.INVTX1_1_.out _045_ vss vss vdd vdd mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold2 mem_bottom_ipin_0.DFF_2_.Q vss vss vdd vdd net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_18 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_45 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_34 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_91 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput14 chanx_right_in[3] vss vss vdd vdd net14 sky130_fd_sc_hd__buf_1
X_101_ net15 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_0_8_59 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_178_ net46 _044_ vss vss vdd vdd mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_150__43 vss vss vdd vdd net43 _150__43/LO sky130_fd_sc_hd__conb_1
Xhold3 mem_top_ipin_2.DFF_0_.Q vss vss vdd vdd net49 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_46 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_40 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_178__46 vss vss vdd vdd net46 _178__46/LO sky130_fd_sc_hd__conb_1
X_100_ net10 vss vss vdd vdd mux_bottom_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
Xinput15 chanx_right_in[4] vss vss vdd vdd net15 sky130_fd_sc_hd__buf_1
X_177_ mux_top_ipin_1.INVTX1_0_.out _043_ vss vss vdd vdd mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold4 mem_top_ipin_1.DFF_0_.Q vss vss vdd vdd net50 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_47 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_52 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput16 chanx_right_in[5] vss vss vdd vdd net16 sky130_fd_sc_hd__buf_1
X_159_ mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out _025_ vss vss vdd vdd mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_176_ mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out _042_ vss vss vdd vdd mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_3_83 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold5 mem_top_ipin_1.DFF_1_.Q vss vss vdd vdd net51 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_48 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XTAP_37 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput17 chanx_right_in[6] vss vss vdd vdd net17 sky130_fd_sc_hd__clkbuf_1
X_175_ mux_top_ipin_1.INVTX1_1_.out _041_ vss vss vdd vdd mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_158_ mux_bottom_ipin_0.INVTX1_4_.out _024_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
Xhold6 mem_bottom_ipin_0.DFF_1_.Q vss vss vdd vdd net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_089_ mem_bottom_ipin_0.DFF_2_.Q vss vss vdd vdd _005_ sky130_fd_sc_hd__clkbuf_1
XTAP_49 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput18 chanx_right_in[7] vss vss vdd vdd net18 sky130_fd_sc_hd__clkbuf_1
X_088_ _004_ vss vss vdd vdd _019_ sky130_fd_sc_hd__clkbuf_1
X_157_ mux_bottom_ipin_0.INVTX1_2_.out _023_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_174_ net45 _040_ vss vss vdd vdd mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
XFILLER_0_3_74 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_8 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xhold7 mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd net53 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_39 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_28 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 chanx_right_in[8] vss vss vdd vdd net19 sky130_fd_sc_hd__buf_1
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_173_ mux_bottom_ipin_0.INVTX1_0_.out _039_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_087_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _004_ sky130_fd_sc_hd__clkbuf_1
Xhold8 mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd net54 sky130_fd_sc_hd__dlygate4sd3_1
X_156_ mux_bottom_ipin_0.INVTX1_0_.out _022_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_139_ net12 vss vss vdd vdd net25 sky130_fd_sc_hd__clkbuf_1
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XTAP_29 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out _021_ vss vss vdd vdd mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_086_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _023_ sky130_fd_sc_hd__inv_2
X_172_ mux_top_ipin_0.INVTX1_2_.out _038_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_069_ _014_ vss vss vdd vdd _030_ sky130_fd_sc_hd__clkbuf_1
X_138_ net13 vss vss vdd vdd net26 sky130_fd_sc_hd__clkbuf_1
Xhold9 mem_top_ipin_0.DFF_1_.Q vss vss vdd vdd net55 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_13 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_171_ mux_top_ipin_0.INVTX1_4_.out _037_ vss vss vdd vdd mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_154_ mux_bottom_ipin_0.INVTX1_5_.out _020_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_085_ _003_ vss vss vdd vdd _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_137_ net14 vss vss vdd vdd net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_98 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_21 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_068_ mem_top_ipin_0.DFF_1_.Q vss vss vdd vdd _014_ sky130_fd_sc_hd__clkbuf_1
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_174__45 vss vss vdd vdd net45 _174__45/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3_12 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_170_ mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out _036_ vss vss vdd vdd mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_136_ net15 vss vss vdd vdd net28 sky130_fd_sc_hd__clkbuf_1
X_153_ mux_bottom_ipin_0.INVTX1_3_.out _019_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_9_55 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_33 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_084_ mem_bottom_ipin_0.DFF_1_.Q vss vss vdd vdd _003_ sky130_fd_sc_hd__clkbuf_1
X_067_ _013_ vss vss vdd vdd _033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_119_ clknet_1_0__leaf_prog_clk net53 vss vss vdd vdd mem_bottom_ipin_0.DFF_1_.Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_45 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_101 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_152_ mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out _018_ vss vss vdd vdd mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_083_ mem_bottom_ipin_0.DFF_0_.Q vss vss vdd vdd _022_ sky130_fd_sc_hd__inv_2
X_118_ clknet_1_1__leaf_prog_clk net52 vss vss vdd vdd mem_bottom_ipin_0.DFF_2_.Q
+ sky130_fd_sc_hd__dfxtp_1
X_135_ net16 vss vss vdd vdd net29 sky130_fd_sc_hd__clkbuf_1
X_066_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _013_ sky130_fd_sc_hd__clkbuf_1
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XANTENNA_1 net45 vss vss vdd vdd sky130_fd_sc_hd__diode_2
XFILLER_0_13_92 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_134_ net17 vss vss vdd vdd net30 sky130_fd_sc_hd__clkbuf_1
X_082_ mem_bottom_ipin_0.DFF_1_.Q vss vss vdd vdd _025_ sky130_fd_sc_hd__inv_2
X_151_ mux_bottom_ipin_0.INVTX1_1_.out _017_ vss vss vdd vdd mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_065_ mem_top_ipin_0.DFF_0_.Q vss vss vdd vdd _039_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_117_ net23 vss vss vdd vdd _046_ sky130_fd_sc_hd__inv_2
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XANTENNA_2 net45 vss vss vdd vdd sky130_fd_sc_hd__diode_2
X_150_ net43 _016_ vss vss vdd vdd mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out sky130_fd_sc_hd__ebufn_1
X_081_ mem_bottom_ipin_0.DFF_2_.Q vss vss vdd vdd _027_ sky130_fd_sc_hd__inv_2
X_133_ net18 vss vss vdd vdd net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_50 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_064_ mem_top_ipin_0.DFF_1_.Q vss vss vdd vdd _036_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_6 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XANTENNA_3 chanx_right_in[4] vss vss vdd vdd sky130_fd_sc_hd__diode_2
X_116_ net14 vss vss vdd vdd mux_top_ipin_2.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_4_9 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xoutput40 net40 vss vss vdd vdd chanx_right_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_72 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_132_ net19 vss vss vdd vdd net32 sky130_fd_sc_hd__clkbuf_1
X_063_ mem_top_ipin_0.DFF_2_.Q vss vss vdd vdd _034_ sky130_fd_sc_hd__inv_2
X_080_ _002_ vss vss vdd vdd _029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_115_ net5 vss vss vdd vdd mux_top_ipin_2.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_0_39 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput30 net30 vss vss vdd vdd chanx_left_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_102 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput41 net41 vss vss vdd vdd chanx_right_out[8] sky130_fd_sc_hd__clkbuf_4
.ends

