magic
tech sky130A
magscale 1 2
timestamp 1708041323
<< obsli1 >>
rect 1104 2159 14812 17425
<< obsm1 >>
rect 474 2128 15074 17808
<< metal2 >>
rect 938 19200 994 20000
rect 1674 19200 1730 20000
rect 2410 19200 2466 20000
rect 3146 19200 3202 20000
rect 3882 19200 3938 20000
rect 4618 19200 4674 20000
rect 5354 19200 5410 20000
rect 6090 19200 6146 20000
rect 6826 19200 6882 20000
rect 7562 19200 7618 20000
rect 8298 19200 8354 20000
rect 9034 19200 9090 20000
rect 9770 19200 9826 20000
rect 10506 19200 10562 20000
rect 11242 19200 11298 20000
rect 11978 19200 12034 20000
rect 12714 19200 12770 20000
rect 13450 19200 13506 20000
rect 14186 19200 14242 20000
rect 14922 19200 14978 20000
rect 478 0 534 800
rect 1306 0 1362 800
rect 2134 0 2190 800
rect 2962 0 3018 800
rect 3790 0 3846 800
rect 4618 0 4674 800
rect 5446 0 5502 800
rect 6274 0 6330 800
rect 7102 0 7158 800
rect 7930 0 7986 800
rect 8758 0 8814 800
rect 9586 0 9642 800
rect 10414 0 10470 800
rect 11242 0 11298 800
rect 12070 0 12126 800
rect 12898 0 12954 800
rect 13726 0 13782 800
rect 14554 0 14610 800
<< obsm2 >>
rect 480 19144 882 19200
rect 1050 19144 1618 19200
rect 1786 19144 2354 19200
rect 2522 19144 3090 19200
rect 3258 19144 3826 19200
rect 3994 19144 4562 19200
rect 4730 19144 5298 19200
rect 5466 19144 6034 19200
rect 6202 19144 6770 19200
rect 6938 19144 7506 19200
rect 7674 19144 8242 19200
rect 8410 19144 8978 19200
rect 9146 19144 9714 19200
rect 9882 19144 10450 19200
rect 10618 19144 11186 19200
rect 11354 19144 11922 19200
rect 12090 19144 12658 19200
rect 12826 19144 13394 19200
rect 13562 19144 14130 19200
rect 14298 19144 14866 19200
rect 15034 19144 15070 19200
rect 480 856 15070 19144
rect 590 734 1250 856
rect 1418 734 2078 856
rect 2246 734 2906 856
rect 3074 734 3734 856
rect 3902 734 4562 856
rect 4730 734 5390 856
rect 5558 734 6218 856
rect 6386 734 7046 856
rect 7214 734 7874 856
rect 8042 734 8702 856
rect 8870 734 9530 856
rect 9698 734 10358 856
rect 10526 734 11186 856
rect 11354 734 12014 856
rect 12182 734 12842 856
rect 13010 734 13670 856
rect 13838 734 14498 856
rect 14666 734 15070 856
<< metal3 >>
rect 0 17960 800 18080
rect 15200 17960 16000 18080
rect 0 16600 800 16720
rect 15200 16600 16000 16720
rect 0 15240 800 15360
rect 15200 15240 16000 15360
rect 0 13880 800 14000
rect 15200 13880 16000 14000
rect 0 12520 800 12640
rect 15200 12520 16000 12640
rect 0 11160 800 11280
rect 15200 11160 16000 11280
rect 0 9800 800 9920
rect 15200 9800 16000 9920
rect 0 8440 800 8560
rect 15200 8440 16000 8560
rect 0 7080 800 7200
rect 15200 7080 16000 7200
rect 0 5720 800 5840
rect 15200 5720 16000 5840
rect 0 4360 800 4480
rect 15200 4360 16000 4480
rect 0 3000 800 3120
rect 15200 3000 16000 3120
rect 15200 1640 16000 1760
<< obsm3 >>
rect 880 17880 15120 18053
rect 798 16800 15210 17880
rect 880 16520 15120 16800
rect 798 15440 15210 16520
rect 880 15160 15120 15440
rect 798 14080 15210 15160
rect 880 13800 15120 14080
rect 798 12720 15210 13800
rect 880 12440 15120 12720
rect 798 11360 15210 12440
rect 880 11080 15120 11360
rect 798 10000 15210 11080
rect 880 9720 15120 10000
rect 798 8640 15210 9720
rect 880 8360 15120 8640
rect 798 7280 15210 8360
rect 880 7000 15120 7280
rect 798 5920 15210 7000
rect 880 5640 15120 5920
rect 798 4560 15210 5640
rect 880 4280 15120 4560
rect 798 3200 15210 4280
rect 880 2920 15120 3200
rect 798 1840 15210 2920
rect 798 1667 15120 1840
<< metal4 >>
rect 2657 2128 2977 17456
rect 4370 2128 4690 17456
rect 6084 2128 6404 17456
rect 7797 2128 8117 17456
rect 9511 2128 9831 17456
rect 11224 2128 11544 17456
rect 12938 2128 13258 17456
rect 14651 2128 14971 17456
<< labels >>
rlabel metal3 s 15200 3000 16000 3120 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 15200 4360 16000 4480 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 chanx_left_in[0]
port 3 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 4 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[2]
port 5 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[3]
port 6 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[4]
port 7 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[5]
port 8 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[6]
port 9 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[7]
port 10 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[8]
port 11 nsew signal input
rlabel metal2 s 478 0 534 800 6 chanx_left_out[0]
port 12 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 chanx_left_out[1]
port 13 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 chanx_left_out[2]
port 14 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 chanx_left_out[3]
port 15 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 chanx_left_out[4]
port 16 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 chanx_left_out[5]
port 17 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 chanx_left_out[6]
port 18 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 chanx_left_out[7]
port 19 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 chanx_left_out[8]
port 20 nsew signal output
rlabel metal3 s 15200 5720 16000 5840 6 chanx_right_in[0]
port 21 nsew signal input
rlabel metal3 s 15200 7080 16000 7200 6 chanx_right_in[1]
port 22 nsew signal input
rlabel metal3 s 15200 8440 16000 8560 6 chanx_right_in[2]
port 23 nsew signal input
rlabel metal3 s 15200 9800 16000 9920 6 chanx_right_in[3]
port 24 nsew signal input
rlabel metal3 s 15200 11160 16000 11280 6 chanx_right_in[4]
port 25 nsew signal input
rlabel metal3 s 15200 12520 16000 12640 6 chanx_right_in[5]
port 26 nsew signal input
rlabel metal3 s 15200 13880 16000 14000 6 chanx_right_in[6]
port 27 nsew signal input
rlabel metal3 s 15200 15240 16000 15360 6 chanx_right_in[7]
port 28 nsew signal input
rlabel metal3 s 15200 16600 16000 16720 6 chanx_right_in[8]
port 29 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 chanx_right_out[0]
port 30 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 chanx_right_out[1]
port 31 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 chanx_right_out[2]
port 32 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 chanx_right_out[3]
port 33 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 chanx_right_out[4]
port 34 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 chanx_right_out[5]
port 35 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 chanx_right_out[6]
port 36 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 chanx_right_out[7]
port 37 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chanx_right_out[8]
port 38 nsew signal output
rlabel metal2 s 1674 19200 1730 20000 6 chany_top_in[0]
port 39 nsew signal input
rlabel metal2 s 2410 19200 2466 20000 6 chany_top_in[1]
port 40 nsew signal input
rlabel metal2 s 3146 19200 3202 20000 6 chany_top_in[2]
port 41 nsew signal input
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_in[3]
port 42 nsew signal input
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_in[4]
port 43 nsew signal input
rlabel metal2 s 5354 19200 5410 20000 6 chany_top_in[5]
port 44 nsew signal input
rlabel metal2 s 6090 19200 6146 20000 6 chany_top_in[6]
port 45 nsew signal input
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_in[7]
port 46 nsew signal input
rlabel metal2 s 7562 19200 7618 20000 6 chany_top_in[8]
port 47 nsew signal input
rlabel metal2 s 9034 19200 9090 20000 6 chany_top_out[0]
port 48 nsew signal output
rlabel metal2 s 9770 19200 9826 20000 6 chany_top_out[1]
port 49 nsew signal output
rlabel metal2 s 10506 19200 10562 20000 6 chany_top_out[2]
port 50 nsew signal output
rlabel metal2 s 11242 19200 11298 20000 6 chany_top_out[3]
port 51 nsew signal output
rlabel metal2 s 11978 19200 12034 20000 6 chany_top_out[4]
port 52 nsew signal output
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_out[5]
port 53 nsew signal output
rlabel metal2 s 13450 19200 13506 20000 6 chany_top_out[6]
port 54 nsew signal output
rlabel metal2 s 14186 19200 14242 20000 6 chany_top_out[7]
port 55 nsew signal output
rlabel metal2 s 14922 19200 14978 20000 6 chany_top_out[8]
port 56 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 57 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 58 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 prog_clk
port 59 nsew signal input
rlabel metal3 s 15200 1640 16000 1760 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 60 nsew signal input
rlabel metal3 s 15200 17960 16000 18080 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 61 nsew signal input
rlabel metal2 s 938 19200 994 20000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 62 nsew signal input
rlabel metal2 s 8298 19200 8354 20000 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 63 nsew signal input
rlabel metal4 s 2657 2128 2977 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 17456 6 vdd
port 64 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 17456 6 vss
port 65 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 17456 6 vss
port 65 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 879826
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_1__0_/runs/24_02_15_17_54/results/signoff/sb_1__0_.magic.gds
string GDS_START 114998
<< end >>

