magic
tech sky130A
magscale 1 2
timestamp 1708121277
<< viali >>
rect 23673 27625 23707 27659
rect 3893 27557 3927 27591
rect 6009 27557 6043 27591
rect 6561 27557 6595 27591
rect 9413 27557 9447 27591
rect 12173 27557 12207 27591
rect 14197 27557 14231 27591
rect 19809 27557 19843 27591
rect 26525 27557 26559 27591
rect 4353 27489 4387 27523
rect 7113 27489 7147 27523
rect 9137 27489 9171 27523
rect 12357 27489 12391 27523
rect 16865 27489 16899 27523
rect 20913 27489 20947 27523
rect 4077 27421 4111 27455
rect 4261 27421 4295 27455
rect 4537 27421 4571 27455
rect 5641 27421 5675 27455
rect 5917 27421 5951 27455
rect 6193 27421 6227 27455
rect 6745 27421 6779 27455
rect 7021 27421 7055 27455
rect 7297 27421 7331 27455
rect 8033 27421 8067 27455
rect 8309 27421 8343 27455
rect 8585 27421 8619 27455
rect 9597 27421 9631 27455
rect 9689 27421 9723 27455
rect 10057 27421 10091 27455
rect 10333 27421 10367 27455
rect 10517 27421 10551 27455
rect 11253 27421 11287 27455
rect 11713 27421 11747 27455
rect 11989 27421 12023 27455
rect 12081 27421 12115 27455
rect 12541 27421 12575 27455
rect 13185 27421 13219 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 14749 27421 14783 27455
rect 15761 27421 15795 27455
rect 17509 27421 17543 27455
rect 17785 27421 17819 27455
rect 18337 27421 18371 27455
rect 19257 27421 19291 27455
rect 19557 27421 19591 27455
rect 19993 27421 20027 27455
rect 20177 27421 20211 27455
rect 21097 27421 21131 27455
rect 22385 27421 22419 27455
rect 23397 27421 23431 27455
rect 23857 27421 23891 27455
rect 23949 27421 23983 27455
rect 26065 27421 26099 27455
rect 28273 27421 28307 27455
rect 1501 27353 1535 27387
rect 17601 27353 17635 27387
rect 23489 27353 23523 27387
rect 26341 27353 26375 27387
rect 1593 27285 1627 27319
rect 4629 27285 4663 27319
rect 4905 27285 4939 27319
rect 5457 27285 5491 27319
rect 5733 27285 5767 27319
rect 6837 27285 6871 27319
rect 7757 27285 7791 27319
rect 8125 27285 8159 27319
rect 8401 27285 8435 27319
rect 8677 27285 8711 27319
rect 9781 27285 9815 27319
rect 10149 27285 10183 27319
rect 10977 27285 11011 27319
rect 11069 27285 11103 27319
rect 11529 27285 11563 27319
rect 11805 27285 11839 27319
rect 13001 27285 13035 27319
rect 13737 27285 13771 27319
rect 14565 27285 14599 27319
rect 15393 27285 15427 27319
rect 16313 27285 16347 27319
rect 17417 27285 17451 27319
rect 17877 27285 17911 27319
rect 18889 27285 18923 27319
rect 19349 27285 19383 27319
rect 19625 27285 19659 27319
rect 20821 27285 20855 27319
rect 21557 27285 21591 27319
rect 22201 27285 22235 27319
rect 25881 27285 25915 27319
rect 28457 27285 28491 27319
rect 1685 27081 1719 27115
rect 8033 27081 8067 27115
rect 10609 27081 10643 27115
rect 11529 27081 11563 27115
rect 12909 27081 12943 27115
rect 14657 27081 14691 27115
rect 16497 27081 16531 27115
rect 18061 27081 18095 27115
rect 19533 27081 19567 27115
rect 21005 27081 21039 27115
rect 21281 27081 21315 27115
rect 21833 27081 21867 27115
rect 25421 27081 25455 27115
rect 2605 27013 2639 27047
rect 2697 27013 2731 27047
rect 4261 27013 4295 27047
rect 11989 27013 12023 27047
rect 13544 27013 13578 27047
rect 18420 27013 18454 27047
rect 19892 27013 19926 27047
rect 1593 26945 1627 26979
rect 2421 26945 2455 26979
rect 3341 26945 3375 26979
rect 4905 26945 4939 26979
rect 5089 26945 5123 26979
rect 5917 26945 5951 26979
rect 6009 26945 6043 26979
rect 6101 26945 6135 26979
rect 7481 26945 7515 26979
rect 8217 26945 8251 26979
rect 8309 26945 8343 26979
rect 8953 26945 8987 26979
rect 9873 26945 9907 26979
rect 10149 26945 10183 26979
rect 10701 26945 10735 26979
rect 11713 26945 11747 26979
rect 12817 26945 12851 26979
rect 13093 26945 13127 26979
rect 14749 26945 14783 26979
rect 15117 26945 15151 26979
rect 15384 26945 15418 26979
rect 16948 26945 16982 26979
rect 18153 26945 18187 26979
rect 21097 26945 21131 26979
rect 21465 26945 21499 26979
rect 21993 26945 22027 26979
rect 22101 26945 22135 26979
rect 22201 26945 22235 26979
rect 22661 26945 22695 26979
rect 23397 26945 23431 26979
rect 24685 26945 24719 26979
rect 25605 26945 25639 26979
rect 25881 26945 25915 26979
rect 25973 26945 26007 26979
rect 26341 26945 26375 26979
rect 27169 26945 27203 26979
rect 27905 26945 27939 26979
rect 28549 26945 28583 26979
rect 3525 26877 3559 26911
rect 4169 26877 4203 26911
rect 6377 26877 6411 26911
rect 6561 26877 6595 26911
rect 7297 26877 7331 26911
rect 8769 26877 8803 26911
rect 9965 26877 9999 26911
rect 10885 26877 10919 26911
rect 11345 26877 11379 26911
rect 11897 26877 11931 26911
rect 13277 26877 13311 26911
rect 16681 26877 16715 26911
rect 19625 26877 19659 26911
rect 22477 26877 22511 26911
rect 23213 26877 23247 26911
rect 23949 26877 23983 26911
rect 24133 26877 24167 26911
rect 24869 26877 24903 26911
rect 26157 26877 26191 26911
rect 26985 26877 27019 26911
rect 27997 26877 28031 26911
rect 3157 26809 3191 26843
rect 3709 26809 3743 26843
rect 4721 26809 4755 26843
rect 5273 26809 5307 26843
rect 5733 26809 5767 26843
rect 7665 26809 7699 26843
rect 12449 26809 12483 26843
rect 12633 26809 12667 26843
rect 23121 26809 23155 26843
rect 23581 26809 23615 26843
rect 2237 26741 2271 26775
rect 6745 26741 6779 26775
rect 8401 26741 8435 26775
rect 9413 26741 9447 26775
rect 9689 26741 9723 26775
rect 14841 26741 14875 26775
rect 21557 26741 21591 26775
rect 24317 26741 24351 26775
rect 25053 26741 25087 26775
rect 26801 26741 26835 26775
rect 27353 26741 27387 26775
rect 27721 26741 27755 26775
rect 28365 26741 28399 26775
rect 2881 26537 2915 26571
rect 3341 26537 3375 26571
rect 4629 26537 4663 26571
rect 7665 26537 7699 26571
rect 9413 26537 9447 26571
rect 11437 26537 11471 26571
rect 13921 26537 13955 26571
rect 15853 26537 15887 26571
rect 18981 26537 19015 26571
rect 20269 26537 20303 26571
rect 21281 26537 21315 26571
rect 23857 26537 23891 26571
rect 28181 26537 28215 26571
rect 5181 26469 5215 26503
rect 7941 26469 7975 26503
rect 12173 26469 12207 26503
rect 16129 26469 16163 26503
rect 17049 26469 17083 26503
rect 17509 26469 17543 26503
rect 19993 26469 20027 26503
rect 23305 26469 23339 26503
rect 24685 26469 24719 26503
rect 28365 26469 28399 26503
rect 5549 26401 5583 26435
rect 6193 26401 6227 26435
rect 6929 26401 6963 26435
rect 7113 26401 7147 26435
rect 9137 26401 9171 26435
rect 9781 26401 9815 26435
rect 9965 26401 9999 26435
rect 14473 26401 14507 26435
rect 16405 26401 16439 26435
rect 16589 26401 16623 26435
rect 17141 26401 17175 26435
rect 18705 26401 18739 26435
rect 19441 26401 19475 26435
rect 20637 26401 20671 26435
rect 20821 26401 20855 26435
rect 21833 26401 21867 26435
rect 22477 26401 22511 26435
rect 25421 26401 25455 26435
rect 26617 26401 26651 26435
rect 27353 26401 27387 26435
rect 27537 26401 27571 26435
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 4537 26333 4571 26367
rect 4813 26333 4847 26367
rect 5365 26333 5399 26367
rect 6561 26333 6595 26367
rect 6837 26333 6871 26367
rect 7573 26333 7607 26367
rect 7849 26333 7883 26367
rect 8125 26333 8159 26367
rect 8493 26333 8527 26367
rect 8769 26333 8803 26367
rect 8953 26333 8987 26367
rect 10517 26333 10551 26367
rect 11253 26333 11287 26367
rect 12541 26333 12575 26367
rect 14197 26333 14231 26367
rect 14740 26333 14774 26367
rect 16313 26333 16347 26367
rect 17325 26333 17359 26367
rect 17877 26333 17911 26367
rect 18061 26333 18095 26367
rect 18613 26333 18647 26367
rect 18889 26333 18923 26367
rect 19257 26333 19291 26367
rect 20177 26333 20211 26367
rect 20453 26333 20487 26367
rect 21649 26333 21683 26367
rect 22385 26333 22419 26367
rect 23489 26333 23523 26367
rect 23765 26333 23799 26367
rect 24041 26333 24075 26367
rect 24869 26333 24903 26367
rect 25605 26333 25639 26367
rect 26249 26333 26283 26367
rect 26801 26333 26835 26367
rect 28089 26333 28123 26367
rect 28549 26333 28583 26367
rect 5641 26265 5675 26299
rect 11621 26265 11655 26299
rect 11713 26265 11747 26299
rect 12786 26265 12820 26299
rect 14289 26265 14323 26299
rect 18521 26265 18555 26299
rect 19901 26265 19935 26299
rect 27261 26265 27295 26299
rect 27997 26265 28031 26299
rect 4353 26197 4387 26231
rect 6377 26197 6411 26231
rect 6653 26197 6687 26231
rect 8309 26197 8343 26231
rect 8585 26197 8619 26231
rect 10425 26197 10459 26231
rect 11161 26197 11195 26231
rect 22293 26197 22327 26231
rect 23581 26197 23615 26231
rect 26065 26197 26099 26231
rect 26341 26197 26375 26231
rect 1777 25993 1811 26027
rect 5273 25993 5307 26027
rect 8033 25993 8067 26027
rect 10425 25993 10459 26027
rect 11345 25993 11379 26027
rect 22477 25993 22511 26027
rect 25053 25993 25087 26027
rect 26157 25993 26191 26027
rect 4997 25925 5031 25959
rect 6469 25925 6503 25959
rect 6561 25925 6595 25959
rect 1593 25857 1627 25891
rect 1961 25857 1995 25891
rect 2237 25857 2271 25891
rect 2605 25857 2639 25891
rect 2697 25857 2731 25891
rect 5189 25857 5223 25891
rect 5549 25857 5583 25891
rect 7941 25857 7975 25891
rect 8493 25857 8527 25891
rect 9965 25857 9999 25891
rect 11805 25857 11839 25891
rect 12357 25857 12391 25891
rect 14565 25857 14599 25891
rect 15209 25857 15243 25891
rect 15945 25857 15979 25891
rect 16865 25857 16899 25891
rect 17141 25857 17175 25891
rect 17233 25857 17267 25891
rect 17601 25857 17635 25891
rect 18521 25857 18555 25891
rect 19993 25857 20027 25891
rect 20269 25857 20303 25891
rect 21281 25857 21315 25891
rect 22753 25857 22787 25891
rect 22937 25857 22971 25891
rect 23857 25857 23891 25891
rect 24409 25857 24443 25891
rect 25237 25857 25271 25891
rect 26341 25857 26375 25891
rect 26985 25857 27019 25891
rect 27721 25857 27755 25891
rect 27905 25857 27939 25891
rect 2881 25789 2915 25823
rect 3433 25789 3467 25823
rect 3617 25789 3651 25823
rect 4353 25789 4387 25823
rect 4537 25789 4571 25823
rect 7205 25789 7239 25823
rect 8309 25789 8343 25823
rect 9045 25789 9079 25823
rect 9229 25789 9263 25823
rect 9781 25789 9815 25823
rect 10793 25789 10827 25823
rect 12449 25789 12483 25823
rect 12633 25789 12667 25823
rect 12909 25789 12943 25823
rect 15025 25789 15059 25823
rect 15761 25789 15795 25823
rect 17785 25789 17819 25823
rect 18705 25789 18739 25823
rect 20545 25789 20579 25823
rect 20729 25789 20763 25823
rect 21189 25789 21223 25823
rect 21833 25789 21867 25823
rect 22017 25789 22051 25823
rect 23121 25789 23155 25823
rect 23673 25789 23707 25823
rect 25513 25789 25547 25823
rect 25697 25789 25731 25823
rect 27169 25789 27203 25823
rect 2421 25721 2455 25755
rect 3341 25721 3375 25755
rect 3801 25721 3835 25755
rect 7021 25721 7055 25755
rect 8953 25721 8987 25755
rect 9413 25721 9447 25755
rect 19809 25721 19843 25755
rect 20085 25721 20119 25755
rect 26617 25721 26651 25755
rect 1409 25653 1443 25687
rect 2053 25653 2087 25687
rect 6101 25653 6135 25687
rect 7849 25653 7883 25687
rect 14381 25653 14415 25687
rect 15669 25653 15703 25687
rect 16129 25653 16163 25687
rect 16681 25653 16715 25687
rect 16957 25653 16991 25687
rect 17325 25653 17359 25687
rect 18245 25653 18279 25687
rect 18889 25653 18923 25687
rect 21373 25653 21407 25687
rect 22569 25653 22603 25687
rect 23581 25653 23615 25687
rect 24041 25653 24075 25687
rect 24593 25653 24627 25687
rect 27353 25653 27387 25687
rect 28089 25653 28123 25687
rect 3525 25449 3559 25483
rect 3985 25449 4019 25483
rect 4813 25449 4847 25483
rect 8401 25449 8435 25483
rect 9873 25449 9907 25483
rect 13921 25449 13955 25483
rect 17049 25449 17083 25483
rect 17601 25449 17635 25483
rect 18521 25449 18555 25483
rect 18705 25449 18739 25483
rect 21189 25449 21223 25483
rect 23121 25449 23155 25483
rect 27261 25449 27295 25483
rect 28089 25449 28123 25483
rect 28365 25449 28399 25483
rect 6469 25381 6503 25415
rect 8585 25381 8619 25415
rect 14841 25381 14875 25415
rect 18889 25381 18923 25415
rect 27997 25381 28031 25415
rect 5089 25313 5123 25347
rect 6837 25313 6871 25347
rect 12541 25313 12575 25347
rect 15393 25313 15427 25347
rect 15577 25313 15611 25347
rect 16129 25313 16163 25347
rect 16313 25313 16347 25347
rect 19257 25313 19291 25347
rect 19441 25313 19475 25347
rect 20913 25313 20947 25347
rect 21925 25313 21959 25347
rect 24501 25313 24535 25347
rect 25881 25313 25915 25347
rect 27353 25313 27387 25347
rect 1593 25245 1627 25279
rect 2053 25245 2087 25279
rect 2513 25245 2547 25279
rect 2605 25245 2639 25279
rect 2881 25245 2915 25279
rect 3157 25245 3191 25279
rect 3433 25245 3467 25279
rect 4169 25245 4203 25279
rect 4445 25245 4479 25279
rect 4721 25245 4755 25279
rect 4997 25245 5031 25279
rect 6745 25245 6779 25279
rect 7104 25245 7138 25279
rect 8309 25245 8343 25279
rect 8769 25245 8803 25279
rect 8953 25245 8987 25279
rect 9781 25245 9815 25279
rect 10241 25245 10275 25279
rect 10333 25245 10367 25279
rect 10600 25245 10634 25279
rect 11805 25245 11839 25279
rect 12797 25245 12831 25279
rect 14105 25245 14139 25279
rect 15025 25245 15059 25279
rect 15117 25245 15151 25279
rect 16957 25245 16991 25279
rect 17509 25241 17543 25275
rect 17785 25245 17819 25279
rect 17877 25245 17911 25279
rect 18613 25245 18647 25279
rect 19073 25245 19107 25279
rect 20729 25245 20763 25279
rect 22753 25245 22787 25279
rect 23029 25245 23063 25279
rect 23397 25245 23431 25279
rect 25789 25245 25823 25279
rect 26065 25245 26099 25279
rect 26617 25245 26651 25279
rect 26801 25245 26835 25279
rect 27537 25245 27571 25279
rect 28273 25245 28307 25279
rect 28549 25245 28583 25279
rect 2697 25177 2731 25211
rect 5356 25177 5390 25211
rect 24593 25177 24627 25211
rect 25513 25177 25547 25211
rect 1685 25109 1719 25143
rect 2145 25109 2179 25143
rect 2329 25109 2363 25143
rect 2973 25109 3007 25143
rect 3249 25109 3283 25143
rect 4261 25109 4295 25143
rect 4537 25109 4571 25143
rect 6561 25109 6595 25143
rect 8217 25109 8251 25143
rect 9597 25109 9631 25143
rect 10057 25109 10091 25143
rect 11713 25109 11747 25143
rect 12449 25109 12483 25143
rect 14749 25109 14783 25143
rect 15209 25109 15243 25143
rect 16037 25109 16071 25143
rect 16773 25109 16807 25143
rect 17325 25109 17359 25143
rect 19901 25109 19935 25143
rect 22477 25109 22511 25143
rect 22569 25109 22603 25143
rect 24041 25109 24075 25143
rect 25605 25109 25639 25143
rect 26525 25109 26559 25143
rect 14289 24905 14323 24939
rect 16129 24905 16163 24939
rect 18705 24905 18739 24939
rect 26341 24905 26375 24939
rect 26617 24905 26651 24939
rect 6653 24837 6687 24871
rect 23572 24837 23606 24871
rect 1593 24769 1627 24803
rect 2053 24769 2087 24803
rect 2513 24769 2547 24803
rect 2973 24769 3007 24803
rect 3065 24769 3099 24803
rect 3249 24769 3283 24803
rect 3801 24769 3835 24803
rect 4344 24769 4378 24803
rect 7389 24769 7423 24803
rect 7849 24769 7883 24803
rect 8309 24769 8343 24803
rect 9045 24769 9079 24803
rect 9312 24769 9346 24803
rect 10793 24769 10827 24803
rect 10885 24769 10919 24803
rect 11345 24769 11379 24803
rect 11621 24769 11655 24803
rect 12081 24769 12115 24803
rect 13176 24769 13210 24803
rect 15301 24769 15335 24803
rect 15853 24769 15887 24803
rect 16313 24769 16347 24803
rect 16865 24769 16899 24803
rect 17509 24769 17543 24803
rect 18429 24769 18463 24803
rect 18889 24769 18923 24803
rect 19717 24769 19751 24803
rect 20352 24769 20386 24803
rect 21833 24769 21867 24803
rect 22100 24769 22134 24803
rect 23305 24769 23339 24803
rect 25513 24769 25547 24803
rect 26249 24769 26283 24803
rect 26801 24769 26835 24803
rect 26985 24769 27019 24803
rect 27077 24769 27111 24803
rect 28089 24769 28123 24803
rect 28549 24769 28583 24803
rect 4077 24701 4111 24735
rect 5549 24701 5583 24735
rect 5733 24701 5767 24735
rect 6561 24701 6595 24735
rect 8585 24701 8619 24735
rect 10977 24701 11011 24735
rect 12173 24701 12207 24735
rect 12909 24701 12943 24735
rect 14381 24701 14415 24735
rect 14565 24701 14599 24735
rect 15117 24701 15151 24735
rect 17693 24701 17727 24735
rect 17877 24701 17911 24735
rect 18521 24701 18555 24735
rect 20085 24701 20119 24735
rect 24777 24701 24811 24735
rect 25697 24701 25731 24735
rect 27353 24701 27387 24735
rect 1869 24633 1903 24667
rect 2329 24633 2363 24667
rect 7113 24633 7147 24667
rect 11897 24633 11931 24667
rect 15945 24633 15979 24667
rect 17325 24633 17359 24667
rect 24685 24633 24719 24667
rect 26157 24633 26191 24667
rect 1685 24565 1719 24599
rect 2789 24565 2823 24599
rect 3709 24565 3743 24599
rect 3893 24565 3927 24599
rect 5457 24565 5491 24599
rect 6101 24565 6135 24599
rect 7481 24565 7515 24599
rect 7941 24565 7975 24599
rect 10425 24565 10459 24599
rect 10609 24565 10643 24599
rect 11161 24565 11195 24599
rect 11713 24565 11747 24599
rect 12817 24565 12851 24599
rect 15025 24565 15059 24599
rect 15485 24565 15519 24599
rect 16957 24565 16991 24599
rect 18245 24565 18279 24599
rect 19533 24565 19567 24599
rect 21465 24565 21499 24599
rect 23213 24565 23247 24599
rect 25421 24565 25455 24599
rect 27997 24565 28031 24599
rect 28181 24565 28215 24599
rect 28365 24565 28399 24599
rect 2789 24361 2823 24395
rect 4537 24361 4571 24395
rect 6101 24361 6135 24395
rect 6561 24361 6595 24395
rect 18245 24361 18279 24395
rect 23949 24361 23983 24395
rect 25513 24361 25547 24395
rect 27537 24361 27571 24395
rect 4169 24293 4203 24327
rect 8033 24293 8067 24327
rect 12541 24293 12575 24327
rect 14749 24293 14783 24327
rect 16129 24293 16163 24327
rect 16497 24293 16531 24327
rect 18521 24293 18555 24327
rect 19257 24293 19291 24327
rect 21925 24293 21959 24327
rect 25145 24293 25179 24327
rect 2881 24225 2915 24259
rect 3985 24225 4019 24259
rect 5549 24225 5583 24259
rect 6377 24225 6411 24259
rect 8677 24225 8711 24259
rect 9781 24225 9815 24259
rect 11161 24225 11195 24259
rect 12633 24225 12667 24259
rect 16957 24225 16991 24259
rect 17969 24225 18003 24259
rect 25973 24225 26007 24259
rect 1409 24157 1443 24191
rect 3801 24157 3835 24191
rect 4721 24157 4755 24191
rect 4813 24157 4847 24191
rect 5181 24157 5215 24191
rect 6193 24157 6227 24191
rect 7297 24157 7331 24191
rect 7665 24157 7699 24191
rect 7941 24157 7975 24191
rect 8217 24157 8251 24191
rect 8309 24157 8343 24191
rect 8585 24157 8619 24191
rect 9321 24157 9355 24191
rect 9597 24157 9631 24191
rect 10793 24157 10827 24191
rect 11069 24157 11103 24191
rect 13553 24133 13587 24167
rect 13921 24157 13955 24191
rect 14105 24157 14139 24191
rect 14381 24157 14415 24191
rect 14565 24157 14599 24191
rect 15197 24157 15231 24191
rect 15393 24157 15427 24191
rect 16313 24157 16347 24191
rect 16681 24157 16715 24191
rect 17141 24157 17175 24191
rect 17785 24157 17819 24191
rect 18705 24157 18739 24191
rect 19073 24157 19107 24191
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 19901 24157 19935 24191
rect 20821 24157 20855 24191
rect 21005 24157 21039 24191
rect 22109 24157 22143 24191
rect 22201 24157 22235 24191
rect 22477 24157 22511 24191
rect 23029 24157 23063 24191
rect 23121 24157 23155 24191
rect 23673 24157 23707 24191
rect 24133 24157 24167 24191
rect 24501 24157 24535 24191
rect 25329 24157 25363 24191
rect 25421 24157 25455 24191
rect 25881 24157 25915 24191
rect 27445 24157 27479 24191
rect 1676 24089 1710 24123
rect 5273 24089 5307 24123
rect 8401 24089 8435 24123
rect 10425 24089 10459 24123
rect 11428 24089 11462 24123
rect 20453 24089 20487 24123
rect 21649 24089 21683 24123
rect 26240 24089 26274 24123
rect 27905 24089 27939 24123
rect 27997 24089 28031 24123
rect 28549 24089 28583 24123
rect 3525 24021 3559 24055
rect 4905 24021 4939 24055
rect 7113 24021 7147 24055
rect 7481 24021 7515 24055
rect 7757 24021 7791 24055
rect 9137 24021 9171 24055
rect 10241 24021 10275 24055
rect 10885 24021 10919 24055
rect 13277 24021 13311 24055
rect 13369 24021 13403 24055
rect 13737 24021 13771 24055
rect 14197 24021 14231 24055
rect 15853 24021 15887 24055
rect 17601 24021 17635 24055
rect 18889 24021 18923 24055
rect 19625 24021 19659 24055
rect 21465 24021 21499 24055
rect 21741 24021 21775 24055
rect 22293 24021 22327 24055
rect 22569 24021 22603 24055
rect 22845 24021 22879 24055
rect 23213 24021 23247 24055
rect 23765 24021 23799 24055
rect 25053 24021 25087 24055
rect 25697 24021 25731 24055
rect 27353 24021 27387 24055
rect 2145 23817 2179 23851
rect 3617 23817 3651 23851
rect 6101 23817 6135 23851
rect 7021 23817 7055 23851
rect 9045 23817 9079 23851
rect 14013 23817 14047 23851
rect 14933 23817 14967 23851
rect 16129 23817 16163 23851
rect 26801 23817 26835 23851
rect 28365 23817 28399 23851
rect 9597 23749 9631 23783
rect 9689 23749 9723 23783
rect 10425 23749 10459 23783
rect 10517 23749 10551 23783
rect 11897 23749 11931 23783
rect 15853 23749 15887 23783
rect 19165 23749 19199 23783
rect 19993 23749 20027 23783
rect 25145 23749 25179 23783
rect 27252 23749 27286 23783
rect 2237 23681 2271 23715
rect 2504 23681 2538 23715
rect 3985 23681 4019 23715
rect 4629 23681 4663 23715
rect 5089 23681 5123 23715
rect 5641 23681 5675 23715
rect 6377 23681 6411 23715
rect 6561 23681 6595 23715
rect 7113 23681 7147 23715
rect 7573 23681 7607 23715
rect 9229 23681 9263 23715
rect 10241 23681 10275 23715
rect 11345 23681 11379 23715
rect 12889 23681 12923 23715
rect 14289 23681 14323 23715
rect 15301 23681 15335 23715
rect 16037 23681 16071 23715
rect 16957 23681 16991 23715
rect 17877 23681 17911 23715
rect 18613 23681 18647 23715
rect 19809 23681 19843 23715
rect 21833 23681 21867 23715
rect 22017 23681 22051 23715
rect 22845 23681 22879 23715
rect 23489 23681 23523 23715
rect 23756 23681 23790 23715
rect 26157 23681 26191 23715
rect 1593 23613 1627 23647
rect 5457 23613 5491 23647
rect 7389 23613 7423 23647
rect 8309 23613 8343 23647
rect 8493 23613 8527 23647
rect 11805 23613 11839 23647
rect 12633 23613 12667 23647
rect 14473 23613 14507 23647
rect 18061 23613 18095 23647
rect 19073 23613 19107 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 22661 23613 22695 23647
rect 25053 23613 25087 23647
rect 25329 23613 25363 23647
rect 26985 23613 27019 23647
rect 4721 23545 4755 23579
rect 10977 23545 11011 23579
rect 12357 23545 12391 23579
rect 18521 23545 18555 23579
rect 4537 23477 4571 23511
rect 5181 23477 5215 23511
rect 7205 23477 7239 23511
rect 7757 23477 7791 23511
rect 8677 23477 8711 23511
rect 11161 23477 11195 23511
rect 17049 23477 17083 23511
rect 18705 23477 18739 23511
rect 22201 23477 22235 23511
rect 23305 23477 23339 23511
rect 24869 23477 24903 23511
rect 2789 23273 2823 23307
rect 5181 23273 5215 23307
rect 5641 23273 5675 23307
rect 7205 23273 7239 23307
rect 7757 23273 7791 23307
rect 8677 23273 8711 23307
rect 8953 23273 8987 23307
rect 17601 23273 17635 23307
rect 18705 23273 18739 23307
rect 21373 23273 21407 23307
rect 22201 23273 22235 23307
rect 23213 23273 23247 23307
rect 23673 23273 23707 23307
rect 24409 23273 24443 23307
rect 26065 23273 26099 23307
rect 9229 23205 9263 23239
rect 17969 23205 18003 23239
rect 23949 23205 23983 23239
rect 26525 23205 26559 23239
rect 28457 23205 28491 23239
rect 3157 23137 3191 23171
rect 7389 23137 7423 23171
rect 7573 23137 7607 23171
rect 8309 23137 8343 23171
rect 10793 23137 10827 23171
rect 11989 23137 12023 23171
rect 12081 23137 12115 23171
rect 12817 23137 12851 23171
rect 15025 23137 15059 23171
rect 17417 23137 17451 23171
rect 19717 23137 19751 23171
rect 20729 23137 20763 23171
rect 20913 23137 20947 23171
rect 22661 23137 22695 23171
rect 22845 23137 22879 23171
rect 24685 23137 24719 23171
rect 1409 23069 1443 23103
rect 2973 23069 3007 23103
rect 3801 23069 3835 23103
rect 5825 23069 5859 23103
rect 8125 23069 8159 23103
rect 9137 23069 9171 23103
rect 9413 23069 9447 23103
rect 9505 23069 9539 23103
rect 9781 23069 9815 23103
rect 14105 23069 14139 23103
rect 14841 23069 14875 23103
rect 15761 23069 15795 23103
rect 17233 23069 17267 23103
rect 18153 23069 18187 23103
rect 18429 23069 18463 23103
rect 18889 23069 18923 23103
rect 20453 23069 20487 23103
rect 21557 23069 21591 23103
rect 21741 23069 21775 23103
rect 22293 23069 22327 23103
rect 23581 23069 23615 23103
rect 23857 23069 23891 23103
rect 24133 23069 24167 23103
rect 24593 23069 24627 23103
rect 24952 23069 24986 23103
rect 26249 23069 26283 23103
rect 26709 23069 26743 23103
rect 26985 23069 27019 23103
rect 27261 23069 27295 23103
rect 27721 23069 27755 23103
rect 1676 23001 1710 23035
rect 4068 23001 4102 23035
rect 5365 23001 5399 23035
rect 6092 23001 6126 23035
rect 10149 23001 10183 23035
rect 10241 23001 10275 23035
rect 10977 23001 11011 23035
rect 11069 23001 11103 23035
rect 12265 23001 12299 23035
rect 16028 23001 16062 23035
rect 19349 23001 19383 23035
rect 19441 23001 19475 23035
rect 27905 23001 27939 23035
rect 27997 23001 28031 23035
rect 3617 22933 3651 22967
rect 9597 22933 9631 22967
rect 9873 22933 9907 22967
rect 14749 22933 14783 22967
rect 15485 22933 15519 22967
rect 17141 22933 17175 22967
rect 18521 22933 18555 22967
rect 20545 22933 20579 22967
rect 22385 22933 22419 22967
rect 23397 22933 23431 22967
rect 26341 22933 26375 22967
rect 26801 22933 26835 22967
rect 27077 22933 27111 22967
rect 27537 22933 27571 22967
rect 2145 22729 2179 22763
rect 3341 22729 3375 22763
rect 4445 22729 4479 22763
rect 5181 22729 5215 22763
rect 7757 22729 7791 22763
rect 8493 22729 8527 22763
rect 14565 22729 14599 22763
rect 16221 22729 16255 22763
rect 17877 22729 17911 22763
rect 23765 22729 23799 22763
rect 24317 22729 24351 22763
rect 27813 22729 27847 22763
rect 28549 22729 28583 22763
rect 7021 22661 7055 22695
rect 8769 22661 8803 22695
rect 9597 22661 9631 22695
rect 10425 22661 10459 22695
rect 11713 22661 11747 22695
rect 13268 22661 13302 22695
rect 19073 22661 19107 22695
rect 19901 22661 19935 22695
rect 22753 22661 22787 22695
rect 1593 22593 1627 22627
rect 2053 22593 2087 22627
rect 2329 22593 2363 22627
rect 2421 22593 2455 22627
rect 3617 22593 3651 22627
rect 3801 22593 3835 22627
rect 4721 22593 4755 22627
rect 6193 22593 6227 22627
rect 6653 22593 6687 22627
rect 7297 22593 7331 22627
rect 8033 22593 8067 22627
rect 14473 22593 14507 22627
rect 15025 22593 15059 22627
rect 16037 22593 16071 22627
rect 16129 22593 16163 22627
rect 17141 22593 17175 22627
rect 17785 22593 17819 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 20913 22593 20947 22627
rect 21557 22593 21591 22627
rect 21833 22593 21867 22627
rect 22293 22593 22327 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 22937 22593 22971 22627
rect 23397 22593 23431 22627
rect 23673 22593 23707 22627
rect 23949 22593 23983 22627
rect 24041 22593 24075 22627
rect 24501 22593 24535 22627
rect 24777 22593 24811 22627
rect 25513 22593 25547 22627
rect 25973 22593 26007 22627
rect 26249 22593 26283 22627
rect 26341 22593 26375 22627
rect 26801 22593 26835 22627
rect 27353 22593 27387 22627
rect 28089 22593 28123 22627
rect 1685 22525 1719 22559
rect 2697 22525 2731 22559
rect 3985 22525 4019 22559
rect 4537 22525 4571 22559
rect 5273 22525 5307 22559
rect 7113 22525 7147 22559
rect 7849 22525 7883 22559
rect 8677 22525 8711 22559
rect 9505 22525 9539 22559
rect 9781 22525 9815 22559
rect 10333 22525 10367 22559
rect 10977 22525 11011 22559
rect 11621 22525 11655 22559
rect 11897 22525 11931 22559
rect 13001 22525 13035 22559
rect 15117 22525 15151 22559
rect 15301 22525 15335 22559
rect 15761 22525 15795 22559
rect 18153 22525 18187 22559
rect 18337 22525 18371 22559
rect 18981 22525 19015 22559
rect 19349 22525 19383 22559
rect 20821 22525 20855 22559
rect 25053 22525 25087 22559
rect 27169 22525 27203 22559
rect 27905 22525 27939 22559
rect 2513 22457 2547 22491
rect 9229 22457 9263 22491
rect 14381 22457 14415 22491
rect 14841 22457 14875 22491
rect 15853 22457 15887 22491
rect 20085 22457 20119 22491
rect 21925 22457 21959 22491
rect 22109 22457 22143 22491
rect 23213 22457 23247 22491
rect 1869 22389 1903 22423
rect 3433 22389 3467 22423
rect 5917 22389 5951 22423
rect 6009 22389 6043 22423
rect 17693 22389 17727 22423
rect 18797 22389 18831 22423
rect 22385 22389 22419 22423
rect 23029 22389 23063 22423
rect 23489 22389 23523 22423
rect 24133 22389 24167 22423
rect 25605 22389 25639 22423
rect 25789 22389 25823 22423
rect 26065 22389 26099 22423
rect 26433 22389 26467 22423
rect 26617 22389 26651 22423
rect 2789 22185 2823 22219
rect 3433 22185 3467 22219
rect 6377 22185 6411 22219
rect 7389 22185 7423 22219
rect 11713 22185 11747 22219
rect 14749 22185 14783 22219
rect 18981 22185 19015 22219
rect 19625 22185 19659 22219
rect 21281 22185 21315 22219
rect 23765 22185 23799 22219
rect 11529 22117 11563 22151
rect 13645 22117 13679 22151
rect 25053 22117 25087 22151
rect 25513 22117 25547 22151
rect 1409 22049 1443 22083
rect 3985 22049 4019 22083
rect 5273 22049 5307 22083
rect 8125 22049 8159 22083
rect 9321 22049 9355 22083
rect 10425 22049 10459 22083
rect 12265 22049 12299 22083
rect 14289 22049 14323 22083
rect 14933 22049 14967 22083
rect 19257 22049 19291 22083
rect 20085 22049 20119 22083
rect 21833 22049 21867 22083
rect 22569 22049 22603 22083
rect 23305 22049 23339 22083
rect 24593 22049 24627 22083
rect 25881 22049 25915 22083
rect 26065 22049 26099 22083
rect 27353 22049 27387 22083
rect 27537 22049 27571 22083
rect 3065 21981 3099 22015
rect 3157 21981 3191 22015
rect 3617 21981 3651 22015
rect 4169 21981 4203 22015
rect 4905 21981 4939 22015
rect 5181 21981 5215 22015
rect 5457 21981 5491 22015
rect 5917 21981 5951 22015
rect 6009 21981 6043 22015
rect 6193 21981 6227 22015
rect 6837 21981 6871 22015
rect 7665 21981 7699 22015
rect 8033 21981 8067 22015
rect 8493 21981 8527 22015
rect 8769 21981 8803 22015
rect 9137 21981 9171 22015
rect 11897 21981 11931 22015
rect 12173 21981 12207 22015
rect 13737 21981 13771 22015
rect 13829 21981 13863 22015
rect 14105 21981 14139 22015
rect 14841 21981 14875 22015
rect 15393 21981 15427 22015
rect 16497 21981 16531 22015
rect 16589 21981 16623 22015
rect 16856 21981 16890 22015
rect 18153 21981 18187 22015
rect 18889 21981 18923 22015
rect 19441 21981 19475 22015
rect 19993 21981 20027 22015
rect 20821 21981 20855 22015
rect 20913 21981 20947 22015
rect 21097 21981 21131 22015
rect 21649 21981 21683 22015
rect 22385 21981 22419 22015
rect 23121 21981 23155 22015
rect 23857 21981 23891 22015
rect 24409 21981 24443 22015
rect 25145 21981 25179 22015
rect 25329 21981 25363 22015
rect 26617 21981 26651 22015
rect 26801 21981 26835 22015
rect 28273 21981 28307 22015
rect 1676 21913 1710 21947
rect 3249 21913 3283 21947
rect 9413 21913 9447 21947
rect 9965 21913 9999 21947
rect 10149 21913 10183 21947
rect 10241 21913 10275 21947
rect 10977 21913 11011 21947
rect 11069 21913 11103 21947
rect 12532 21913 12566 21947
rect 15761 21913 15795 21947
rect 20361 21913 20395 21947
rect 27261 21913 27295 21947
rect 27997 21913 28031 21947
rect 2881 21845 2915 21879
rect 4629 21845 4663 21879
rect 4721 21845 4755 21879
rect 4997 21845 5031 21879
rect 7757 21845 7791 21879
rect 8309 21845 8343 21879
rect 8585 21845 8619 21879
rect 8953 21845 8987 21879
rect 11989 21845 12023 21879
rect 16313 21845 16347 21879
rect 17969 21845 18003 21879
rect 18705 21845 18739 21879
rect 20453 21845 20487 21879
rect 20637 21845 20671 21879
rect 22293 21845 22327 21879
rect 23029 21845 23063 21879
rect 23949 21845 23983 21879
rect 26525 21845 26559 21879
rect 28089 21845 28123 21879
rect 28365 21845 28399 21879
rect 2237 21641 2271 21675
rect 4813 21641 4847 21675
rect 6193 21641 6227 21675
rect 6377 21641 6411 21675
rect 13829 21641 13863 21675
rect 15393 21641 15427 21675
rect 17325 21641 17359 21675
rect 23305 21641 23339 21675
rect 24133 21641 24167 21675
rect 24961 21641 24995 21675
rect 25329 21641 25363 21675
rect 26249 21641 26283 21675
rect 26709 21641 26743 21675
rect 7113 21573 7147 21607
rect 10793 21573 10827 21607
rect 12532 21573 12566 21607
rect 27414 21573 27448 21607
rect 1685 21505 1719 21539
rect 2329 21505 2363 21539
rect 2789 21505 2823 21539
rect 3525 21505 3559 21539
rect 4169 21505 4203 21539
rect 5089 21505 5123 21539
rect 5457 21505 5491 21539
rect 5733 21505 5767 21539
rect 6561 21505 6595 21539
rect 6745 21505 6779 21539
rect 7849 21505 7883 21539
rect 8125 21505 8159 21539
rect 8677 21505 8711 21539
rect 9873 21505 9907 21539
rect 10517 21505 10551 21539
rect 11621 21505 11655 21539
rect 13737 21505 13771 21539
rect 14841 21505 14875 21539
rect 15117 21505 15151 21539
rect 15209 21505 15243 21539
rect 15577 21505 15611 21539
rect 17509 21505 17543 21539
rect 17877 21505 17911 21539
rect 18144 21505 18178 21539
rect 19533 21505 19567 21539
rect 20269 21505 20303 21539
rect 20453 21505 20487 21539
rect 21189 21505 21223 21539
rect 22017 21505 22051 21539
rect 22109 21505 22143 21539
rect 22845 21505 22879 21539
rect 25237 21505 25271 21539
rect 25513 21505 25547 21539
rect 26525 21505 26559 21539
rect 26617 21505 26651 21539
rect 27169 21505 27203 21539
rect 2605 21437 2639 21471
rect 3341 21437 3375 21471
rect 4353 21437 4387 21471
rect 5549 21437 5583 21471
rect 8217 21437 8251 21471
rect 9045 21437 9079 21471
rect 10701 21437 10735 21471
rect 12265 21437 12299 21471
rect 15761 21437 15795 21471
rect 21005 21437 21039 21471
rect 22385 21437 22419 21471
rect 22661 21437 22695 21471
rect 23489 21437 23523 21471
rect 23673 21437 23707 21471
rect 24317 21437 24351 21471
rect 24501 21437 24535 21471
rect 25605 21437 25639 21471
rect 25789 21437 25823 21471
rect 2421 21369 2455 21403
rect 7665 21369 7699 21403
rect 9597 21369 9631 21403
rect 11253 21369 11287 21403
rect 14657 21369 14691 21403
rect 19257 21369 19291 21403
rect 21833 21369 21867 21403
rect 25053 21369 25087 21403
rect 26341 21369 26375 21403
rect 3249 21301 3283 21335
rect 3709 21301 3743 21335
rect 7941 21301 7975 21335
rect 8493 21301 8527 21335
rect 12173 21301 12207 21335
rect 13645 21301 13679 21335
rect 14933 21301 14967 21335
rect 16129 21301 16163 21335
rect 20085 21301 20119 21335
rect 20913 21301 20947 21335
rect 21373 21301 21407 21335
rect 22293 21301 22327 21335
rect 28549 21301 28583 21335
rect 2789 21097 2823 21131
rect 3525 21097 3559 21131
rect 4537 21097 4571 21131
rect 4813 21097 4847 21131
rect 6469 21097 6503 21131
rect 8769 21097 8803 21131
rect 13277 21097 13311 21131
rect 15301 21097 15335 21131
rect 16129 21097 16163 21131
rect 21741 21097 21775 21131
rect 22293 21097 22327 21131
rect 24133 21097 24167 21131
rect 24961 21097 24995 21131
rect 12541 21029 12575 21063
rect 18337 21029 18371 21063
rect 18705 21029 18739 21063
rect 20729 21029 20763 21063
rect 26985 21029 27019 21063
rect 1409 20961 1443 20995
rect 3249 20961 3283 20995
rect 3985 20961 4019 20995
rect 6653 20961 6687 20995
rect 10885 20961 10919 20995
rect 12725 20961 12759 20995
rect 15669 20961 15703 20995
rect 16313 20961 16347 20995
rect 21097 20961 21131 20995
rect 22017 20961 22051 20995
rect 22753 20961 22787 20995
rect 23213 20961 23247 20995
rect 23489 20961 23523 20995
rect 26801 20961 26835 20995
rect 27997 20961 28031 20995
rect 3065 20893 3099 20927
rect 3157 20893 3191 20927
rect 3433 20893 3467 20927
rect 3801 20893 3835 20927
rect 4721 20893 4755 20927
rect 4997 20893 5031 20927
rect 5089 20893 5123 20927
rect 5356 20893 5390 20927
rect 7389 20893 7423 20927
rect 11161 20893 11195 20927
rect 13829 20893 13863 20927
rect 15209 20893 15243 20927
rect 15485 20893 15519 20927
rect 16497 20893 16531 20927
rect 16957 20893 16991 20927
rect 17325 20893 17359 20927
rect 17509 20893 17543 20927
rect 18153 20893 18187 20927
rect 18429 20893 18463 20927
rect 18889 20893 18923 20927
rect 19257 20893 19291 20927
rect 20913 20893 20947 20927
rect 21281 20893 21315 20927
rect 21833 20893 21867 20927
rect 22569 20893 22603 20927
rect 23305 20893 23339 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24593 20893 24627 20927
rect 24869 20893 24903 20927
rect 25145 20893 25179 20927
rect 26617 20893 26651 20927
rect 27353 20893 27387 20927
rect 27813 20893 27847 20927
rect 27905 20893 27939 20927
rect 28549 20893 28583 20927
rect 1676 20825 1710 20859
rect 7656 20825 7690 20859
rect 9045 20825 9079 20859
rect 9137 20825 9171 20859
rect 10057 20825 10091 20859
rect 10149 20825 10183 20859
rect 11406 20825 11440 20859
rect 18521 20825 18555 20859
rect 19524 20825 19558 20859
rect 2881 20757 2915 20791
rect 4445 20757 4479 20791
rect 7297 20757 7331 20791
rect 13369 20757 13403 20791
rect 13645 20757 13679 20791
rect 17049 20757 17083 20791
rect 17969 20757 18003 20791
rect 20637 20757 20671 20791
rect 24409 20757 24443 20791
rect 24685 20757 24719 20791
rect 27445 20757 27479 20791
rect 27629 20757 27663 20791
rect 28365 20757 28399 20791
rect 2605 20553 2639 20587
rect 3525 20553 3559 20587
rect 8217 20553 8251 20587
rect 8769 20553 8803 20587
rect 13185 20553 13219 20587
rect 16037 20553 16071 20587
rect 17325 20553 17359 20587
rect 17417 20553 17451 20587
rect 24041 20553 24075 20587
rect 24317 20553 24351 20587
rect 26617 20553 26651 20587
rect 27629 20553 27663 20587
rect 28365 20553 28399 20587
rect 7104 20485 7138 20519
rect 18245 20485 18279 20519
rect 20729 20485 20763 20519
rect 21925 20485 21959 20519
rect 22017 20485 22051 20519
rect 23857 20485 23891 20519
rect 1409 20417 1443 20451
rect 1685 20417 1719 20451
rect 3709 20417 3743 20451
rect 3985 20417 4019 20451
rect 4077 20417 4111 20451
rect 4537 20417 4571 20451
rect 4629 20417 4663 20451
rect 4905 20417 4939 20451
rect 5825 20417 5859 20451
rect 6009 20417 6043 20451
rect 6561 20417 6595 20451
rect 6837 20417 6871 20451
rect 8677 20417 8711 20451
rect 8953 20417 8987 20451
rect 9045 20417 9079 20451
rect 9588 20417 9622 20451
rect 10793 20417 10827 20451
rect 11161 20417 11195 20451
rect 11529 20417 11563 20451
rect 11796 20417 11830 20451
rect 13369 20417 13403 20451
rect 13645 20417 13679 20451
rect 13921 20417 13955 20451
rect 14197 20417 14231 20451
rect 14933 20417 14967 20451
rect 15945 20417 15979 20451
rect 16405 20417 16439 20451
rect 16681 20417 16715 20451
rect 17601 20417 17635 20451
rect 18061 20417 18095 20451
rect 19993 20417 20027 20451
rect 23029 20417 23063 20451
rect 24225 20417 24259 20451
rect 24501 20417 24535 20451
rect 24777 20417 24811 20451
rect 25053 20417 25087 20451
rect 26525 20417 26559 20451
rect 26801 20417 26835 20451
rect 27169 20417 27203 20451
rect 27905 20417 27939 20451
rect 2053 20349 2087 20383
rect 2789 20349 2823 20383
rect 5089 20349 5123 20383
rect 9321 20349 9355 20383
rect 11253 20349 11287 20383
rect 14381 20349 14415 20383
rect 15025 20349 15059 20383
rect 15209 20349 15243 20383
rect 15393 20349 15427 20383
rect 16865 20349 16899 20383
rect 18981 20349 19015 20383
rect 21005 20349 21039 20383
rect 22201 20349 22235 20383
rect 24869 20349 24903 20383
rect 25605 20349 25639 20383
rect 25789 20349 25823 20383
rect 26985 20349 27019 20383
rect 27721 20349 27755 20383
rect 1777 20281 1811 20315
rect 4721 20281 4755 20315
rect 8493 20281 8527 20315
rect 12909 20281 12943 20315
rect 14841 20281 14875 20315
rect 24593 20281 24627 20315
rect 1501 20213 1535 20247
rect 3341 20213 3375 20247
rect 3801 20213 3835 20247
rect 4169 20213 4203 20247
rect 4353 20213 4387 20247
rect 5273 20213 5307 20247
rect 5641 20213 5675 20247
rect 6101 20213 6135 20247
rect 6653 20213 6687 20247
rect 9229 20213 9263 20247
rect 10701 20213 10735 20247
rect 10977 20213 11011 20247
rect 13461 20213 13495 20247
rect 13737 20213 13771 20247
rect 15853 20213 15887 20247
rect 16221 20213 16255 20247
rect 21649 20213 21683 20247
rect 25513 20213 25547 20247
rect 25973 20213 26007 20247
rect 26341 20213 26375 20247
rect 2789 20009 2823 20043
rect 4261 20009 4295 20043
rect 4537 20009 4571 20043
rect 7849 20009 7883 20043
rect 14841 20009 14875 20043
rect 16037 20009 16071 20043
rect 16497 20009 16531 20043
rect 17969 20009 18003 20043
rect 20637 20009 20671 20043
rect 25605 20009 25639 20043
rect 26709 20009 26743 20043
rect 27261 20009 27295 20043
rect 9781 19941 9815 19975
rect 10241 19941 10275 19975
rect 13737 19941 13771 19975
rect 15853 19941 15887 19975
rect 18797 19941 18831 19975
rect 24133 19941 24167 19975
rect 26617 19941 26651 19975
rect 6377 19873 6411 19907
rect 7389 19873 7423 19907
rect 12725 19873 12759 19907
rect 13185 19873 13219 19907
rect 14197 19873 14231 19907
rect 14381 19873 14415 19907
rect 17141 19873 17175 19907
rect 17509 19873 17543 19907
rect 20821 19873 20855 19907
rect 25973 19873 26007 19907
rect 26157 19873 26191 19907
rect 1409 19805 1443 19839
rect 2973 19805 3007 19839
rect 3157 19805 3191 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 4721 19805 4755 19839
rect 5641 19805 5675 19839
rect 6653 19805 6687 19839
rect 8033 19805 8067 19839
rect 8125 19805 8159 19839
rect 8309 19805 8343 19839
rect 9137 19805 9171 19839
rect 9321 19805 9355 19839
rect 9873 19805 9907 19839
rect 10057 19805 10091 19839
rect 13001 19805 13035 19839
rect 13921 19805 13955 19839
rect 15209 19805 15243 19839
rect 15393 19805 15427 19839
rect 15945 19805 15979 19839
rect 16681 19805 16715 19839
rect 17049 19805 17083 19839
rect 17325 19805 17359 19839
rect 18153 19805 18187 19839
rect 18981 19805 19015 19839
rect 19257 19805 19291 19839
rect 22017 19805 22051 19839
rect 22753 19805 22787 19839
rect 24593 19805 24627 19839
rect 24685 19805 24719 19839
rect 25145 19805 25179 19839
rect 25421 19805 25455 19839
rect 25513 19805 25547 19839
rect 26893 19805 26927 19839
rect 26985 19805 27019 19839
rect 27445 19805 27479 19839
rect 27537 19805 27571 19839
rect 27905 19805 27939 19839
rect 28181 19805 28215 19839
rect 1676 19737 1710 19771
rect 4905 19737 4939 19771
rect 4997 19737 5031 19771
rect 5549 19737 5583 19771
rect 10885 19737 10919 19771
rect 10977 19737 11011 19771
rect 11897 19737 11931 19771
rect 11989 19737 12023 19771
rect 19524 19737 19558 19771
rect 20913 19737 20947 19771
rect 21833 19737 21867 19771
rect 22569 19737 22603 19771
rect 23020 19737 23054 19771
rect 28273 19737 28307 19771
rect 3617 19669 3651 19703
rect 8769 19669 8803 19703
rect 13645 19669 13679 19703
rect 18705 19669 18739 19703
rect 24409 19669 24443 19703
rect 24777 19669 24811 19703
rect 24961 19669 24995 19703
rect 25237 19669 25271 19703
rect 27077 19669 27111 19703
rect 27721 19669 27755 19703
rect 27997 19669 28031 19703
rect 2789 19465 2823 19499
rect 3525 19465 3559 19499
rect 3893 19465 3927 19499
rect 5365 19465 5399 19499
rect 5733 19465 5767 19499
rect 13001 19465 13035 19499
rect 14933 19465 14967 19499
rect 15761 19465 15795 19499
rect 16037 19465 16071 19499
rect 18061 19465 18095 19499
rect 21465 19465 21499 19499
rect 22477 19465 22511 19499
rect 22569 19465 22603 19499
rect 6561 19397 6595 19431
rect 7849 19397 7883 19431
rect 9689 19397 9723 19431
rect 10425 19397 10459 19431
rect 11345 19397 11379 19431
rect 12265 19397 12299 19431
rect 13369 19397 13403 19431
rect 20821 19397 20855 19431
rect 23213 19397 23247 19431
rect 1409 19329 1443 19363
rect 1676 19329 1710 19363
rect 2881 19329 2915 19363
rect 3801 19329 3835 19363
rect 4077 19329 4111 19363
rect 4721 19329 4755 19363
rect 4905 19329 4939 19363
rect 5641 19329 5675 19363
rect 5917 19329 5951 19363
rect 6009 19329 6043 19363
rect 7573 19329 7607 19363
rect 7665 19329 7699 19363
rect 9505 19329 9539 19363
rect 9597 19329 9631 19363
rect 10057 19329 10091 19363
rect 11621 19329 11655 19363
rect 12357 19329 12391 19363
rect 13277 19329 13311 19363
rect 14197 19329 14231 19363
rect 15669 19329 15703 19363
rect 15945 19329 15979 19363
rect 16221 19329 16255 19363
rect 16948 19329 16982 19363
rect 18153 19329 18187 19363
rect 20085 19329 20119 19363
rect 21097 19329 21131 19363
rect 21365 19335 21399 19369
rect 22753 19329 22787 19363
rect 23029 19329 23063 19363
rect 24041 19329 24075 19363
rect 24225 19329 24259 19363
rect 25881 19329 25915 19363
rect 26433 19329 26467 19363
rect 26985 19329 27019 19363
rect 27169 19329 27203 19363
rect 27629 19329 27663 19363
rect 28365 19329 28399 19363
rect 3065 19261 3099 19295
rect 6469 19261 6503 19295
rect 10333 19261 10367 19295
rect 11805 19261 11839 19295
rect 12541 19261 12575 19295
rect 13645 19261 13679 19295
rect 14289 19261 14323 19295
rect 14473 19261 14507 19295
rect 15025 19261 15059 19295
rect 15209 19261 15243 19295
rect 16681 19261 16715 19295
rect 18337 19261 18371 19295
rect 18981 19261 19015 19295
rect 21833 19261 21867 19295
rect 24409 19261 24443 19295
rect 24961 19261 24995 19295
rect 25697 19261 25731 19295
rect 27721 19261 27755 19295
rect 27905 19261 27939 19295
rect 7021 19193 7055 19227
rect 22845 19193 22879 19227
rect 3617 19125 3651 19159
rect 5457 19125 5491 19159
rect 6101 19125 6135 19159
rect 7389 19125 7423 19159
rect 9873 19125 9907 19159
rect 21189 19125 21223 19159
rect 24869 19125 24903 19159
rect 25605 19125 25639 19159
rect 26341 19125 26375 19159
rect 26525 19125 26559 19159
rect 2237 18921 2271 18955
rect 5457 18921 5491 18955
rect 6193 18921 6227 18955
rect 9045 18921 9079 18955
rect 10241 18921 10275 18955
rect 10977 18921 11011 18955
rect 12449 18921 12483 18955
rect 13093 18921 13127 18955
rect 14105 18921 14139 18955
rect 18889 18921 18923 18955
rect 23489 18921 23523 18955
rect 25513 18921 25547 18955
rect 26341 18921 26375 18955
rect 4537 18853 4571 18887
rect 24225 18853 24259 18887
rect 25053 18853 25087 18887
rect 28365 18853 28399 18887
rect 1685 18785 1719 18819
rect 4997 18785 5031 18819
rect 5549 18785 5583 18819
rect 6653 18785 6687 18819
rect 7113 18785 7147 18819
rect 7573 18785 7607 18819
rect 9781 18785 9815 18819
rect 12817 18785 12851 18819
rect 13461 18785 13495 18819
rect 19625 18785 19659 18819
rect 20913 18785 20947 18819
rect 23581 18785 23615 18819
rect 25145 18785 25179 18819
rect 25881 18785 25915 18819
rect 26065 18785 26099 18819
rect 26617 18785 26651 18819
rect 26801 18785 26835 18819
rect 27445 18785 27479 18819
rect 27629 18785 27663 18819
rect 2421 18717 2455 18751
rect 2697 18717 2731 18751
rect 3433 18717 3467 18751
rect 3525 18717 3559 18751
rect 3801 18717 3835 18751
rect 3985 18717 4019 18751
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 5733 18717 5767 18751
rect 6469 18717 6503 18751
rect 8585 18717 8619 18751
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 9597 18717 9631 18751
rect 10333 18717 10367 18751
rect 11161 18717 11195 18751
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 12633 18717 12667 18751
rect 13369 18717 13403 18751
rect 13829 18717 13863 18751
rect 14289 18717 14323 18751
rect 15393 18717 15427 18751
rect 15577 18717 15611 18751
rect 17417 18717 17451 18751
rect 17509 18717 17543 18751
rect 17776 18717 17810 18751
rect 19441 18717 19475 18751
rect 21373 18717 21407 18751
rect 22845 18717 22879 18751
rect 23765 18717 23799 18751
rect 24409 18717 24443 18751
rect 24593 18717 24627 18751
rect 25329 18717 25363 18751
rect 28549 18717 28583 18751
rect 3341 18649 3375 18683
rect 7297 18649 7331 18683
rect 7389 18649 7423 18683
rect 11713 18649 11747 18683
rect 21640 18649 21674 18683
rect 2513 18581 2547 18615
rect 4445 18581 4479 18615
rect 8401 18581 8435 18615
rect 9413 18581 9447 18615
rect 13645 18581 13679 18615
rect 16037 18581 16071 18615
rect 17233 18581 17267 18615
rect 22753 18581 22787 18615
rect 27261 18581 27295 18615
rect 28089 18581 28123 18615
rect 2789 18377 2823 18411
rect 3801 18377 3835 18411
rect 5089 18377 5123 18411
rect 8401 18377 8435 18411
rect 9597 18377 9631 18411
rect 10609 18377 10643 18411
rect 11621 18377 11655 18411
rect 12541 18377 12575 18411
rect 13185 18377 13219 18411
rect 14933 18377 14967 18411
rect 16129 18377 16163 18411
rect 17325 18377 17359 18411
rect 21005 18377 21039 18411
rect 21373 18377 21407 18411
rect 22477 18377 22511 18411
rect 23949 18377 23983 18411
rect 24225 18377 24259 18411
rect 24869 18377 24903 18411
rect 25145 18377 25179 18411
rect 28365 18377 28399 18411
rect 1676 18309 1710 18343
rect 3617 18309 3651 18343
rect 4629 18309 4663 18343
rect 21189 18309 21223 18343
rect 25688 18309 25722 18343
rect 1409 18241 1443 18275
rect 2973 18241 3007 18275
rect 3709 18241 3743 18275
rect 3985 18241 4019 18275
rect 4721 18241 4755 18275
rect 4997 18241 5031 18275
rect 5457 18241 5491 18275
rect 6009 18241 6043 18275
rect 6745 18241 6779 18275
rect 8217 18241 8251 18275
rect 9505 18241 9539 18275
rect 9965 18241 9999 18275
rect 10701 18241 10735 18275
rect 11345 18241 11379 18275
rect 11805 18241 11839 18275
rect 12081 18241 12115 18275
rect 13093 18241 13127 18275
rect 14841 18241 14875 18275
rect 15117 18241 15151 18275
rect 15209 18241 15243 18275
rect 15301 18241 15335 18275
rect 15669 18241 15703 18275
rect 16221 18241 16255 18275
rect 16681 18241 16715 18275
rect 17601 18241 17635 18275
rect 17693 18241 17727 18275
rect 18337 18241 18371 18275
rect 19809 18241 19843 18275
rect 20545 18241 20579 18275
rect 21097 18241 21131 18275
rect 21557 18241 21591 18275
rect 21833 18241 21867 18275
rect 22937 18241 22971 18275
rect 24133 18241 24167 18275
rect 24409 18241 24443 18275
rect 24685 18241 24719 18275
rect 24777 18241 24811 18275
rect 25053 18241 25087 18275
rect 27077 18241 27111 18275
rect 27721 18241 27755 18275
rect 3157 18173 3191 18207
rect 4169 18173 4203 18207
rect 4813 18173 4847 18207
rect 5549 18173 5583 18207
rect 6377 18173 6411 18207
rect 8769 18173 8803 18207
rect 8953 18173 8987 18207
rect 9413 18173 9447 18207
rect 10149 18173 10183 18207
rect 10793 18173 10827 18207
rect 11897 18173 11931 18207
rect 15485 18173 15519 18207
rect 17969 18173 18003 18207
rect 20361 18173 20395 18207
rect 23213 18173 23247 18207
rect 23397 18173 23431 18207
rect 25421 18173 25455 18207
rect 27905 18173 27939 18207
rect 6101 18105 6135 18139
rect 11161 18105 11195 18139
rect 14657 18105 14691 18139
rect 17417 18105 17451 18139
rect 19993 18105 20027 18139
rect 26801 18105 26835 18139
rect 16313 18037 16347 18071
rect 17785 18037 17819 18071
rect 22753 18037 22787 18071
rect 23857 18037 23891 18071
rect 24501 18037 24535 18071
rect 27629 18037 27663 18071
rect 2789 17833 2823 17867
rect 2973 17833 3007 17867
rect 4813 17833 4847 17867
rect 6561 17833 6595 17867
rect 6837 17833 6871 17867
rect 7021 17833 7055 17867
rect 7389 17833 7423 17867
rect 9321 17833 9355 17867
rect 19349 17833 19383 17867
rect 21097 17833 21131 17867
rect 24041 17833 24075 17867
rect 25881 17833 25915 17867
rect 4905 17765 4939 17799
rect 8769 17765 8803 17799
rect 9965 17765 9999 17799
rect 14749 17765 14783 17799
rect 15209 17765 15243 17799
rect 16589 17765 16623 17799
rect 17049 17765 17083 17799
rect 18061 17765 18095 17799
rect 21649 17765 21683 17799
rect 21925 17765 21959 17799
rect 22845 17765 22879 17799
rect 23305 17765 23339 17799
rect 25789 17765 25823 17799
rect 1409 17697 1443 17731
rect 4353 17697 4387 17731
rect 8309 17697 8343 17731
rect 9137 17697 9171 17731
rect 10333 17697 10367 17731
rect 13829 17697 13863 17731
rect 15025 17697 15059 17731
rect 15945 17697 15979 17731
rect 16865 17697 16899 17731
rect 18337 17697 18371 17731
rect 18613 17697 18647 17731
rect 22385 17697 22419 17731
rect 24409 17697 24443 17731
rect 24593 17697 24627 17731
rect 26249 17697 26283 17731
rect 26893 17697 26927 17731
rect 3157 17629 3191 17663
rect 4077 17629 4111 17663
rect 4169 17629 4203 17663
rect 5089 17629 5123 17663
rect 6469 17629 6503 17663
rect 6653 17629 6687 17663
rect 6745 17629 6779 17663
rect 7205 17629 7239 17663
rect 7297 17629 7331 17663
rect 7757 17629 7791 17663
rect 8033 17629 8067 17663
rect 8125 17629 8159 17663
rect 8953 17629 8987 17663
rect 9873 17629 9907 17663
rect 10149 17629 10183 17663
rect 12449 17629 12483 17663
rect 13645 17605 13679 17639
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 14841 17629 14875 17663
rect 15853 17629 15887 17663
rect 16129 17629 16163 17663
rect 16681 17629 16715 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 19717 17629 19751 17663
rect 19984 17629 20018 17663
rect 21833 17629 21867 17663
rect 22109 17629 22143 17663
rect 22201 17629 22235 17663
rect 22937 17629 22971 17663
rect 23121 17629 23155 17663
rect 23857 17629 23891 17663
rect 23949 17629 23983 17663
rect 25145 17629 25179 17663
rect 25329 17629 25363 17663
rect 26065 17629 26099 17663
rect 26157 17629 26191 17663
rect 26433 17629 26467 17663
rect 28549 17629 28583 17663
rect 1676 17561 1710 17595
rect 10600 17561 10634 17595
rect 17509 17561 17543 17595
rect 17601 17561 17635 17595
rect 18429 17561 18463 17595
rect 26617 17561 26651 17595
rect 3893 17493 3927 17527
rect 7573 17493 7607 17527
rect 7849 17493 7883 17527
rect 9689 17493 9723 17527
rect 11713 17493 11747 17527
rect 12265 17493 12299 17527
rect 13461 17493 13495 17527
rect 15669 17493 15703 17527
rect 23673 17493 23707 17527
rect 25053 17493 25087 17527
rect 28365 17493 28399 17527
rect 2329 17289 2363 17323
rect 4721 17289 4755 17323
rect 6009 17289 6043 17323
rect 10149 17289 10183 17323
rect 12541 17289 12575 17323
rect 13277 17289 13311 17323
rect 14013 17289 14047 17323
rect 16681 17289 16715 17323
rect 16957 17289 16991 17323
rect 17877 17289 17911 17323
rect 20085 17289 20119 17323
rect 22661 17289 22695 17323
rect 23857 17289 23891 17323
rect 27629 17289 27663 17323
rect 25320 17221 25354 17255
rect 2513 17153 2547 17187
rect 2973 17153 3007 17187
rect 3065 17153 3099 17187
rect 3433 17153 3467 17187
rect 3985 17153 4019 17187
rect 4905 17153 4939 17187
rect 5365 17153 5399 17187
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 7941 17153 7975 17187
rect 8217 17153 8251 17187
rect 10241 17153 10275 17187
rect 11621 17153 11655 17187
rect 11713 17153 11747 17187
rect 12081 17153 12115 17187
rect 13553 17153 13587 17187
rect 14197 17153 14231 17187
rect 15025 17153 15059 17187
rect 16313 17153 16347 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 17233 17153 17267 17187
rect 17693 17153 17727 17187
rect 17785 17153 17819 17187
rect 19165 17153 19199 17187
rect 19901 17153 19935 17187
rect 20269 17153 20303 17187
rect 20453 17153 20487 17187
rect 21649 17153 21683 17187
rect 22569 17153 22603 17187
rect 23397 17153 23431 17187
rect 25053 17153 25087 17187
rect 26709 17153 26743 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 27905 17153 27939 17187
rect 1777 17085 1811 17119
rect 3249 17085 3283 17119
rect 4169 17085 4203 17119
rect 6561 17085 6595 17119
rect 8033 17085 8067 17119
rect 8769 17085 8803 17119
rect 8953 17085 8987 17119
rect 9505 17085 9539 17119
rect 9689 17085 9723 17119
rect 10333 17085 10367 17119
rect 10701 17085 10735 17119
rect 10885 17085 10919 17119
rect 11345 17085 11379 17119
rect 11897 17085 11931 17119
rect 12633 17085 12667 17119
rect 12817 17085 12851 17119
rect 15577 17085 15611 17119
rect 15761 17085 15795 17119
rect 20637 17085 20671 17119
rect 20729 17085 20763 17119
rect 20913 17085 20947 17119
rect 23213 17085 23247 17119
rect 24225 17085 24259 17119
rect 27721 17085 27755 17119
rect 3893 17017 3927 17051
rect 4353 17017 4387 17051
rect 5181 17017 5215 17051
rect 7757 17017 7791 17051
rect 8677 17017 8711 17051
rect 9137 17017 9171 17051
rect 13369 17017 13403 17051
rect 21465 17017 21499 17051
rect 28181 17017 28215 17051
rect 2789 16949 2823 16983
rect 6929 16949 6963 16983
rect 7113 16949 7147 16983
rect 7573 16949 7607 16983
rect 14841 16949 14875 16983
rect 16221 16949 16255 16983
rect 16405 16949 16439 16983
rect 17325 16949 17359 16983
rect 17509 16949 17543 16983
rect 19349 16949 19383 16983
rect 19717 16949 19751 16983
rect 21097 16949 21131 16983
rect 24777 16949 24811 16983
rect 26433 16949 26467 16983
rect 26525 16949 26559 16983
rect 3065 16745 3099 16779
rect 3249 16745 3283 16779
rect 4629 16745 4663 16779
rect 9045 16745 9079 16779
rect 10057 16745 10091 16779
rect 10977 16745 11011 16779
rect 11805 16745 11839 16779
rect 12725 16745 12759 16779
rect 15485 16745 15519 16779
rect 16221 16745 16255 16779
rect 17233 16745 17267 16779
rect 27077 16745 27111 16779
rect 27721 16745 27755 16779
rect 23673 16677 23707 16711
rect 1685 16609 1719 16643
rect 3801 16609 3835 16643
rect 5733 16609 5767 16643
rect 5917 16609 5951 16643
rect 6561 16609 6595 16643
rect 7481 16609 7515 16643
rect 8217 16609 8251 16643
rect 9873 16609 9907 16643
rect 11161 16609 11195 16643
rect 14105 16609 14139 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 16865 16609 16899 16643
rect 17601 16609 17635 16643
rect 19533 16609 19567 16643
rect 20085 16609 20119 16643
rect 20821 16609 20855 16643
rect 25053 16609 25087 16643
rect 27997 16609 28031 16643
rect 3157 16541 3191 16575
rect 3617 16541 3651 16575
rect 4537 16541 4571 16575
rect 6469 16541 6503 16575
rect 7297 16541 7331 16575
rect 8033 16541 8067 16575
rect 8953 16541 8987 16575
rect 9689 16541 9723 16575
rect 10885 16541 10919 16575
rect 11345 16541 11379 16575
rect 12173 16541 12207 16575
rect 13277 16541 13311 16575
rect 13737 16541 13771 16575
rect 14361 16541 14395 16575
rect 16681 16541 16715 16575
rect 19349 16541 19383 16575
rect 20269 16541 20303 16575
rect 21005 16541 21039 16575
rect 21557 16541 21591 16575
rect 21925 16541 21959 16575
rect 22192 16541 22226 16575
rect 23581 16557 23615 16591
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 26985 16541 27019 16575
rect 1952 16473 1986 16507
rect 4445 16473 4479 16507
rect 6377 16473 6411 16507
rect 17868 16473 17902 16507
rect 25237 16473 25271 16507
rect 26893 16473 26927 16507
rect 27445 16473 27479 16507
rect 3433 16405 3467 16439
rect 7941 16405 7975 16439
rect 8677 16405 8711 16439
rect 18981 16405 19015 16439
rect 19993 16405 20027 16439
rect 20729 16405 20763 16439
rect 21465 16405 21499 16439
rect 21649 16405 21683 16439
rect 23305 16405 23339 16439
rect 23397 16405 23431 16439
rect 24593 16405 24627 16439
rect 28549 16405 28583 16439
rect 2789 16201 2823 16235
rect 3985 16201 4019 16235
rect 9873 16201 9907 16235
rect 10609 16201 10643 16235
rect 12817 16201 12851 16235
rect 13553 16201 13587 16235
rect 14105 16201 14139 16235
rect 14657 16201 14691 16235
rect 17417 16201 17451 16235
rect 19073 16201 19107 16235
rect 19533 16201 19567 16235
rect 21373 16201 21407 16235
rect 25053 16201 25087 16235
rect 26249 16201 26283 16235
rect 26985 16201 27019 16235
rect 3525 16133 3559 16167
rect 22569 16133 22603 16167
rect 1409 16065 1443 16099
rect 1676 16065 1710 16099
rect 2973 16065 3007 16099
rect 3893 16065 3927 16099
rect 4169 16065 4203 16099
rect 4537 16065 4571 16099
rect 6377 16065 6411 16099
rect 7573 16065 7607 16099
rect 8861 16065 8895 16099
rect 8953 16065 8987 16099
rect 9045 16065 9079 16099
rect 9413 16065 9447 16099
rect 9965 16065 9999 16099
rect 11069 16065 11103 16099
rect 11345 16065 11379 16099
rect 11805 16065 11839 16099
rect 11897 16065 11931 16099
rect 12173 16065 12207 16099
rect 12909 16065 12943 16099
rect 13829 16065 13863 16099
rect 14289 16065 14323 16099
rect 14541 16065 14575 16099
rect 14841 16065 14875 16099
rect 15117 16065 15151 16099
rect 15393 16065 15427 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 15945 16065 15979 16099
rect 16773 16065 16807 16099
rect 16957 16065 16991 16099
rect 17693 16065 17727 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 19993 16065 20027 16099
rect 20361 16065 20395 16099
rect 20545 16065 20579 16099
rect 21089 16055 21123 16089
rect 21557 16065 21591 16099
rect 22017 16065 22051 16099
rect 23673 16065 23707 16099
rect 24593 16065 24627 16099
rect 25145 16065 25179 16099
rect 26065 16065 26099 16099
rect 26341 16065 26375 16099
rect 26617 16065 26651 16099
rect 27177 16065 27211 16099
rect 27353 16065 27387 16099
rect 27905 16065 27939 16099
rect 4629 15997 4663 16031
rect 4813 15997 4847 16031
rect 6561 15997 6595 16031
rect 7757 15997 7791 16031
rect 9229 15997 9263 16031
rect 10149 15997 10183 16031
rect 12357 15997 12391 16031
rect 13093 15997 13127 16031
rect 15761 15997 15795 16031
rect 18245 15997 18279 16031
rect 20085 15997 20119 16031
rect 22845 15997 22879 16031
rect 23489 15997 23523 16031
rect 24409 15997 24443 16031
rect 25329 15997 25363 16031
rect 27721 15997 27755 16031
rect 3709 15929 3743 15963
rect 4353 15929 4387 15963
rect 11161 15929 11195 15963
rect 11989 15929 12023 15963
rect 15209 15929 15243 15963
rect 20729 15929 20763 15963
rect 21189 15929 21223 15963
rect 26709 15929 26743 15963
rect 5181 15861 5215 15895
rect 6745 15861 6779 15895
rect 7941 15861 7975 15895
rect 8677 15861 8711 15895
rect 10885 15861 10919 15895
rect 11621 15861 11655 15895
rect 13921 15861 13955 15895
rect 14381 15861 14415 15895
rect 14933 15861 14967 15895
rect 16405 15861 16439 15895
rect 23397 15861 23431 15895
rect 24041 15861 24075 15895
rect 25789 15861 25823 15895
rect 26433 15861 26467 15895
rect 27537 15861 27571 15895
rect 28089 15861 28123 15895
rect 2237 15657 2271 15691
rect 5181 15657 5215 15691
rect 6653 15657 6687 15691
rect 8493 15657 8527 15691
rect 9321 15657 9355 15691
rect 17233 15657 17267 15691
rect 21281 15657 21315 15691
rect 22293 15657 22327 15691
rect 24041 15657 24075 15691
rect 24869 15657 24903 15691
rect 25789 15657 25823 15691
rect 26893 15657 26927 15691
rect 28365 15657 28399 15691
rect 3433 15589 3467 15623
rect 13921 15589 13955 15623
rect 27997 15589 28031 15623
rect 5273 15521 5307 15555
rect 6009 15521 6043 15555
rect 6837 15521 6871 15555
rect 7481 15521 7515 15555
rect 7941 15521 7975 15555
rect 10057 15521 10091 15555
rect 12541 15521 12575 15555
rect 17049 15521 17083 15555
rect 18153 15521 18187 15555
rect 18337 15521 18371 15555
rect 18981 15521 19015 15555
rect 20177 15521 20211 15555
rect 20361 15521 20395 15555
rect 20913 15521 20947 15555
rect 21097 15521 21131 15555
rect 23397 15521 23431 15555
rect 25145 15521 25179 15555
rect 25329 15521 25363 15555
rect 26433 15521 26467 15555
rect 26985 15521 27019 15555
rect 27813 15521 27847 15555
rect 1685 15453 1719 15487
rect 2329 15453 2363 15487
rect 3341 15453 3375 15487
rect 3617 15453 3651 15487
rect 3985 15453 4019 15487
rect 4445 15453 4479 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 5457 15453 5491 15487
rect 6193 15453 6227 15487
rect 8401 15453 8435 15487
rect 9505 15453 9539 15487
rect 9781 15453 9815 15487
rect 10977 15453 11011 15487
rect 14105 15453 14139 15487
rect 16865 15453 16899 15487
rect 17785 15453 17819 15487
rect 18889 15453 18923 15487
rect 19441 15453 19475 15487
rect 21649 15453 21683 15487
rect 22385 15453 22419 15487
rect 22569 15453 22603 15487
rect 23305 15453 23339 15487
rect 23581 15453 23615 15487
rect 24501 15453 24535 15487
rect 25053 15453 25087 15487
rect 25881 15453 25915 15487
rect 26249 15453 26283 15487
rect 27169 15453 27203 15487
rect 27721 15453 27755 15487
rect 28181 15453 28215 15487
rect 28273 15453 28307 15487
rect 6929 15385 6963 15419
rect 7665 15385 7699 15419
rect 7757 15385 7791 15419
rect 12808 15385 12842 15419
rect 14749 15385 14783 15419
rect 15025 15385 15059 15419
rect 25973 15385 26007 15419
rect 2973 15317 3007 15351
rect 3157 15317 3191 15351
rect 4077 15317 4111 15351
rect 4261 15317 4295 15351
rect 5917 15317 5951 15351
rect 10793 15317 10827 15351
rect 16313 15317 16347 15351
rect 17601 15317 17635 15351
rect 18797 15317 18831 15351
rect 20085 15317 20119 15351
rect 20821 15317 20855 15351
rect 23029 15317 23063 15351
rect 23121 15317 23155 15351
rect 24593 15317 24627 15351
rect 27629 15317 27663 15351
rect 2789 15113 2823 15147
rect 4813 15113 4847 15147
rect 5273 15113 5307 15147
rect 6009 15113 6043 15147
rect 6377 15113 6411 15147
rect 6745 15113 6779 15147
rect 7021 15113 7055 15147
rect 7481 15113 7515 15147
rect 10425 15113 10459 15147
rect 16681 15113 16715 15147
rect 20545 15113 20579 15147
rect 21373 15113 21407 15147
rect 26709 15113 26743 15147
rect 28365 15113 28399 15147
rect 1676 15045 1710 15079
rect 3065 14977 3099 15011
rect 4445 14977 4479 15011
rect 4721 14977 4755 15011
rect 5457 14977 5491 15011
rect 5917 14977 5951 15011
rect 6193 14977 6227 15011
rect 6653 14977 6687 15011
rect 7205 14977 7239 15011
rect 7389 14977 7423 15011
rect 7849 14977 7883 15011
rect 8033 14977 8067 15011
rect 8309 14977 8343 15011
rect 10609 14977 10643 15011
rect 10885 14977 10919 15011
rect 12081 14977 12115 15011
rect 12348 14977 12382 15011
rect 13737 14977 13771 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 17509 14977 17543 15011
rect 18153 14977 18187 15011
rect 18981 14977 19015 15011
rect 20637 14977 20671 15011
rect 21557 14977 21591 15011
rect 21833 14977 21867 15011
rect 22569 14977 22603 15011
rect 22836 14977 22870 15011
rect 24225 14977 24259 15011
rect 25881 14977 25915 15011
rect 27169 14977 27203 15011
rect 27445 14977 27479 15011
rect 27721 14977 27755 15011
rect 27997 14977 28031 15011
rect 28273 14977 28307 15011
rect 28549 14977 28583 15011
rect 1409 14909 1443 14943
rect 2881 14909 2915 14943
rect 3709 14909 3743 14943
rect 3893 14909 3927 14943
rect 4537 14909 4571 14943
rect 8493 14909 8527 14943
rect 10057 14909 10091 14943
rect 14013 14909 14047 14943
rect 14197 14909 14231 14943
rect 14565 14909 14599 14943
rect 15945 14909 15979 14943
rect 17325 14909 17359 14943
rect 18337 14909 18371 14943
rect 19165 14909 19199 14943
rect 19901 14909 19935 14943
rect 20085 14909 20119 14943
rect 20821 14909 20855 14943
rect 22017 14909 22051 14943
rect 24409 14909 24443 14943
rect 24961 14909 24995 14943
rect 25145 14909 25179 14943
rect 26065 14909 26099 14943
rect 26249 14909 26283 14943
rect 5733 14841 5767 14875
rect 7665 14841 7699 14875
rect 8217 14841 8251 14875
rect 13921 14841 13955 14875
rect 17141 14841 17175 14875
rect 25697 14841 25731 14875
rect 27261 14841 27295 14875
rect 27537 14841 27571 14875
rect 3249 14773 3283 14807
rect 4353 14773 4387 14807
rect 10701 14773 10735 14807
rect 13461 14773 13495 14807
rect 17969 14773 18003 14807
rect 18521 14773 18555 14807
rect 19625 14773 19659 14807
rect 21005 14773 21039 14807
rect 22477 14773 22511 14807
rect 23949 14773 23983 14807
rect 24869 14773 24903 14807
rect 25329 14773 25363 14807
rect 26985 14773 27019 14807
rect 27813 14773 27847 14807
rect 28089 14773 28123 14807
rect 2329 14569 2363 14603
rect 3157 14569 3191 14603
rect 3249 14569 3283 14603
rect 4353 14569 4387 14603
rect 8401 14569 8435 14603
rect 12081 14569 12115 14603
rect 13001 14569 13035 14603
rect 13921 14569 13955 14603
rect 16589 14569 16623 14603
rect 17141 14569 17175 14603
rect 17969 14569 18003 14603
rect 18521 14569 18555 14603
rect 19349 14569 19383 14603
rect 19901 14569 19935 14603
rect 20177 14569 20211 14603
rect 20453 14569 20487 14603
rect 22477 14569 22511 14603
rect 22845 14569 22879 14603
rect 25053 14569 25087 14603
rect 26617 14569 26651 14603
rect 27445 14569 27479 14603
rect 4537 14501 4571 14535
rect 19625 14501 19659 14535
rect 20729 14501 20763 14535
rect 24041 14501 24075 14535
rect 27353 14501 27387 14535
rect 28089 14501 28123 14535
rect 2053 14433 2087 14467
rect 2513 14433 2547 14467
rect 2697 14433 2731 14467
rect 3801 14433 3835 14467
rect 3985 14433 4019 14467
rect 10425 14433 10459 14467
rect 10609 14433 10643 14467
rect 12449 14433 12483 14467
rect 14565 14433 14599 14467
rect 16221 14433 16255 14467
rect 17509 14433 17543 14467
rect 21189 14433 21223 14467
rect 21741 14433 21775 14467
rect 25237 14433 25271 14467
rect 27721 14433 27755 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2237 14365 2271 14399
rect 3433 14365 3467 14399
rect 4721 14365 4755 14399
rect 5089 14365 5123 14399
rect 5273 14365 5307 14399
rect 6929 14365 6963 14399
rect 8585 14365 8619 14399
rect 8953 14365 8987 14399
rect 11161 14365 11195 14399
rect 11345 14365 11379 14399
rect 11805 14365 11839 14399
rect 11997 14365 12031 14399
rect 12265 14365 12299 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 14105 14365 14139 14399
rect 16037 14365 16071 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 17693 14365 17727 14399
rect 18429 14365 18463 14399
rect 18705 14365 18739 14399
rect 19257 14365 19291 14399
rect 19809 14365 19843 14399
rect 20085 14365 20119 14399
rect 20361 14365 20395 14399
rect 20637 14365 20671 14399
rect 20913 14365 20947 14399
rect 21005 14365 21039 14399
rect 21925 14365 21959 14399
rect 22661 14365 22695 14399
rect 22753 14365 22787 14399
rect 24225 14365 24259 14399
rect 24961 14365 24995 14399
rect 26709 14365 26743 14399
rect 26893 14365 26927 14399
rect 27629 14365 27663 14399
rect 27905 14365 27939 14399
rect 5529 14297 5563 14331
rect 7196 14297 7230 14331
rect 9220 14297 9254 14331
rect 14289 14297 14323 14331
rect 24501 14297 24535 14331
rect 25504 14297 25538 14331
rect 1777 14229 1811 14263
rect 4905 14229 4939 14263
rect 6653 14229 6687 14263
rect 8309 14229 8343 14263
rect 10333 14229 10367 14263
rect 11069 14229 11103 14263
rect 12909 14229 12943 14263
rect 18245 14229 18279 14263
rect 21649 14229 21683 14263
rect 22385 14229 22419 14263
rect 24593 14229 24627 14263
rect 2789 14025 2823 14059
rect 6653 14025 6687 14059
rect 7573 14025 7607 14059
rect 8125 14025 8159 14059
rect 10885 14025 10919 14059
rect 12173 14025 12207 14059
rect 12265 14025 12299 14059
rect 13185 14025 13219 14059
rect 14657 14025 14691 14059
rect 15117 14025 15151 14059
rect 16129 14025 16163 14059
rect 16221 14025 16255 14059
rect 17601 14025 17635 14059
rect 18061 14025 18095 14059
rect 21097 14025 21131 14059
rect 21465 14025 21499 14059
rect 28457 14025 28491 14059
rect 6469 13957 6503 13991
rect 17509 13957 17543 13991
rect 19892 13957 19926 13991
rect 24133 13957 24167 13991
rect 1676 13889 1710 13923
rect 3617 13889 3651 13923
rect 4077 13889 4111 13923
rect 4445 13889 4479 13923
rect 6009 13889 6043 13923
rect 6377 13889 6411 13923
rect 6837 13889 6871 13923
rect 7849 13889 7883 13923
rect 8033 13889 8067 13923
rect 10241 13889 10275 13923
rect 11345 13889 11379 13923
rect 12449 13889 12483 13923
rect 13277 13889 13311 13923
rect 13544 13889 13578 13923
rect 14933 13889 14967 13923
rect 15025 13889 15059 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 16405 13889 16439 13923
rect 17969 13889 18003 13923
rect 18521 13889 18555 13923
rect 18613 13889 18647 13923
rect 18797 13889 18831 13923
rect 19533 13889 19567 13923
rect 19625 13889 19659 13923
rect 21281 13889 21315 13923
rect 21373 13889 21407 13923
rect 22201 13889 22235 13923
rect 23029 13889 23063 13923
rect 23121 13889 23155 13923
rect 23489 13889 23523 13923
rect 24593 13889 24627 13923
rect 25237 13889 25271 13923
rect 25881 13889 25915 13923
rect 26341 13889 26375 13923
rect 26433 13889 26467 13923
rect 27077 13889 27111 13923
rect 27169 13889 27203 13923
rect 27537 13889 27571 13923
rect 28273 13889 28307 13923
rect 28365 13889 28399 13923
rect 1409 13821 1443 13855
rect 2881 13821 2915 13855
rect 3065 13821 3099 13855
rect 3709 13821 3743 13855
rect 4261 13821 4295 13855
rect 5089 13821 5123 13855
rect 5273 13821 5307 13855
rect 7021 13821 7055 13855
rect 8309 13821 8343 13855
rect 8493 13821 8527 13855
rect 10057 13821 10091 13855
rect 10425 13821 10459 13855
rect 11529 13821 11563 13855
rect 11713 13821 11747 13855
rect 12541 13821 12575 13855
rect 12725 13821 12759 13855
rect 23305 13821 23339 13855
rect 24409 13821 24443 13855
rect 27353 13821 27387 13855
rect 27997 13821 28031 13855
rect 11161 13753 11195 13787
rect 14749 13753 14783 13787
rect 19349 13753 19383 13787
rect 21005 13753 21039 13787
rect 28089 13753 28123 13787
rect 3249 13685 3283 13719
rect 3893 13685 3927 13719
rect 4813 13685 4847 13719
rect 5733 13685 5767 13719
rect 6101 13685 6135 13719
rect 7665 13685 7699 13719
rect 18337 13685 18371 13719
rect 19257 13685 19291 13719
rect 22017 13685 22051 13719
rect 23673 13685 23707 13719
rect 25053 13685 25087 13719
rect 25789 13685 25823 13719
rect 25973 13685 26007 13719
rect 26157 13685 26191 13719
rect 26525 13685 26559 13719
rect 3893 13481 3927 13515
rect 4813 13481 4847 13515
rect 5549 13481 5583 13515
rect 6009 13481 6043 13515
rect 7113 13481 7147 13515
rect 7941 13481 7975 13515
rect 8309 13481 8343 13515
rect 9965 13481 9999 13515
rect 12725 13481 12759 13515
rect 13737 13481 13771 13515
rect 16037 13481 16071 13515
rect 19625 13481 19659 13515
rect 24777 13481 24811 13515
rect 25513 13481 25547 13515
rect 1777 13413 1811 13447
rect 3433 13413 3467 13447
rect 7389 13413 7423 13447
rect 9137 13413 9171 13447
rect 16681 13413 16715 13447
rect 16957 13413 16991 13447
rect 18061 13413 18095 13447
rect 18521 13413 18555 13447
rect 22937 13413 22971 13447
rect 23397 13413 23431 13447
rect 2237 13345 2271 13379
rect 2697 13345 2731 13379
rect 4169 13345 4203 13379
rect 5825 13345 5859 13379
rect 6469 13345 6503 13379
rect 7757 13345 7791 13379
rect 9321 13345 9355 13379
rect 10149 13345 10183 13379
rect 11621 13345 11655 13379
rect 11805 13345 11839 13379
rect 13185 13345 13219 13379
rect 14473 13345 14507 13379
rect 14841 13345 14875 13379
rect 15577 13345 15611 13379
rect 16221 13345 16255 13379
rect 17417 13345 17451 13379
rect 17601 13345 17635 13379
rect 18981 13345 19015 13379
rect 19441 13345 19475 13379
rect 20729 13345 20763 13379
rect 22293 13345 22327 13379
rect 24133 13345 24167 13379
rect 24593 13345 24627 13379
rect 25145 13345 25179 13379
rect 25329 13345 25363 13379
rect 27169 13345 27203 13379
rect 1961 13277 1995 13311
rect 2053 13277 2087 13311
rect 2881 13277 2915 13311
rect 3801 13277 3835 13311
rect 4353 13277 4387 13311
rect 4905 13277 4939 13311
rect 5641 13277 5675 13311
rect 6653 13277 6687 13311
rect 7297 13277 7331 13311
rect 7573 13277 7607 13311
rect 8493 13277 8527 13311
rect 8769 13277 8803 13311
rect 9045 13277 9079 13311
rect 10793 13277 10827 13311
rect 10977 13277 11011 13311
rect 12357 13277 12391 13311
rect 12541 13277 12575 13311
rect 14289 13277 14323 13311
rect 14381 13277 14415 13311
rect 14657 13277 14691 13311
rect 15301 13277 15335 13311
rect 15393 13277 15427 13311
rect 16129 13277 16163 13311
rect 16865 13277 16899 13311
rect 17141 13277 17175 13311
rect 18153 13277 18187 13311
rect 18337 13277 18371 13311
rect 18889 13277 18923 13311
rect 19257 13277 19291 13311
rect 20913 13277 20947 13311
rect 21465 13277 21499 13311
rect 22477 13277 22511 13311
rect 23029 13277 23063 13311
rect 23213 13277 23247 13311
rect 23949 13277 23983 13311
rect 24041 13277 24075 13311
rect 24409 13277 24443 13311
rect 25881 13277 25915 13311
rect 26709 13277 26743 13311
rect 1501 13209 1535 13243
rect 22109 13209 22143 13243
rect 26893 13209 26927 13243
rect 1593 13141 1627 13175
rect 8585 13141 8619 13175
rect 10701 13141 10735 13175
rect 11437 13141 11471 13175
rect 12265 13141 12299 13175
rect 14105 13141 14139 13175
rect 19993 13141 20027 13175
rect 21373 13141 21407 13175
rect 23765 13141 23799 13175
rect 26525 13141 26559 13175
rect 2973 12937 3007 12971
rect 3985 12937 4019 12971
rect 6009 12937 6043 12971
rect 6561 12937 6595 12971
rect 8125 12937 8159 12971
rect 8953 12937 8987 12971
rect 9229 12937 9263 12971
rect 10793 12937 10827 12971
rect 12173 12937 12207 12971
rect 12265 12937 12299 12971
rect 12909 12937 12943 12971
rect 13093 12937 13127 12971
rect 13461 12937 13495 12971
rect 13645 12937 13679 12971
rect 15301 12937 15335 12971
rect 15485 12937 15519 12971
rect 17325 12937 17359 12971
rect 17601 12937 17635 12971
rect 21557 12937 21591 12971
rect 22385 12937 22419 12971
rect 22753 12937 22787 12971
rect 24593 12937 24627 12971
rect 27629 12937 27663 12971
rect 28365 12937 28399 12971
rect 25412 12869 25446 12903
rect 1860 12801 1894 12835
rect 3709 12801 3743 12835
rect 3893 12801 3927 12835
rect 4261 12801 4295 12835
rect 4353 12801 4387 12835
rect 4721 12801 4755 12835
rect 6193 12801 6227 12835
rect 6469 12801 6503 12835
rect 6929 12801 6963 12835
rect 7665 12801 7699 12835
rect 8493 12801 8527 12835
rect 9413 12801 9447 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10701 12801 10735 12835
rect 10977 12801 11011 12835
rect 11345 12801 11379 12835
rect 12449 12801 12483 12835
rect 12725 12801 12759 12835
rect 12817 12801 12851 12835
rect 13277 12801 13311 12835
rect 13369 12801 13403 12835
rect 13837 12801 13871 12835
rect 14841 12801 14875 12835
rect 15669 12801 15703 12835
rect 16037 12801 16071 12835
rect 17509 12801 17543 12835
rect 17969 12801 18003 12835
rect 19073 12801 19107 12835
rect 20545 12801 20579 12835
rect 21465 12801 21499 12835
rect 22017 12801 22051 12835
rect 22293 12801 22327 12835
rect 22569 12801 22603 12835
rect 22661 12801 22695 12835
rect 23121 12801 23155 12835
rect 23213 12801 23247 12835
rect 23397 12801 23431 12835
rect 23949 12801 23983 12835
rect 24869 12801 24903 12835
rect 26617 12801 26651 12835
rect 27905 12801 27939 12835
rect 1593 12733 1627 12767
rect 3065 12733 3099 12767
rect 4537 12733 4571 12767
rect 5273 12733 5307 12767
rect 5457 12733 5491 12767
rect 6745 12733 6779 12767
rect 7481 12733 7515 12767
rect 8309 12733 8343 12767
rect 10057 12733 10091 12767
rect 10241 12733 10275 12767
rect 11529 12733 11563 12767
rect 11713 12733 11747 12767
rect 14657 12733 14691 12767
rect 16681 12733 16715 12767
rect 16865 12733 16899 12767
rect 18337 12733 18371 12767
rect 18521 12733 18555 12767
rect 19257 12733 19291 12767
rect 19809 12733 19843 12767
rect 19993 12733 20027 12767
rect 20729 12733 20763 12767
rect 24133 12733 24167 12767
rect 25145 12733 25179 12767
rect 27077 12733 27111 12767
rect 27721 12733 27755 12767
rect 9597 12665 9631 12699
rect 11161 12665 11195 12699
rect 15853 12665 15887 12699
rect 18981 12665 19015 12699
rect 19441 12665 19475 12699
rect 23673 12665 23707 12699
rect 24685 12665 24719 12699
rect 26525 12665 26559 12699
rect 5181 12597 5215 12631
rect 5641 12597 5675 12631
rect 7389 12597 7423 12631
rect 9873 12597 9907 12631
rect 12541 12597 12575 12631
rect 17785 12597 17819 12631
rect 20453 12597 20487 12631
rect 20913 12597 20947 12631
rect 21833 12597 21867 12631
rect 22109 12597 22143 12631
rect 22937 12597 22971 12631
rect 26709 12597 26743 12631
rect 2789 12393 2823 12427
rect 5181 12393 5215 12427
rect 6101 12393 6135 12427
rect 7389 12393 7423 12427
rect 8585 12393 8619 12427
rect 9321 12393 9355 12427
rect 11069 12393 11103 12427
rect 12817 12393 12851 12427
rect 15301 12393 15335 12427
rect 17785 12393 17819 12427
rect 18797 12393 18831 12427
rect 19625 12393 19659 12427
rect 20085 12393 20119 12427
rect 23857 12393 23891 12427
rect 25053 12393 25087 12427
rect 6469 12325 6503 12359
rect 7573 12325 7607 12359
rect 16037 12325 16071 12359
rect 16497 12325 16531 12359
rect 21373 12325 21407 12359
rect 25329 12325 25363 12359
rect 28089 12325 28123 12359
rect 6929 12257 6963 12291
rect 8309 12257 8343 12291
rect 8953 12257 8987 12291
rect 11897 12257 11931 12291
rect 14473 12257 14507 12291
rect 14841 12257 14875 12291
rect 16129 12257 16163 12291
rect 20821 12257 20855 12291
rect 21005 12257 21039 12291
rect 21741 12257 21775 12291
rect 25605 12257 25639 12291
rect 25789 12257 25823 12291
rect 26801 12257 26835 12291
rect 27721 12257 27755 12291
rect 27905 12257 27939 12291
rect 1409 12189 1443 12223
rect 2973 12189 3007 12223
rect 3525 12189 3559 12223
rect 3801 12189 3835 12223
rect 5365 12189 5399 12223
rect 6285 12189 6319 12223
rect 6653 12189 6687 12223
rect 6745 12189 6779 12223
rect 7757 12189 7791 12223
rect 7849 12189 7883 12223
rect 8125 12189 8159 12223
rect 9137 12189 9171 12223
rect 9689 12189 9723 12223
rect 9956 12189 9990 12223
rect 11437 12189 11471 12223
rect 11713 12189 11747 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14105 12189 14139 12223
rect 14381 12189 14415 12223
rect 14657 12189 14691 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 16313 12189 16347 12223
rect 17969 12189 18003 12223
rect 18705 12189 18739 12223
rect 19533 12189 19567 12223
rect 19993 12189 20027 12223
rect 20269 12189 20303 12223
rect 22845 12189 22879 12223
rect 23305 12189 23339 12223
rect 23581 12189 23615 12223
rect 24041 12189 24075 12223
rect 24501 12189 24535 12223
rect 24777 12189 24811 12223
rect 25237 12189 25271 12223
rect 25513 12189 25547 12223
rect 1676 12121 1710 12155
rect 4068 12121 4102 12155
rect 6009 12121 6043 12155
rect 7941 12121 7975 12155
rect 13921 12121 13955 12155
rect 21833 12121 21867 12155
rect 22753 12121 22787 12155
rect 11253 12053 11287 12087
rect 12357 12053 12391 12087
rect 14197 12053 14231 12087
rect 19809 12053 19843 12087
rect 23029 12053 23063 12087
rect 23397 12053 23431 12087
rect 23673 12053 23707 12087
rect 24593 12053 24627 12087
rect 24869 12053 24903 12087
rect 4721 11849 4755 11883
rect 7113 11849 7147 11883
rect 10701 11849 10735 11883
rect 12173 11849 12207 11883
rect 12449 11849 12483 11883
rect 12817 11849 12851 11883
rect 13093 11849 13127 11883
rect 13553 11849 13587 11883
rect 14749 11849 14783 11883
rect 15853 11849 15887 11883
rect 16037 11849 16071 11883
rect 16313 11849 16347 11883
rect 24409 11849 24443 11883
rect 26065 11849 26099 11883
rect 28181 11849 28215 11883
rect 28365 11849 28399 11883
rect 2053 11781 2087 11815
rect 20536 11781 20570 11815
rect 21925 11781 21959 11815
rect 22017 11781 22051 11815
rect 24952 11781 24986 11815
rect 3985 11713 4019 11747
rect 4077 11713 4111 11747
rect 5080 11713 5114 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 7757 11713 7791 11747
rect 7941 11713 7975 11747
rect 8677 11713 8711 11747
rect 9689 11713 9723 11747
rect 10885 11713 10919 11747
rect 11713 11713 11747 11747
rect 12633 11713 12667 11747
rect 12725 11713 12759 11747
rect 13277 11713 13311 11747
rect 13737 11713 13771 11747
rect 14289 11713 14323 11747
rect 15761 11713 15795 11747
rect 16221 11713 16255 11747
rect 16497 11713 16531 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 20177 11713 20211 11747
rect 23213 11713 23247 11747
rect 23489 11713 23523 11747
rect 24593 11713 24627 11747
rect 27169 11713 27203 11747
rect 27445 11713 27479 11747
rect 27537 11713 27571 11747
rect 28273 11713 28307 11747
rect 1593 11645 1627 11679
rect 1961 11645 1995 11679
rect 2973 11645 3007 11679
rect 3065 11645 3099 11679
rect 3249 11645 3283 11679
rect 4813 11645 4847 11679
rect 6377 11645 6411 11679
rect 10057 11645 10091 11679
rect 11529 11645 11563 11679
rect 14105 11645 14139 11679
rect 20269 11645 20303 11679
rect 22753 11645 22787 11679
rect 23673 11645 23707 11679
rect 24685 11645 24719 11679
rect 26249 11645 26283 11679
rect 27721 11645 27755 11679
rect 19993 11577 20027 11611
rect 26985 11577 27019 11611
rect 3433 11509 3467 11543
rect 3801 11509 3835 11543
rect 6193 11509 6227 11543
rect 7573 11509 7607 11543
rect 7849 11509 7883 11543
rect 8769 11509 8803 11543
rect 18613 11509 18647 11543
rect 21649 11509 21683 11543
rect 23029 11509 23063 11543
rect 24133 11509 24167 11543
rect 26801 11509 26835 11543
rect 27261 11509 27295 11543
rect 2053 11305 2087 11339
rect 2513 11305 2547 11339
rect 2697 11305 2731 11339
rect 5457 11305 5491 11339
rect 9413 11305 9447 11339
rect 11529 11305 11563 11339
rect 11989 11305 12023 11339
rect 21005 11305 21039 11339
rect 22661 11305 22695 11339
rect 23029 11305 23063 11339
rect 24133 11305 24167 11339
rect 26893 11305 26927 11339
rect 2145 11237 2179 11271
rect 3617 11237 3651 11271
rect 4721 11237 4755 11271
rect 5181 11237 5215 11271
rect 8309 11237 8343 11271
rect 8585 11237 8619 11271
rect 9873 11237 9907 11271
rect 10333 11237 10367 11271
rect 14749 11237 14783 11271
rect 26617 11237 26651 11271
rect 3157 11169 3191 11203
rect 4169 11169 4203 11203
rect 4537 11169 4571 11203
rect 9045 11169 9079 11203
rect 9229 11169 9263 11203
rect 11621 11169 11655 11203
rect 11805 11169 11839 11203
rect 17509 11169 17543 11203
rect 19441 11169 19475 11203
rect 19625 11169 19659 11203
rect 25237 11169 25271 11203
rect 27169 11169 27203 11203
rect 1869 11101 1903 11135
rect 2329 11101 2363 11135
rect 2421 11101 2455 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4353 11101 4387 11135
rect 5365 11101 5399 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 6101 11101 6135 11135
rect 7573 11101 7607 11135
rect 8493 11101 8527 11135
rect 8769 11101 8803 11135
rect 10057 11101 10091 11135
rect 10517 11101 10551 11135
rect 10885 11101 10919 11135
rect 11069 11101 11103 11135
rect 12541 11101 12575 11135
rect 12817 11101 12851 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 15301 11101 15335 11135
rect 16037 11101 16071 11135
rect 17693 11101 17727 11135
rect 18245 11101 18279 11135
rect 18889 11101 18923 11135
rect 19349 11101 19383 11135
rect 21097 11101 21131 11135
rect 21833 11101 21867 11135
rect 22569 11101 22603 11135
rect 23213 11101 23247 11135
rect 23489 11101 23523 11135
rect 23673 11101 23707 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 27077 11101 27111 11135
rect 27436 11101 27470 11135
rect 15577 11033 15611 11067
rect 19892 11033 19926 11067
rect 22477 11033 22511 11067
rect 25504 11033 25538 11067
rect 3801 10965 3835 10999
rect 7757 10965 7791 10999
rect 15853 10965 15887 10999
rect 18153 10965 18187 10999
rect 18337 10965 18371 10999
rect 18705 10965 18739 10999
rect 21741 10965 21775 10999
rect 25053 10965 25087 10999
rect 28549 10965 28583 10999
rect 2605 10761 2639 10795
rect 5641 10761 5675 10795
rect 7757 10761 7791 10795
rect 10425 10761 10459 10795
rect 10977 10761 11011 10795
rect 11529 10761 11563 10795
rect 13645 10761 13679 10795
rect 13921 10761 13955 10795
rect 15117 10761 15151 10795
rect 15209 10761 15243 10795
rect 17693 10761 17727 10795
rect 24225 10761 24259 10795
rect 27261 10761 27295 10795
rect 13369 10693 13403 10727
rect 20444 10693 20478 10727
rect 23121 10693 23155 10727
rect 24593 10693 24627 10727
rect 25145 10693 25179 10727
rect 25596 10693 25630 10727
rect 28181 10693 28215 10727
rect 1593 10625 1627 10659
rect 1869 10625 1903 10659
rect 2697 10625 2731 10659
rect 2964 10625 2998 10659
rect 4169 10625 4203 10659
rect 4436 10625 4470 10659
rect 5825 10625 5859 10659
rect 6101 10625 6135 10659
rect 6644 10625 6678 10659
rect 9965 10625 9999 10659
rect 10885 10625 10919 10659
rect 11345 10625 11379 10659
rect 11713 10625 11747 10659
rect 11989 10625 12023 10659
rect 13277 10625 13311 10659
rect 13829 10625 13863 10659
rect 14105 10625 14139 10659
rect 14197 10625 14231 10659
rect 14289 10625 14323 10659
rect 14657 10625 14691 10659
rect 15393 10625 15427 10659
rect 15853 10625 15887 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 17785 10625 17819 10659
rect 19625 10625 19659 10659
rect 22017 10625 22051 10659
rect 22385 10625 22419 10659
rect 22845 10625 22879 10659
rect 23029 10625 23063 10659
rect 24133 10625 24167 10659
rect 27169 10625 27203 10659
rect 27445 10625 27479 10659
rect 28273 10625 28307 10659
rect 1961 10557 1995 10591
rect 2145 10557 2179 10591
rect 6377 10557 6411 10591
rect 7849 10557 7883 10591
rect 8033 10557 8067 10591
rect 8401 10557 8435 10591
rect 9781 10557 9815 10591
rect 11805 10557 11839 10591
rect 12541 10557 12575 10591
rect 12725 10557 12759 10591
rect 14473 10557 14507 10591
rect 15669 10557 15703 10591
rect 17233 10557 17267 10591
rect 18153 10557 18187 10591
rect 20177 10557 20211 10591
rect 23305 10557 23339 10591
rect 23489 10557 23523 10591
rect 23949 10557 23983 10591
rect 24501 10557 24535 10591
rect 25329 10557 25363 10591
rect 27537 10557 27571 10591
rect 1409 10489 1443 10523
rect 1685 10489 1719 10523
rect 5549 10489 5583 10523
rect 11161 10489 11195 10523
rect 21833 10489 21867 10523
rect 22201 10489 22235 10523
rect 22661 10489 22695 10523
rect 4077 10421 4111 10455
rect 5917 10421 5951 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 16037 10421 16071 10455
rect 16773 10421 16807 10455
rect 19809 10421 19843 10455
rect 21557 10421 21591 10455
rect 26709 10421 26743 10455
rect 26985 10421 27019 10455
rect 28365 10421 28399 10455
rect 2329 10217 2363 10251
rect 4905 10217 4939 10251
rect 5457 10217 5491 10251
rect 7849 10217 7883 10251
rect 8309 10217 8343 10251
rect 16037 10217 16071 10251
rect 17601 10217 17635 10251
rect 21189 10217 21223 10251
rect 22293 10217 22327 10251
rect 23305 10217 23339 10251
rect 23673 10217 23707 10251
rect 24777 10217 24811 10251
rect 1593 10149 1627 10183
rect 3157 10149 3191 10183
rect 6653 10149 6687 10183
rect 19073 10149 19107 10183
rect 19625 10149 19659 10183
rect 21373 10149 21407 10183
rect 21925 10149 21959 10183
rect 22937 10149 22971 10183
rect 5181 10081 5215 10115
rect 11529 10081 11563 10115
rect 12357 10081 12391 10115
rect 15577 10081 15611 10115
rect 16221 10081 16255 10115
rect 17969 10081 18003 10115
rect 18613 10081 18647 10115
rect 19257 10081 19291 10115
rect 22661 10081 22695 10115
rect 24593 10081 24627 10115
rect 25237 10081 25271 10115
rect 26157 10081 26191 10115
rect 26341 10081 26375 10115
rect 27077 10081 27111 10115
rect 27813 10081 27847 10115
rect 1409 10013 1443 10047
rect 2513 10013 2547 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3433 10013 3467 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 5089 10013 5123 10047
rect 5365 10013 5399 10047
rect 5641 10013 5675 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 8217 10013 8251 10047
rect 9413 10013 9447 10047
rect 9597 10013 9631 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 11713 10013 11747 10047
rect 12541 10013 12575 10047
rect 13745 10013 13779 10047
rect 15393 10013 15427 10047
rect 16129 10013 16163 10047
rect 17417 10013 17451 10047
rect 17509 10013 17543 10047
rect 17877 10013 17911 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 19441 10013 19475 10047
rect 20177 10013 20211 10047
rect 21097 10013 21131 10047
rect 21557 10013 21591 10047
rect 21649 10013 21683 10047
rect 22109 10013 22143 10047
rect 22201 10013 22235 10047
rect 22477 10013 22511 10047
rect 23213 10013 23247 10047
rect 23857 10013 23891 10047
rect 24133 10013 24167 10047
rect 24409 10013 24443 10047
rect 26525 10013 26559 10047
rect 27997 10013 28031 10047
rect 2605 9945 2639 9979
rect 3525 9945 3559 9979
rect 6377 9945 6411 9979
rect 7297 9945 7331 9979
rect 11161 9945 11195 9979
rect 20729 9945 20763 9979
rect 25329 9945 25363 9979
rect 2881 9877 2915 9911
rect 3985 9877 4019 9911
rect 7021 9877 7055 9911
rect 10057 9877 10091 9911
rect 10149 9877 10183 9911
rect 12173 9877 12207 9911
rect 13001 9877 13035 9911
rect 13553 9877 13587 9911
rect 17233 9877 17267 9911
rect 18153 9877 18187 9911
rect 21833 9877 21867 9911
rect 23949 9877 23983 9911
rect 26985 9877 27019 9911
rect 27721 9877 27755 9911
rect 28457 9877 28491 9911
rect 7205 9673 7239 9707
rect 8861 9673 8895 9707
rect 11805 9673 11839 9707
rect 12357 9673 12391 9707
rect 21833 9673 21867 9707
rect 28181 9673 28215 9707
rect 3065 9605 3099 9639
rect 3893 9605 3927 9639
rect 5273 9605 5307 9639
rect 6101 9605 6135 9639
rect 6561 9605 6595 9639
rect 7665 9605 7699 9639
rect 8585 9605 8619 9639
rect 25421 9605 25455 9639
rect 28089 9605 28123 9639
rect 1593 9537 1627 9571
rect 1869 9537 1903 9571
rect 4721 9537 4755 9571
rect 7389 9537 7423 9571
rect 9045 9537 9079 9571
rect 9137 9537 9171 9571
rect 9505 9537 9539 9571
rect 10977 9537 11011 9571
rect 11713 9537 11747 9571
rect 12173 9537 12207 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 13737 9537 13771 9571
rect 14657 9537 14691 9571
rect 14933 9537 14967 9571
rect 15669 9537 15703 9571
rect 17049 9537 17083 9571
rect 17141 9537 17175 9571
rect 17877 9537 17911 9571
rect 18613 9537 18647 9571
rect 20269 9537 20303 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 20913 9537 20947 9571
rect 21005 9537 21039 9571
rect 21189 9537 21223 9571
rect 21465 9537 21499 9571
rect 22017 9537 22051 9571
rect 22845 9537 22879 9571
rect 23029 9537 23063 9571
rect 23673 9537 23707 9571
rect 24685 9537 24719 9571
rect 25881 9537 25915 9571
rect 26249 9537 26283 9571
rect 26525 9537 26559 9571
rect 26801 9537 26835 9571
rect 26985 9537 27019 9571
rect 27445 9537 27479 9571
rect 28365 9537 28399 9571
rect 2145 9469 2179 9503
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 2973 9469 3007 9503
rect 3801 9469 3835 9503
rect 4537 9469 4571 9503
rect 6469 9469 6503 9503
rect 7573 9469 7607 9503
rect 9689 9469 9723 9503
rect 10241 9469 10275 9503
rect 10425 9469 10459 9503
rect 13001 9469 13035 9503
rect 13185 9469 13219 9503
rect 13921 9469 13955 9503
rect 15117 9469 15151 9503
rect 15853 9469 15887 9503
rect 17325 9469 17359 9503
rect 18061 9469 18095 9503
rect 18797 9469 18831 9503
rect 19349 9469 19383 9503
rect 19533 9469 19567 9503
rect 22109 9469 22143 9503
rect 22293 9469 22327 9503
rect 24501 9469 24535 9503
rect 27629 9469 27663 9503
rect 1409 9401 1443 9435
rect 3525 9401 3559 9435
rect 4353 9401 4387 9435
rect 4905 9401 4939 9435
rect 7021 9401 7055 9435
rect 11989 9401 12023 9435
rect 12633 9401 12667 9435
rect 14473 9401 14507 9435
rect 19257 9401 19291 9435
rect 19993 9401 20027 9435
rect 23213 9401 23247 9435
rect 26065 9401 26099 9435
rect 26617 9401 26651 9435
rect 1685 9333 1719 9367
rect 9229 9333 9263 9367
rect 10149 9333 10183 9367
rect 10609 9333 10643 9367
rect 13645 9333 13679 9367
rect 14105 9333 14139 9367
rect 15485 9333 15519 9367
rect 16037 9333 16071 9367
rect 16865 9333 16899 9367
rect 17785 9333 17819 9367
rect 18245 9333 18279 9367
rect 20085 9333 20119 9367
rect 20453 9333 20487 9367
rect 20729 9333 20763 9367
rect 21281 9333 21315 9367
rect 21649 9333 21683 9367
rect 22753 9333 22787 9367
rect 25697 9333 25731 9367
rect 26341 9333 26375 9367
rect 27077 9333 27111 9367
rect 2789 9129 2823 9163
rect 3525 9129 3559 9163
rect 5365 9129 5399 9163
rect 6285 9129 6319 9163
rect 8401 9129 8435 9163
rect 8585 9129 8619 9163
rect 9781 9129 9815 9163
rect 13829 9129 13863 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 17049 9129 17083 9163
rect 17417 9129 17451 9163
rect 18245 9129 18279 9163
rect 18889 9129 18923 9163
rect 20177 9129 20211 9163
rect 22201 9129 22235 9163
rect 23673 9129 23707 9163
rect 24041 9129 24075 9163
rect 25237 9129 25271 9163
rect 27629 9129 27663 9163
rect 7205 9061 7239 9095
rect 14473 9061 14507 9095
rect 21005 9061 21039 9095
rect 21465 9061 21499 9095
rect 3985 8993 4019 9027
rect 4721 8993 4755 9027
rect 5549 8993 5583 9027
rect 6193 8993 6227 9027
rect 7389 8993 7423 9027
rect 7665 8993 7699 9027
rect 9321 8993 9355 9027
rect 10885 8993 10919 9027
rect 11621 8993 11655 9027
rect 14105 8993 14139 9027
rect 14289 8993 14323 9027
rect 14933 8993 14967 9027
rect 20361 8993 20395 9027
rect 21281 8993 21315 9027
rect 23305 8993 23339 9027
rect 24409 8993 24443 9027
rect 25421 8993 25455 9027
rect 26985 8993 27019 9027
rect 27721 8993 27755 9027
rect 2053 8925 2087 8959
rect 2145 8925 2179 8959
rect 2329 8925 2363 8959
rect 2881 8925 2915 8959
rect 4169 8925 4203 8959
rect 4905 8925 4939 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 8309 8925 8343 8959
rect 8769 8925 8803 8959
rect 9137 8925 9171 8959
rect 9873 8925 9907 8959
rect 11069 8925 11103 8959
rect 11805 8925 11839 8959
rect 13737 8925 13771 8959
rect 14841 8925 14875 8959
rect 15209 8925 15243 8959
rect 15853 8925 15887 8959
rect 16129 8925 16163 8959
rect 16405 8925 16439 8959
rect 16681 8925 16715 8959
rect 16773 8925 16807 8959
rect 17233 8925 17267 8959
rect 17325 8925 17359 8959
rect 17785 8925 17819 8959
rect 17877 8925 17911 8959
rect 18153 8925 18187 8959
rect 18797 8925 18831 8959
rect 19073 8925 19107 8959
rect 19441 8925 19475 8959
rect 19901 8925 19935 8959
rect 20085 8925 20119 8959
rect 20545 8925 20579 8959
rect 21097 8925 21131 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 22569 8925 22603 8959
rect 23489 8925 23523 8959
rect 24225 8925 24259 8959
rect 24593 8925 24627 8959
rect 25145 8925 25179 8959
rect 27169 8925 27203 8959
rect 27905 8925 27939 8959
rect 4629 8857 4663 8891
rect 5641 8857 5675 8891
rect 7481 8857 7515 8891
rect 10609 8857 10643 8891
rect 25688 8857 25722 8891
rect 1869 8789 1903 8823
rect 11529 8789 11563 8823
rect 12265 8789 12299 8823
rect 15945 8789 15979 8823
rect 16221 8789 16255 8823
rect 16497 8789 16531 8823
rect 16957 8789 16991 8823
rect 17601 8789 17635 8823
rect 18061 8789 18095 8823
rect 18613 8789 18647 8823
rect 19625 8789 19659 8823
rect 19717 8789 19751 8823
rect 23213 8789 23247 8823
rect 25053 8789 25087 8823
rect 26801 8789 26835 8823
rect 28365 8789 28399 8823
rect 1685 8585 1719 8619
rect 2145 8585 2179 8619
rect 2421 8585 2455 8619
rect 3617 8585 3651 8619
rect 4721 8585 4755 8619
rect 4905 8585 4939 8619
rect 5641 8585 5675 8619
rect 8033 8585 8067 8619
rect 10885 8585 10919 8619
rect 11161 8585 11195 8619
rect 11621 8585 11655 8619
rect 11805 8585 11839 8619
rect 17969 8585 18003 8619
rect 20453 8585 20487 8619
rect 21005 8585 21039 8619
rect 21281 8585 21315 8619
rect 22477 8585 22511 8619
rect 22661 8585 22695 8619
rect 23857 8585 23891 8619
rect 28457 8585 28491 8619
rect 4537 8517 4571 8551
rect 7389 8517 7423 8551
rect 9781 8517 9815 8551
rect 19165 8517 19199 8551
rect 19993 8517 20027 8551
rect 25053 8517 25087 8551
rect 1593 8449 1627 8483
rect 2053 8449 2087 8483
rect 2329 8449 2363 8483
rect 2605 8449 2639 8483
rect 2697 8449 2731 8483
rect 3157 8449 3191 8483
rect 4077 8449 4111 8483
rect 4629 8449 4663 8483
rect 5089 8449 5123 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 6101 8449 6135 8483
rect 6653 8449 6687 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 9045 8449 9079 8483
rect 9505 8449 9539 8483
rect 10793 8449 10827 8483
rect 11345 8449 11379 8483
rect 11529 8449 11563 8483
rect 11989 8449 12023 8483
rect 13001 8449 13035 8483
rect 14933 8449 14967 8483
rect 15117 8449 15151 8483
rect 15393 8449 15427 8483
rect 16129 8449 16163 8483
rect 16773 8449 16807 8483
rect 17049 8449 17083 8483
rect 17325 8449 17359 8483
rect 18061 8449 18095 8483
rect 18429 8449 18463 8483
rect 20177 8449 20211 8483
rect 20637 8449 20671 8483
rect 20913 8449 20947 8483
rect 21189 8449 21223 8483
rect 21465 8449 21499 8483
rect 22017 8449 22051 8483
rect 22569 8449 22603 8483
rect 23029 8449 23063 8483
rect 23765 8449 23799 8483
rect 24225 8449 24259 8483
rect 26065 8449 26099 8483
rect 26249 8449 26283 8483
rect 27077 8449 27111 8483
rect 2973 8381 3007 8415
rect 3893 8381 3927 8415
rect 6469 8381 6503 8415
rect 7297 8381 7331 8415
rect 7573 8381 7607 8415
rect 8493 8381 8527 8415
rect 9137 8381 9171 8415
rect 9689 8381 9723 8415
rect 10701 8381 10735 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 13093 8381 13127 8415
rect 15577 8381 15611 8415
rect 16221 8381 16255 8415
rect 17509 8381 17543 8415
rect 18153 8381 18187 8415
rect 18613 8381 18647 8415
rect 20269 8381 20303 8415
rect 21833 8381 21867 8415
rect 23213 8381 23247 8415
rect 24409 8381 24443 8415
rect 24593 8381 24627 8415
rect 25329 8381 25363 8415
rect 27261 8381 27295 8415
rect 27813 8381 27847 8415
rect 27997 8381 28031 8415
rect 1869 8313 1903 8347
rect 8677 8313 8711 8347
rect 9321 8313 9355 8347
rect 15209 8313 15243 8347
rect 16865 8313 16899 8347
rect 20729 8313 20763 8347
rect 23581 8313 23615 8347
rect 24041 8313 24075 8347
rect 2789 8245 2823 8279
rect 5457 8245 5491 8279
rect 6837 8245 6871 8279
rect 12725 8245 12759 8279
rect 14749 8245 14783 8279
rect 15853 8245 15887 8279
rect 17141 8245 17175 8279
rect 19073 8245 19107 8279
rect 25973 8245 26007 8279
rect 26433 8245 26467 8279
rect 27537 8245 27571 8279
rect 2789 8041 2823 8075
rect 4997 8041 5031 8075
rect 12725 8041 12759 8075
rect 14197 8041 14231 8075
rect 15853 8041 15887 8075
rect 19625 8041 19659 8075
rect 21557 8041 21591 8075
rect 23489 8041 23523 8075
rect 24409 8041 24443 8075
rect 24777 8041 24811 8075
rect 28273 8041 28307 8075
rect 7021 7973 7055 8007
rect 17693 7973 17727 8007
rect 27169 7973 27203 8007
rect 27629 7973 27663 8007
rect 4813 7905 4847 7939
rect 5917 7905 5951 7939
rect 6837 7905 6871 7939
rect 8125 7905 8159 7939
rect 8309 7905 8343 7939
rect 11621 7905 11655 7939
rect 12081 7905 12115 7939
rect 12817 7905 12851 7939
rect 13001 7905 13035 7939
rect 13645 7905 13679 7939
rect 15945 7905 15979 7939
rect 16129 7905 16163 7939
rect 16773 7905 16807 7939
rect 18429 7905 18463 7939
rect 19257 7905 19291 7939
rect 22293 7905 22327 7939
rect 24961 7905 24995 7939
rect 26525 7905 26559 7939
rect 1409 7837 1443 7871
rect 3893 7837 3927 7871
rect 4629 7837 4663 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 6561 7837 6595 7871
rect 6653 7837 6687 7871
rect 7481 7837 7515 7871
rect 8769 7837 8803 7871
rect 9137 7837 9171 7871
rect 9788 7837 9822 7871
rect 11437 7837 11471 7871
rect 11529 7837 11563 7871
rect 12265 7837 12299 7871
rect 13553 7837 13587 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 16681 7837 16715 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 18613 7837 18647 7871
rect 19441 7837 19475 7871
rect 20361 7837 20395 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 21925 7837 21959 7871
rect 22109 7837 22143 7871
rect 22845 7837 22879 7871
rect 23397 7837 23431 7871
rect 23673 7837 23707 7871
rect 24133 7837 24167 7871
rect 24593 7837 24627 7871
rect 24685 7837 24719 7871
rect 25228 7837 25262 7871
rect 26709 7837 26743 7871
rect 27261 7837 27295 7871
rect 27445 7837 27479 7871
rect 28089 7837 28123 7871
rect 28549 7837 28583 7871
rect 1676 7769 1710 7803
rect 3249 7769 3283 7803
rect 4537 7769 4571 7803
rect 10048 7769 10082 7803
rect 20545 7769 20579 7803
rect 3525 7701 3559 7735
rect 5365 7701 5399 7735
rect 5641 7701 5675 7735
rect 8033 7701 8067 7735
rect 9689 7701 9723 7735
rect 11161 7701 11195 7735
rect 11253 7701 11287 7735
rect 13461 7701 13495 7735
rect 15117 7701 15151 7735
rect 16589 7701 16623 7735
rect 16957 7701 16991 7735
rect 17509 7701 17543 7735
rect 17969 7701 18003 7735
rect 19073 7701 19107 7735
rect 20177 7701 20211 7735
rect 21005 7701 21039 7735
rect 21741 7701 21775 7735
rect 22753 7701 22787 7735
rect 22937 7701 22971 7735
rect 23213 7701 23247 7735
rect 23949 7701 23983 7735
rect 26341 7701 26375 7735
rect 28365 7701 28399 7735
rect 5089 7497 5123 7531
rect 5825 7497 5859 7531
rect 6377 7497 6411 7531
rect 14105 7497 14139 7531
rect 15301 7497 15335 7531
rect 16865 7497 16899 7531
rect 19533 7497 19567 7531
rect 19717 7497 19751 7531
rect 22477 7497 22511 7531
rect 23213 7497 23247 7531
rect 25513 7497 25547 7531
rect 2145 7429 2179 7463
rect 7012 7429 7046 7463
rect 9873 7429 9907 7463
rect 10793 7429 10827 7463
rect 13737 7429 13771 7463
rect 20361 7429 20395 7463
rect 21097 7429 21131 7463
rect 1593 7361 1627 7395
rect 2513 7361 2547 7395
rect 2789 7361 2823 7395
rect 2881 7361 2915 7395
rect 3617 7361 3651 7395
rect 4629 7361 4663 7395
rect 5181 7361 5215 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 8217 7361 8251 7395
rect 8484 7361 8518 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 14013 7361 14047 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 15577 7361 15611 7395
rect 15669 7361 15703 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 17049 7361 17083 7395
rect 17417 7361 17451 7395
rect 18153 7361 18187 7395
rect 18889 7361 18923 7395
rect 19441 7361 19475 7395
rect 19901 7361 19935 7395
rect 20269 7361 20303 7395
rect 21373 7361 21407 7395
rect 23489 7361 23523 7395
rect 25697 7361 25731 7395
rect 25973 7361 26007 7395
rect 26157 7361 26191 7395
rect 27169 7361 27203 7395
rect 27445 7361 27479 7395
rect 28181 7361 28215 7395
rect 3065 7293 3099 7327
rect 3801 7293 3835 7327
rect 4445 7293 4479 7327
rect 5365 7293 5399 7327
rect 9781 7293 9815 7327
rect 11713 7293 11747 7327
rect 12357 7293 12391 7327
rect 12541 7293 12575 7327
rect 13001 7293 13035 7327
rect 13093 7293 13127 7327
rect 13277 7293 13311 7327
rect 14657 7293 14691 7327
rect 15853 7293 15887 7327
rect 17233 7293 17267 7327
rect 17969 7293 18003 7327
rect 18705 7293 18739 7327
rect 21833 7293 21867 7327
rect 22017 7293 22051 7327
rect 22569 7293 22603 7327
rect 22753 7293 22787 7327
rect 23581 7293 23615 7327
rect 23765 7293 23799 7327
rect 24225 7293 24259 7327
rect 27629 7293 27663 7327
rect 2329 7225 2363 7259
rect 2605 7225 2639 7259
rect 3525 7225 3559 7259
rect 3985 7225 4019 7259
rect 9597 7225 9631 7259
rect 10977 7225 11011 7259
rect 13829 7225 13863 7259
rect 15393 7225 15427 7259
rect 17877 7225 17911 7259
rect 18337 7225 18371 7259
rect 19349 7225 19383 7259
rect 20085 7225 20119 7259
rect 26985 7225 27019 7259
rect 6101 7157 6135 7191
rect 8125 7157 8159 7191
rect 11897 7157 11931 7191
rect 14381 7157 14415 7191
rect 16129 7157 16163 7191
rect 21465 7157 21499 7191
rect 23305 7157 23339 7191
rect 25789 7157 25823 7191
rect 26709 7157 26743 7191
rect 27905 7157 27939 7191
rect 28273 7157 28307 7191
rect 3893 6953 3927 6987
rect 4169 6953 4203 6987
rect 5181 6953 5215 6987
rect 6837 6953 6871 6987
rect 7389 6953 7423 6987
rect 9873 6953 9907 6987
rect 11161 6953 11195 6987
rect 11529 6953 11563 6987
rect 12449 6953 12483 6987
rect 13093 6953 13127 6987
rect 14749 6953 14783 6987
rect 15577 6953 15611 6987
rect 17325 6953 17359 6987
rect 18889 6953 18923 6987
rect 22753 6953 22787 6987
rect 26709 6953 26743 6987
rect 14381 6885 14415 6919
rect 16773 6885 16807 6919
rect 22293 6885 22327 6919
rect 24501 6885 24535 6919
rect 28181 6885 28215 6919
rect 5457 6817 5491 6851
rect 7205 6817 7239 6851
rect 10977 6817 11011 6851
rect 11805 6817 11839 6851
rect 12541 6817 12575 6851
rect 20913 6817 20947 6851
rect 21833 6817 21867 6851
rect 22385 6817 22419 6851
rect 22569 6817 22603 6851
rect 23581 6817 23615 6851
rect 26157 6817 26191 6851
rect 27077 6817 27111 6851
rect 2421 6749 2455 6783
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 5365 6749 5399 6783
rect 7021 6749 7055 6783
rect 8309 6749 8343 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 9781 6749 9815 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 10793 6749 10827 6783
rect 11713 6749 11747 6783
rect 12725 6749 12759 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 16221 6749 16255 6783
rect 16497 6749 16531 6783
rect 16957 6749 16991 6783
rect 17073 6749 17107 6783
rect 17509 6749 17543 6783
rect 17785 6749 17819 6783
rect 18061 6749 18095 6783
rect 18337 6749 18371 6783
rect 18797 6749 18831 6783
rect 19073 6749 19107 6783
rect 19257 6749 19291 6783
rect 19993 6749 20027 6783
rect 21649 6749 21683 6783
rect 23121 6749 23155 6783
rect 24225 6749 24259 6783
rect 24433 6749 24467 6783
rect 24685 6749 24719 6783
rect 25881 6749 25915 6783
rect 27261 6749 27295 6783
rect 27813 6749 27847 6783
rect 27997 6749 28031 6783
rect 5724 6681 5758 6715
rect 13737 6681 13771 6715
rect 16589 6681 16623 6715
rect 20085 6681 20119 6715
rect 20545 6681 20579 6715
rect 20637 6681 20671 6715
rect 23673 6681 23707 6715
rect 25145 6681 25179 6715
rect 25237 6681 25271 6715
rect 25789 6681 25823 6715
rect 2513 6613 2547 6647
rect 3525 6613 3559 6647
rect 4997 6613 5031 6647
rect 8125 6613 8159 6647
rect 9229 6613 9263 6647
rect 9689 6613 9723 6647
rect 10057 6613 10091 6647
rect 10609 6613 10643 6647
rect 14197 6613 14231 6647
rect 15025 6613 15059 6647
rect 15393 6613 15427 6647
rect 16037 6613 16071 6647
rect 16313 6613 16347 6647
rect 17141 6613 17175 6647
rect 17601 6613 17635 6647
rect 18245 6613 18279 6647
rect 18429 6613 18463 6647
rect 18613 6613 18647 6647
rect 19901 6613 19935 6647
rect 23213 6613 23247 6647
rect 24777 6613 24811 6647
rect 25973 6613 26007 6647
rect 27721 6613 27755 6647
rect 5641 6409 5675 6443
rect 6009 6409 6043 6443
rect 7021 6409 7055 6443
rect 8769 6409 8803 6443
rect 11713 6409 11747 6443
rect 12081 6409 12115 6443
rect 12265 6409 12299 6443
rect 12725 6409 12759 6443
rect 13829 6409 13863 6443
rect 15393 6409 15427 6443
rect 20729 6409 20763 6443
rect 21465 6409 21499 6443
rect 26801 6409 26835 6443
rect 28365 6409 28399 6443
rect 22928 6341 22962 6375
rect 24777 6341 24811 6375
rect 2789 6273 2823 6307
rect 3056 6273 3090 6307
rect 4261 6273 4295 6307
rect 4528 6273 4562 6307
rect 5733 6273 5767 6307
rect 6193 6273 6227 6307
rect 6377 6273 6411 6307
rect 7297 6273 7331 6307
rect 7389 6273 7423 6307
rect 7849 6273 7883 6307
rect 8493 6273 8527 6307
rect 8953 6273 8987 6307
rect 9045 6273 9079 6307
rect 9229 6273 9263 6307
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 12449 6273 12483 6307
rect 12909 6273 12943 6307
rect 14013 6273 14047 6307
rect 14565 6273 14599 6307
rect 14933 6273 14967 6307
rect 15301 6273 15335 6307
rect 15577 6273 15611 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 17224 6273 17258 6307
rect 18797 6273 18831 6307
rect 19349 6273 19383 6307
rect 19616 6273 19650 6307
rect 21005 6273 21039 6307
rect 21925 6273 21959 6307
rect 22661 6273 22695 6307
rect 24133 6273 24167 6307
rect 25421 6273 25455 6307
rect 25688 6273 25722 6307
rect 26985 6273 27019 6307
rect 1961 6205 1995 6239
rect 9781 6205 9815 6239
rect 9965 6205 9999 6239
rect 10517 6205 10551 6239
rect 10701 6205 10735 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 15761 6205 15795 6239
rect 18613 6205 18647 6239
rect 20821 6205 20855 6239
rect 22477 6205 22511 6239
rect 24685 6205 24719 6239
rect 27721 6205 27755 6239
rect 27905 6205 27939 6239
rect 7113 6137 7147 6171
rect 10425 6137 10459 6171
rect 10885 6137 10919 6171
rect 15025 6137 15059 6171
rect 16313 6137 16347 6171
rect 25237 6137 25271 6171
rect 2513 6069 2547 6103
rect 4169 6069 4203 6103
rect 5825 6069 5859 6103
rect 7481 6069 7515 6103
rect 7665 6069 7699 6103
rect 8585 6069 8619 6103
rect 9597 6069 9631 6103
rect 16221 6069 16255 6103
rect 16773 6069 16807 6103
rect 18337 6069 18371 6103
rect 19257 6069 19291 6103
rect 24041 6069 24075 6103
rect 24225 6069 24259 6103
rect 27629 6069 27663 6103
rect 3433 5865 3467 5899
rect 4445 5865 4479 5899
rect 7665 5865 7699 5899
rect 8401 5865 8435 5899
rect 9597 5865 9631 5899
rect 10885 5865 10919 5899
rect 11161 5865 11195 5899
rect 12817 5865 12851 5899
rect 13093 5865 13127 5899
rect 13277 5865 13311 5899
rect 16221 5865 16255 5899
rect 19625 5865 19659 5899
rect 20913 5865 20947 5899
rect 23581 5865 23615 5899
rect 25513 5865 25547 5899
rect 26249 5865 26283 5899
rect 27813 5865 27847 5899
rect 14105 5797 14139 5831
rect 16681 5797 16715 5831
rect 18613 5797 18647 5831
rect 19993 5797 20027 5831
rect 23765 5797 23799 5831
rect 25881 5797 25915 5831
rect 2053 5729 2087 5763
rect 3801 5729 3835 5763
rect 5825 5729 5859 5763
rect 8217 5729 8251 5763
rect 9137 5729 9171 5763
rect 10057 5729 10091 5763
rect 11437 5729 11471 5763
rect 13553 5729 13587 5763
rect 14841 5729 14875 5763
rect 15025 5729 15059 5763
rect 15761 5729 15795 5763
rect 16313 5729 16347 5763
rect 18429 5729 18463 5763
rect 19441 5729 19475 5763
rect 20269 5729 20303 5763
rect 21005 5729 21039 5763
rect 21189 5729 21223 5763
rect 23029 5729 23063 5763
rect 23213 5729 23247 5763
rect 26433 5729 26467 5763
rect 27905 5729 27939 5763
rect 1593 5661 1627 5695
rect 1961 5661 1995 5695
rect 2320 5661 2354 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 5641 5661 5675 5695
rect 6561 5661 6595 5695
rect 6745 5661 6779 5695
rect 7297 5661 7331 5695
rect 7481 5661 7515 5695
rect 8033 5661 8067 5695
rect 8953 5661 8987 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 11069 5661 11103 5695
rect 11345 5661 11379 5695
rect 13001 5661 13035 5695
rect 13461 5661 13495 5695
rect 14289 5661 14323 5695
rect 14749 5661 14783 5695
rect 15577 5661 15611 5695
rect 16497 5661 16531 5695
rect 17325 5661 17359 5695
rect 17509 5661 17543 5695
rect 18245 5661 18279 5695
rect 19257 5661 19291 5695
rect 20177 5661 20211 5695
rect 20453 5661 20487 5695
rect 23949 5661 23983 5695
rect 24041 5661 24075 5695
rect 24409 5661 24443 5695
rect 25145 5661 25179 5695
rect 25329 5661 25363 5695
rect 26065 5661 26099 5695
rect 26157 5661 26191 5695
rect 26700 5661 26734 5695
rect 11682 5593 11716 5627
rect 18061 5593 18095 5627
rect 22845 5593 22879 5627
rect 28549 5593 28583 5627
rect 1409 5525 1443 5559
rect 1777 5525 1811 5559
rect 5549 5525 5583 5559
rect 6285 5525 6319 5559
rect 7205 5525 7239 5559
rect 9781 5525 9815 5559
rect 10701 5525 10735 5559
rect 14565 5525 14599 5559
rect 15485 5525 15519 5559
rect 17141 5525 17175 5559
rect 24133 5525 24167 5559
rect 25053 5525 25087 5559
rect 2789 5321 2823 5355
rect 4721 5321 4755 5355
rect 5733 5321 5767 5355
rect 6009 5321 6043 5355
rect 7113 5321 7147 5355
rect 7481 5321 7515 5355
rect 9137 5321 9171 5355
rect 9781 5321 9815 5355
rect 10609 5321 10643 5355
rect 11345 5321 11379 5355
rect 15485 5321 15519 5355
rect 16313 5321 16347 5355
rect 16681 5321 16715 5355
rect 18429 5321 18463 5355
rect 21925 5321 21959 5355
rect 24133 5321 24167 5355
rect 24869 5321 24903 5355
rect 25789 5321 25823 5355
rect 28549 5321 28583 5355
rect 12081 5253 12115 5287
rect 13829 5253 13863 5287
rect 14197 5253 14231 5287
rect 16221 5253 16255 5287
rect 19809 5253 19843 5287
rect 19901 5253 19935 5287
rect 22477 5253 22511 5287
rect 23020 5253 23054 5287
rect 27436 5253 27470 5287
rect 1409 5185 1443 5219
rect 1676 5185 1710 5219
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 3801 5185 3835 5219
rect 4905 5185 4939 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 5925 5185 5959 5219
rect 6193 5185 6227 5219
rect 6469 5185 6503 5219
rect 7413 5185 7447 5219
rect 7849 5185 7883 5219
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 8493 5185 8527 5219
rect 8953 5185 8987 5219
rect 9321 5185 9355 5219
rect 9597 5185 9631 5219
rect 9689 5185 9723 5219
rect 10793 5185 10827 5219
rect 11713 5185 11747 5219
rect 13185 5185 13219 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 15025 5185 15059 5219
rect 15577 5185 15611 5219
rect 16497 5185 16531 5219
rect 16865 5185 16899 5219
rect 17785 5185 17819 5219
rect 18521 5185 18555 5219
rect 18981 5185 19015 5219
rect 21281 5185 21315 5219
rect 21373 5185 21407 5219
rect 21833 5185 21867 5219
rect 22109 5185 22143 5219
rect 22393 5185 22427 5219
rect 22753 5185 22787 5219
rect 24409 5185 24443 5219
rect 25973 5185 26007 5219
rect 26341 5185 26375 5219
rect 27169 5185 27203 5219
rect 3985 5117 4019 5151
rect 6653 5117 6687 5151
rect 9965 5117 9999 5151
rect 10149 5117 10183 5151
rect 12449 5117 12483 5151
rect 12633 5117 12667 5151
rect 14105 5117 14139 5151
rect 14381 5117 14415 5151
rect 14841 5117 14875 5151
rect 15761 5117 15795 5151
rect 17141 5117 17175 5151
rect 17969 5117 18003 5151
rect 19165 5117 19199 5151
rect 20637 5117 20671 5151
rect 24225 5117 24259 5151
rect 25145 5117 25179 5151
rect 25329 5117 25363 5151
rect 4997 5049 5031 5083
rect 7665 5049 7699 5083
rect 8217 5049 8251 5083
rect 9413 5049 9447 5083
rect 13461 5049 13495 5083
rect 18613 5049 18647 5083
rect 20361 5049 20395 5083
rect 22201 5049 22235 5083
rect 3525 4981 3559 5015
rect 4445 4981 4479 5015
rect 5273 4981 5307 5015
rect 7941 4981 7975 5015
rect 8585 4981 8619 5015
rect 8769 4981 8803 5015
rect 12817 4981 12851 5015
rect 13369 4981 13403 5015
rect 17693 4981 17727 5015
rect 19349 4981 19383 5015
rect 21189 4981 21223 5015
rect 2145 4777 2179 4811
rect 3893 4777 3927 4811
rect 7205 4777 7239 4811
rect 8493 4777 8527 4811
rect 13001 4777 13035 4811
rect 19257 4777 19291 4811
rect 22201 4777 22235 4811
rect 25053 4777 25087 4811
rect 25789 4777 25823 4811
rect 26525 4777 26559 4811
rect 28273 4777 28307 4811
rect 6837 4709 6871 4743
rect 9413 4709 9447 4743
rect 9781 4709 9815 4743
rect 11069 4709 11103 4743
rect 13829 4709 13863 4743
rect 21189 4709 21223 4743
rect 23213 4709 23247 4743
rect 23673 4709 23707 4743
rect 24041 4709 24075 4743
rect 2237 4641 2271 4675
rect 4353 4641 4387 4675
rect 5733 4641 5767 4675
rect 6377 4641 6411 4675
rect 7389 4641 7423 4675
rect 8309 4641 8343 4675
rect 9229 4641 9263 4675
rect 10425 4641 10459 4675
rect 10793 4641 10827 4675
rect 11345 4641 11379 4675
rect 13277 4641 13311 4675
rect 14289 4641 14323 4675
rect 15301 4641 15335 4675
rect 16129 4641 16163 4675
rect 17049 4641 17083 4675
rect 17601 4641 17635 4675
rect 22569 4641 22603 4675
rect 26985 4641 27019 4675
rect 27169 4641 27203 4675
rect 27353 4641 27387 4675
rect 27905 4641 27939 4675
rect 28089 4641 28123 4675
rect 1593 4573 1627 4607
rect 3801 4573 3835 4607
rect 4169 4573 4203 4607
rect 4905 4573 4939 4607
rect 5549 4573 5583 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6193 4573 6227 4607
rect 7113 4573 7147 4607
rect 7573 4573 7607 4607
rect 8033 4573 8067 4607
rect 8125 4573 8159 4607
rect 9045 4573 9079 4607
rect 9965 4573 9999 4607
rect 10057 4573 10091 4607
rect 10333 4573 10367 4607
rect 10609 4573 10643 4607
rect 12909 4573 12943 4607
rect 14105 4573 14139 4607
rect 16313 4573 16347 4607
rect 16865 4573 16899 4607
rect 17785 4573 17819 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 21557 4573 21591 4607
rect 22385 4573 22419 4607
rect 22753 4573 22787 4607
rect 23305 4573 23339 4607
rect 23489 4573 23523 4607
rect 24225 4573 24259 4607
rect 24409 4573 24443 4607
rect 24593 4573 24627 4607
rect 25329 4573 25363 4607
rect 25421 4573 25455 4607
rect 25605 4573 25639 4607
rect 26157 4573 26191 4607
rect 26341 4573 26375 4607
rect 26893 4573 26927 4607
rect 2504 4505 2538 4539
rect 11612 4505 11646 4539
rect 13362 4505 13396 4539
rect 18429 4505 18463 4539
rect 18521 4505 18555 4539
rect 19073 4505 19107 4539
rect 20076 4505 20110 4539
rect 27813 4505 27847 4539
rect 3617 4437 3651 4471
rect 4813 4437 4847 4471
rect 4997 4437 5031 4471
rect 5365 4437 5399 4471
rect 6009 4437 6043 4471
rect 10149 4437 10183 4471
rect 12725 4437 12759 4471
rect 16773 4437 16807 4471
rect 17509 4437 17543 4471
rect 18245 4437 18279 4471
rect 19533 4437 19567 4471
rect 22109 4437 22143 4471
rect 25145 4437 25179 4471
rect 4261 4233 4295 4267
rect 5273 4233 5307 4267
rect 5457 4233 5491 4267
rect 7021 4233 7055 4267
rect 11161 4233 11195 4267
rect 13185 4233 13219 4267
rect 16221 4233 16255 4267
rect 17417 4233 17451 4267
rect 24685 4233 24719 4267
rect 24777 4233 24811 4267
rect 27721 4233 27755 4267
rect 13461 4165 13495 4199
rect 17969 4165 18003 4199
rect 1593 4097 1627 4131
rect 2145 4097 2179 4131
rect 2412 4097 2446 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 6193 4097 6227 4131
rect 8125 4101 8159 4135
rect 8401 4097 8435 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 11345 4097 11379 4131
rect 11713 4097 11747 4131
rect 12072 4097 12106 4131
rect 16129 4097 16163 4131
rect 17601 4097 17635 4131
rect 18705 4097 18739 4131
rect 19625 4097 19659 4131
rect 19901 4097 19935 4131
rect 20168 4097 20202 4131
rect 21557 4097 21591 4131
rect 22100 4097 22134 4131
rect 24961 4097 24995 4131
rect 25237 4097 25271 4131
rect 27261 4097 27295 4131
rect 28181 4097 28215 4131
rect 4353 4029 4387 4063
rect 6377 4029 6411 4063
rect 6561 4029 6595 4063
rect 7113 4029 7147 4063
rect 7297 4029 7331 4063
rect 8217 4029 8251 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 10057 4029 10091 4063
rect 10425 4029 10459 4063
rect 11805 4029 11839 4063
rect 13277 4029 13311 4063
rect 13829 4029 13863 4063
rect 15209 4029 15243 4063
rect 16773 4029 16807 4063
rect 17877 4029 17911 4063
rect 19257 4029 19291 4063
rect 21833 4029 21867 4063
rect 23305 4029 23339 4063
rect 24041 4029 24075 4063
rect 24225 4029 24259 4063
rect 25329 4029 25363 4063
rect 26065 4029 26099 4063
rect 26249 4029 26283 4063
rect 27077 4029 27111 4063
rect 28273 4029 28307 4063
rect 3525 3961 3559 3995
rect 4813 3961 4847 3995
rect 6009 3961 6043 3995
rect 7481 3961 7515 3995
rect 7941 3961 7975 3995
rect 15853 3961 15887 3995
rect 18429 3961 18463 3995
rect 21281 3961 21315 3995
rect 23949 3961 23983 3995
rect 25053 3961 25087 3995
rect 26433 3961 26467 3995
rect 27997 3961 28031 3995
rect 1409 3893 1443 3927
rect 5825 3893 5859 3927
rect 8585 3893 8619 3927
rect 9321 3893 9355 3927
rect 9689 3893 9723 3927
rect 10609 3893 10643 3927
rect 11529 3893 11563 3927
rect 17325 3893 17359 3927
rect 19441 3893 19475 3927
rect 21373 3893 21407 3927
rect 23213 3893 23247 3927
rect 25973 3893 26007 3927
rect 1869 3689 1903 3723
rect 3249 3689 3283 3723
rect 4537 3689 4571 3723
rect 5457 3689 5491 3723
rect 8585 3689 8619 3723
rect 9873 3689 9907 3723
rect 12817 3689 12851 3723
rect 14105 3689 14139 3723
rect 16865 3689 16899 3723
rect 24777 3689 24811 3723
rect 26249 3689 26283 3723
rect 26617 3689 26651 3723
rect 26985 3689 27019 3723
rect 2145 3621 2179 3655
rect 5733 3621 5767 3655
rect 6009 3621 6043 3655
rect 6285 3621 6319 3655
rect 11345 3621 11379 3655
rect 11805 3621 11839 3655
rect 13001 3621 13035 3655
rect 15761 3621 15795 3655
rect 22569 3621 22603 3655
rect 2605 3553 2639 3587
rect 3525 3553 3559 3587
rect 6929 3553 6963 3587
rect 7941 3553 7975 3587
rect 8125 3553 8159 3587
rect 9413 3553 9447 3587
rect 19717 3553 19751 3587
rect 21189 3553 21223 3587
rect 23397 3553 23431 3587
rect 25789 3553 25823 3587
rect 25881 3553 25915 3587
rect 26065 3553 26099 3587
rect 27169 3553 27203 3587
rect 1501 3485 1535 3519
rect 1777 3485 1811 3519
rect 2053 3485 2087 3519
rect 2513 3485 2547 3519
rect 3433 3487 3467 3521
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 4721 3485 4755 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 6561 3485 6595 3519
rect 6837 3485 6871 3519
rect 7113 3485 7147 3519
rect 8953 3485 8987 3519
rect 9045 3485 9079 3519
rect 9229 3485 9263 3519
rect 9965 3485 9999 3519
rect 10701 3485 10735 3519
rect 10885 3485 10919 3519
rect 11437 3485 11471 3519
rect 11621 3485 11655 3519
rect 12265 3485 12299 3519
rect 13185 3485 13219 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 14381 3485 14415 3519
rect 16037 3485 16071 3519
rect 16681 3485 16715 3519
rect 17141 3485 17175 3519
rect 17233 3485 17267 3519
rect 19257 3485 19291 3519
rect 22753 3485 22787 3519
rect 24409 3485 24443 3519
rect 24593 3485 24627 3519
rect 25145 3485 25179 3519
rect 26801 3485 26835 3519
rect 26893 3485 26927 3519
rect 1593 3417 1627 3451
rect 5181 3417 5215 3451
rect 6653 3417 6687 3451
rect 13921 3417 13955 3451
rect 14626 3417 14660 3451
rect 17500 3417 17534 3451
rect 19441 3417 19475 3451
rect 21456 3417 21490 3451
rect 24041 3417 24075 3451
rect 27436 3417 27470 3451
rect 2329 3349 2363 3383
rect 7757 3349 7791 3383
rect 10609 3349 10643 3383
rect 16589 3349 16623 3383
rect 16957 3349 16991 3383
rect 18613 3349 18647 3383
rect 18797 3349 18831 3383
rect 23305 3349 23339 3383
rect 28549 3349 28583 3383
rect 4077 3145 4111 3179
rect 4537 3145 4571 3179
rect 6469 3145 6503 3179
rect 9505 3145 9539 3179
rect 11805 3145 11839 3179
rect 14841 3145 14875 3179
rect 16313 3145 16347 3179
rect 17417 3145 17451 3179
rect 17509 3145 17543 3179
rect 21557 3145 21591 3179
rect 23765 3145 23799 3179
rect 26801 3145 26835 3179
rect 5080 3077 5114 3111
rect 12256 3077 12290 3111
rect 19901 3077 19935 3111
rect 1409 3009 1443 3043
rect 1685 3009 1719 3043
rect 1777 3009 1811 3043
rect 2697 3009 2731 3043
rect 2953 3009 2987 3043
rect 4261 3009 4295 3043
rect 4721 3009 4755 3043
rect 4813 3009 4847 3043
rect 6377 3009 6411 3043
rect 6745 3009 6779 3043
rect 8033 3009 8067 3043
rect 8125 3009 8159 3043
rect 8381 3009 8415 3043
rect 9781 3009 9815 3043
rect 10048 3009 10082 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 13461 3009 13495 3043
rect 13728 3009 13762 3043
rect 14933 3009 14967 3043
rect 15200 3009 15234 3043
rect 17693 3009 17727 3043
rect 17969 3009 18003 3043
rect 18061 3009 18095 3043
rect 19993 3009 20027 3043
rect 20260 3009 20294 3043
rect 21465 3009 21499 3043
rect 21925 3009 21959 3043
rect 22192 3009 22226 3043
rect 23581 3009 23615 3043
rect 23673 3009 23707 3043
rect 24216 3009 24250 3043
rect 25421 3009 25455 3043
rect 25688 3009 25722 3043
rect 26985 3009 27019 3043
rect 27252 3009 27286 3043
rect 1501 2941 1535 2975
rect 2053 2941 2087 2975
rect 2605 2941 2639 2975
rect 7389 2941 7423 2975
rect 16773 2941 16807 2975
rect 16957 2941 16991 2975
rect 18245 2941 18279 2975
rect 23949 2941 23983 2975
rect 4353 2873 4387 2907
rect 7297 2873 7331 2907
rect 21373 2873 21407 2907
rect 23305 2873 23339 2907
rect 6193 2805 6227 2839
rect 11161 2805 11195 2839
rect 13369 2805 13403 2839
rect 17785 2805 17819 2839
rect 23397 2805 23431 2839
rect 25329 2805 25363 2839
rect 28365 2805 28399 2839
rect 3617 2601 3651 2635
rect 5365 2601 5399 2635
rect 7021 2601 7055 2635
rect 8585 2601 8619 2635
rect 9137 2601 9171 2635
rect 10701 2601 10735 2635
rect 10977 2601 11011 2635
rect 11161 2601 11195 2635
rect 15025 2601 15059 2635
rect 15209 2601 15243 2635
rect 16497 2601 16531 2635
rect 18153 2601 18187 2635
rect 19257 2601 19291 2635
rect 21281 2601 21315 2635
rect 24501 2601 24535 2635
rect 25513 2601 25547 2635
rect 25973 2601 26007 2635
rect 26801 2601 26835 2635
rect 28549 2601 28583 2635
rect 1961 2533 1995 2567
rect 13093 2533 13127 2567
rect 19073 2533 19107 2567
rect 24777 2533 24811 2567
rect 27629 2533 27663 2567
rect 2237 2465 2271 2499
rect 4077 2465 4111 2499
rect 4721 2465 4755 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 9321 2465 9355 2499
rect 11713 2465 11747 2499
rect 16681 2465 16715 2499
rect 19717 2465 19751 2499
rect 19993 2465 20027 2499
rect 20637 2465 20671 2499
rect 21097 2465 21131 2499
rect 21925 2465 21959 2499
rect 22845 2465 22879 2499
rect 26157 2465 26191 2499
rect 27077 2465 27111 2499
rect 27997 2465 28031 2499
rect 1593 2397 1627 2431
rect 1685 2397 1719 2431
rect 2145 2397 2179 2431
rect 4905 2397 4939 2431
rect 5733 2397 5767 2431
rect 6193 2397 6227 2431
rect 7205 2397 7239 2431
rect 9045 2397 9079 2431
rect 9588 2397 9622 2431
rect 10885 2397 10919 2431
rect 11345 2397 11379 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 14749 2397 14783 2431
rect 14841 2397 14875 2431
rect 15393 2397 15427 2431
rect 15669 2397 15703 2431
rect 15945 2397 15979 2431
rect 16948 2397 16982 2431
rect 18337 2397 18371 2431
rect 18429 2397 18463 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 20821 2397 20855 2431
rect 21465 2397 21499 2431
rect 23029 2397 23063 2431
rect 23305 2397 23339 2431
rect 23765 2397 23799 2431
rect 23857 2397 23891 2431
rect 24409 2397 24443 2431
rect 24961 2397 24995 2431
rect 25145 2397 25179 2431
rect 25421 2397 25455 2431
rect 25881 2397 25915 2431
rect 2504 2329 2538 2363
rect 7472 2329 7506 2363
rect 11980 2329 12014 2363
rect 13829 2329 13863 2363
rect 20085 2329 20119 2363
rect 22017 2329 22051 2363
rect 1409 2261 1443 2295
rect 1777 2261 1811 2295
rect 4629 2261 4663 2295
rect 6009 2261 6043 2295
rect 15485 2261 15519 2295
rect 18061 2261 18095 2295
rect 23121 2261 23155 2295
rect 23489 2261 23523 2295
rect 23581 2261 23615 2295
rect 25237 2261 25271 2295
<< metal1 >>
rect 9674 27820 9680 27872
rect 9732 27860 9738 27872
rect 11974 27860 11980 27872
rect 9732 27832 11980 27860
rect 9732 27820 9738 27832
rect 11974 27820 11980 27832
rect 12032 27820 12038 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 23658 27616 23664 27668
rect 23716 27616 23722 27668
rect 3786 27548 3792 27600
rect 3844 27548 3850 27600
rect 3881 27591 3939 27597
rect 3881 27557 3893 27591
rect 3927 27557 3939 27591
rect 3881 27551 3939 27557
rect 5997 27591 6055 27597
rect 5997 27557 6009 27591
rect 6043 27557 6055 27591
rect 5997 27551 6055 27557
rect 6549 27591 6607 27597
rect 6549 27557 6561 27591
rect 6595 27588 6607 27591
rect 8478 27588 8484 27600
rect 6595 27560 8484 27588
rect 6595 27557 6607 27560
rect 6549 27551 6607 27557
rect 3804 27452 3832 27548
rect 3896 27520 3924 27551
rect 4341 27523 4399 27529
rect 3896 27492 4292 27520
rect 4264 27461 4292 27492
rect 4341 27489 4353 27523
rect 4387 27520 4399 27523
rect 5350 27520 5356 27532
rect 4387 27492 5356 27520
rect 4387 27489 4399 27492
rect 4341 27483 4399 27489
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 6012 27520 6040 27551
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 9401 27591 9459 27597
rect 9401 27557 9413 27591
rect 9447 27588 9459 27591
rect 9674 27588 9680 27600
rect 9447 27560 9680 27588
rect 9447 27557 9459 27560
rect 9401 27551 9459 27557
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 12161 27591 12219 27597
rect 11256 27560 12112 27588
rect 7101 27523 7159 27529
rect 6012 27492 7052 27520
rect 4065 27455 4123 27461
rect 4065 27452 4077 27455
rect 3804 27424 4077 27452
rect 4065 27421 4077 27424
rect 4111 27421 4123 27455
rect 4065 27415 4123 27421
rect 4249 27455 4307 27461
rect 4249 27421 4261 27455
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 4571 27424 4844 27452
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 1486 27344 1492 27396
rect 1544 27344 1550 27396
rect 4816 27328 4844 27424
rect 5074 27412 5080 27464
rect 5132 27452 5138 27464
rect 5629 27455 5687 27461
rect 5629 27452 5641 27455
rect 5132 27424 5641 27452
rect 5132 27412 5138 27424
rect 5629 27421 5641 27424
rect 5675 27421 5687 27455
rect 5629 27415 5687 27421
rect 5905 27455 5963 27461
rect 5905 27421 5917 27455
rect 5951 27452 5963 27455
rect 6181 27455 6239 27461
rect 5951 27424 6040 27452
rect 5951 27421 5963 27424
rect 5905 27415 5963 27421
rect 6012 27328 6040 27424
rect 6181 27421 6193 27455
rect 6227 27421 6239 27455
rect 6181 27415 6239 27421
rect 934 27276 940 27328
rect 992 27316 998 27328
rect 1581 27319 1639 27325
rect 1581 27316 1593 27319
rect 992 27288 1593 27316
rect 992 27276 998 27288
rect 1581 27285 1593 27288
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 4614 27276 4620 27328
rect 4672 27276 4678 27328
rect 4798 27276 4804 27328
rect 4856 27276 4862 27328
rect 4890 27276 4896 27328
rect 4948 27276 4954 27328
rect 5442 27276 5448 27328
rect 5500 27276 5506 27328
rect 5718 27276 5724 27328
rect 5776 27276 5782 27328
rect 5994 27276 6000 27328
rect 6052 27276 6058 27328
rect 6196 27316 6224 27415
rect 6730 27412 6736 27464
rect 6788 27412 6794 27464
rect 7024 27461 7052 27492
rect 7101 27489 7113 27523
rect 7147 27520 7159 27523
rect 8938 27520 8944 27532
rect 7147 27492 8944 27520
rect 7147 27489 7159 27492
rect 7101 27483 7159 27489
rect 8938 27480 8944 27492
rect 8996 27480 9002 27532
rect 9125 27523 9183 27529
rect 9125 27489 9137 27523
rect 9171 27520 9183 27523
rect 11256 27520 11284 27560
rect 9171 27492 11284 27520
rect 9171 27489 9183 27492
rect 9125 27483 9183 27489
rect 11422 27480 11428 27532
rect 11480 27520 11486 27532
rect 12084 27520 12112 27560
rect 12161 27557 12173 27591
rect 12207 27588 12219 27591
rect 14185 27591 14243 27597
rect 12207 27560 13308 27588
rect 12207 27557 12219 27560
rect 12161 27551 12219 27557
rect 12345 27523 12403 27529
rect 12345 27520 12357 27523
rect 11480 27492 11744 27520
rect 12084 27492 12357 27520
rect 11480 27480 11486 27492
rect 7009 27455 7067 27461
rect 7009 27421 7021 27455
rect 7055 27421 7067 27455
rect 7009 27415 7067 27421
rect 7285 27455 7343 27461
rect 7285 27421 7297 27455
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27452 8079 27455
rect 8297 27455 8355 27461
rect 8297 27452 8309 27455
rect 8067 27424 8309 27452
rect 8067 27421 8079 27424
rect 8021 27415 8079 27421
rect 8297 27421 8309 27424
rect 8343 27421 8355 27455
rect 8297 27415 8355 27421
rect 8573 27455 8631 27461
rect 8573 27421 8585 27455
rect 8619 27452 8631 27455
rect 9585 27455 9643 27461
rect 9585 27452 9597 27455
rect 8619 27424 9597 27452
rect 8619 27421 8631 27424
rect 8573 27415 8631 27421
rect 9585 27421 9597 27424
rect 9631 27452 9643 27455
rect 9677 27455 9735 27461
rect 9677 27452 9689 27455
rect 9631 27424 9689 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 9677 27421 9689 27424
rect 9723 27421 9735 27455
rect 9677 27415 9735 27421
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27421 10103 27455
rect 10045 27415 10103 27421
rect 6270 27344 6276 27396
rect 6328 27384 6334 27396
rect 7300 27384 7328 27415
rect 6328 27356 7328 27384
rect 8312 27384 8340 27415
rect 8312 27356 8616 27384
rect 6328 27344 6334 27356
rect 8588 27328 8616 27356
rect 9600 27328 9628 27415
rect 10060 27384 10088 27415
rect 10134 27412 10140 27464
rect 10192 27452 10198 27464
rect 10321 27455 10379 27461
rect 10321 27452 10333 27455
rect 10192 27424 10333 27452
rect 10192 27412 10198 27424
rect 10321 27421 10333 27424
rect 10367 27421 10379 27455
rect 10321 27415 10379 27421
rect 10410 27412 10416 27464
rect 10468 27452 10474 27464
rect 10505 27455 10563 27461
rect 10505 27452 10517 27455
rect 10468 27424 10517 27452
rect 10468 27412 10474 27424
rect 10505 27421 10517 27424
rect 10551 27421 10563 27455
rect 10505 27415 10563 27421
rect 11146 27412 11152 27464
rect 11204 27452 11210 27464
rect 11716 27461 11744 27492
rect 12345 27489 12357 27492
rect 12391 27489 12403 27523
rect 13280 27520 13308 27560
rect 14185 27557 14197 27591
rect 14231 27588 14243 27591
rect 15378 27588 15384 27600
rect 14231 27560 15384 27588
rect 14231 27557 14243 27560
rect 14185 27551 14243 27557
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 15746 27548 15752 27600
rect 15804 27548 15810 27600
rect 19150 27548 19156 27600
rect 19208 27588 19214 27600
rect 19797 27591 19855 27597
rect 19797 27588 19809 27591
rect 19208 27560 19809 27588
rect 19208 27548 19214 27560
rect 19797 27557 19809 27560
rect 19843 27557 19855 27591
rect 19797 27551 19855 27557
rect 21358 27548 21364 27600
rect 21416 27588 21422 27600
rect 21416 27560 24348 27588
rect 21416 27548 21422 27560
rect 15764 27520 15792 27548
rect 12345 27483 12403 27489
rect 12452 27492 13216 27520
rect 13280 27492 15792 27520
rect 11241 27455 11299 27461
rect 11241 27452 11253 27455
rect 11204 27424 11253 27452
rect 11204 27412 11210 27424
rect 11241 27421 11253 27424
rect 11287 27421 11299 27455
rect 11241 27415 11299 27421
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 11974 27412 11980 27464
rect 12032 27412 12038 27464
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27454 12127 27455
rect 12115 27426 12204 27454
rect 12115 27421 12127 27426
rect 12069 27415 12127 27421
rect 12176 27384 12204 27426
rect 12452 27384 12480 27492
rect 13188 27461 13216 27492
rect 16850 27480 16856 27532
rect 16908 27520 16914 27532
rect 16908 27492 17816 27520
rect 16908 27480 16914 27492
rect 12529 27455 12587 27461
rect 12529 27421 12541 27455
rect 12575 27421 12587 27455
rect 12529 27415 12587 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27452 13231 27455
rect 13906 27452 13912 27464
rect 13219 27424 13912 27452
rect 13219 27421 13231 27424
rect 13173 27415 13231 27421
rect 10060 27356 11192 27384
rect 12176 27356 12480 27384
rect 6638 27316 6644 27328
rect 6196 27288 6644 27316
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 6822 27276 6828 27328
rect 6880 27276 6886 27328
rect 6914 27276 6920 27328
rect 6972 27316 6978 27328
rect 7745 27319 7803 27325
rect 7745 27316 7757 27319
rect 6972 27288 7757 27316
rect 6972 27276 6978 27288
rect 7745 27285 7757 27288
rect 7791 27285 7803 27319
rect 7745 27279 7803 27285
rect 8113 27319 8171 27325
rect 8113 27285 8125 27319
rect 8159 27316 8171 27319
rect 8294 27316 8300 27328
rect 8159 27288 8300 27316
rect 8159 27285 8171 27288
rect 8113 27279 8171 27285
rect 8294 27276 8300 27288
rect 8352 27276 8358 27328
rect 8386 27276 8392 27328
rect 8444 27276 8450 27328
rect 8570 27276 8576 27328
rect 8628 27276 8634 27328
rect 8665 27319 8723 27325
rect 8665 27285 8677 27319
rect 8711 27316 8723 27319
rect 9030 27316 9036 27328
rect 8711 27288 9036 27316
rect 8711 27285 8723 27288
rect 8665 27279 8723 27285
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 9582 27276 9588 27328
rect 9640 27276 9646 27328
rect 9766 27276 9772 27328
rect 9824 27276 9830 27328
rect 10137 27319 10195 27325
rect 10137 27285 10149 27319
rect 10183 27316 10195 27319
rect 10502 27316 10508 27328
rect 10183 27288 10508 27316
rect 10183 27285 10195 27288
rect 10137 27279 10195 27285
rect 10502 27276 10508 27288
rect 10560 27276 10566 27328
rect 10962 27276 10968 27328
rect 11020 27276 11026 27328
rect 11054 27276 11060 27328
rect 11112 27276 11118 27328
rect 11164 27316 11192 27356
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 11164 27288 11529 27316
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 11517 27279 11575 27285
rect 11793 27319 11851 27325
rect 11793 27285 11805 27319
rect 11839 27316 11851 27319
rect 12544 27316 12572 27415
rect 13906 27412 13912 27424
rect 13964 27412 13970 27464
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27452 14519 27455
rect 14642 27452 14648 27464
rect 14507 27424 14648 27452
rect 14507 27421 14519 27424
rect 14461 27415 14519 27421
rect 12894 27344 12900 27396
rect 12952 27384 12958 27396
rect 14384 27384 14412 27415
rect 14642 27412 14648 27424
rect 14700 27452 14706 27464
rect 14737 27455 14795 27461
rect 14737 27452 14749 27455
rect 14700 27424 14749 27452
rect 14700 27412 14706 27424
rect 14737 27421 14749 27424
rect 14783 27421 14795 27455
rect 14737 27415 14795 27421
rect 15749 27455 15807 27461
rect 15749 27421 15761 27455
rect 15795 27452 15807 27455
rect 15838 27452 15844 27464
rect 15795 27424 15844 27452
rect 15795 27421 15807 27424
rect 15749 27415 15807 27421
rect 15838 27412 15844 27424
rect 15896 27452 15902 27464
rect 17788 27461 17816 27492
rect 18690 27480 18696 27532
rect 18748 27520 18754 27532
rect 20901 27523 20959 27529
rect 18748 27492 20024 27520
rect 18748 27480 18754 27492
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 15896 27424 17509 27452
rect 15896 27412 15902 27424
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 18322 27412 18328 27464
rect 18380 27452 18386 27464
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 18380 27424 19257 27452
rect 18380 27412 18386 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 19518 27412 19524 27464
rect 19576 27461 19582 27464
rect 19996 27461 20024 27492
rect 20901 27489 20913 27523
rect 20947 27520 20959 27523
rect 24320 27520 24348 27560
rect 26234 27548 26240 27600
rect 26292 27588 26298 27600
rect 26513 27591 26571 27597
rect 26513 27588 26525 27591
rect 26292 27560 26525 27588
rect 26292 27548 26298 27560
rect 26513 27557 26525 27560
rect 26559 27557 26571 27591
rect 26513 27551 26571 27557
rect 26602 27548 26608 27600
rect 26660 27548 26666 27600
rect 26620 27520 26648 27548
rect 20947 27492 24256 27520
rect 24320 27492 26648 27520
rect 20947 27489 20959 27492
rect 20901 27483 20959 27489
rect 19576 27455 19603 27461
rect 19591 27452 19603 27455
rect 19981 27455 20039 27461
rect 19591 27424 19748 27452
rect 19591 27421 19603 27424
rect 19576 27415 19603 27421
rect 19576 27412 19582 27415
rect 12952 27356 14412 27384
rect 12952 27344 12958 27356
rect 16482 27344 16488 27396
rect 16540 27384 16546 27396
rect 17589 27387 17647 27393
rect 17589 27384 17601 27387
rect 16540 27356 17601 27384
rect 16540 27344 16546 27356
rect 17589 27353 17601 27356
rect 17635 27353 17647 27387
rect 19720 27384 19748 27424
rect 19981 27421 19993 27455
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 20180 27384 20208 27415
rect 21082 27412 21088 27464
rect 21140 27412 21146 27464
rect 22370 27412 22376 27464
rect 22428 27412 22434 27464
rect 22830 27412 22836 27464
rect 22888 27452 22894 27464
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 22888 27424 23397 27452
rect 22888 27412 22894 27424
rect 23385 27421 23397 27424
rect 23431 27452 23443 27455
rect 23845 27455 23903 27461
rect 23845 27452 23857 27455
rect 23431 27424 23857 27452
rect 23431 27421 23443 27424
rect 23385 27415 23443 27421
rect 23845 27421 23857 27424
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27452 23995 27455
rect 24118 27452 24124 27464
rect 23983 27424 24124 27452
rect 23983 27421 23995 27424
rect 23937 27415 23995 27421
rect 24118 27412 24124 27424
rect 24176 27412 24182 27464
rect 24228 27452 24256 27492
rect 25038 27452 25044 27464
rect 24228 27424 25044 27452
rect 25038 27412 25044 27424
rect 25096 27412 25102 27464
rect 26050 27412 26056 27464
rect 26108 27412 26114 27464
rect 28166 27412 28172 27464
rect 28224 27452 28230 27464
rect 28261 27455 28319 27461
rect 28261 27452 28273 27455
rect 28224 27424 28273 27452
rect 28224 27412 28230 27424
rect 28261 27421 28273 27424
rect 28307 27421 28319 27455
rect 28261 27415 28319 27421
rect 19720 27356 20208 27384
rect 23477 27387 23535 27393
rect 17589 27347 17647 27353
rect 23477 27353 23489 27387
rect 23523 27384 23535 27387
rect 24026 27384 24032 27396
rect 23523 27356 24032 27384
rect 23523 27353 23535 27356
rect 23477 27347 23535 27353
rect 24026 27344 24032 27356
rect 24084 27344 24090 27396
rect 26329 27387 26387 27393
rect 26329 27353 26341 27387
rect 26375 27384 26387 27387
rect 27798 27384 27804 27396
rect 26375 27356 27804 27384
rect 26375 27353 26387 27356
rect 26329 27347 26387 27353
rect 27798 27344 27804 27356
rect 27856 27344 27862 27396
rect 11839 27288 12572 27316
rect 11839 27285 11851 27288
rect 11793 27279 11851 27285
rect 12986 27276 12992 27328
rect 13044 27276 13050 27328
rect 13722 27276 13728 27328
rect 13780 27276 13786 27328
rect 14553 27319 14611 27325
rect 14553 27285 14565 27319
rect 14599 27316 14611 27319
rect 14734 27316 14740 27328
rect 14599 27288 14740 27316
rect 14599 27285 14611 27288
rect 14553 27279 14611 27285
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 15194 27276 15200 27328
rect 15252 27316 15258 27328
rect 15381 27319 15439 27325
rect 15381 27316 15393 27319
rect 15252 27288 15393 27316
rect 15252 27276 15258 27288
rect 15381 27285 15393 27288
rect 15427 27285 15439 27319
rect 15381 27279 15439 27285
rect 16298 27276 16304 27328
rect 16356 27276 16362 27328
rect 17402 27276 17408 27328
rect 17460 27276 17466 27328
rect 17678 27276 17684 27328
rect 17736 27316 17742 27328
rect 17865 27319 17923 27325
rect 17865 27316 17877 27319
rect 17736 27288 17877 27316
rect 17736 27276 17742 27288
rect 17865 27285 17877 27288
rect 17911 27285 17923 27319
rect 17865 27279 17923 27285
rect 18874 27276 18880 27328
rect 18932 27276 18938 27328
rect 19334 27276 19340 27328
rect 19392 27276 19398 27328
rect 19610 27276 19616 27328
rect 19668 27276 19674 27328
rect 20806 27276 20812 27328
rect 20864 27276 20870 27328
rect 21266 27276 21272 27328
rect 21324 27316 21330 27328
rect 21545 27319 21603 27325
rect 21545 27316 21557 27319
rect 21324 27288 21557 27316
rect 21324 27276 21330 27288
rect 21545 27285 21557 27288
rect 21591 27285 21603 27319
rect 21545 27279 21603 27285
rect 22189 27319 22247 27325
rect 22189 27285 22201 27319
rect 22235 27316 22247 27319
rect 22738 27316 22744 27328
rect 22235 27288 22744 27316
rect 22235 27285 22247 27288
rect 22189 27279 22247 27285
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 25869 27319 25927 27325
rect 25869 27285 25881 27319
rect 25915 27316 25927 27319
rect 26510 27316 26516 27328
rect 25915 27288 26516 27316
rect 25915 27285 25927 27288
rect 25869 27279 25927 27285
rect 26510 27276 26516 27288
rect 26568 27276 26574 27328
rect 28442 27276 28448 27328
rect 28500 27276 28506 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1486 27072 1492 27124
rect 1544 27112 1550 27124
rect 1673 27115 1731 27121
rect 1673 27112 1685 27115
rect 1544 27084 1685 27112
rect 1544 27072 1550 27084
rect 1673 27081 1685 27084
rect 1719 27081 1731 27115
rect 4614 27112 4620 27124
rect 1673 27075 1731 27081
rect 4264 27084 4620 27112
rect 2590 27004 2596 27056
rect 2648 27004 2654 27056
rect 2682 27004 2688 27056
rect 2740 27004 2746 27056
rect 4264 27053 4292 27084
rect 4614 27072 4620 27084
rect 4672 27072 4678 27124
rect 4890 27072 4896 27124
rect 4948 27072 4954 27124
rect 5442 27072 5448 27124
rect 5500 27072 5506 27124
rect 5718 27072 5724 27124
rect 5776 27072 5782 27124
rect 6730 27072 6736 27124
rect 6788 27112 6794 27124
rect 8021 27115 8079 27121
rect 8021 27112 8033 27115
rect 6788 27084 8033 27112
rect 6788 27072 6794 27084
rect 8021 27081 8033 27084
rect 8067 27081 8079 27115
rect 8021 27075 8079 27081
rect 8294 27072 8300 27124
rect 8352 27072 8358 27124
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 10597 27115 10655 27121
rect 8444 27084 10180 27112
rect 8444 27072 8450 27084
rect 4249 27047 4307 27053
rect 4249 27013 4261 27047
rect 4295 27013 4307 27047
rect 4249 27007 4307 27013
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26976 1639 26979
rect 2314 26976 2320 26988
rect 1627 26948 2320 26976
rect 1627 26945 1639 26948
rect 1581 26939 1639 26945
rect 2314 26936 2320 26948
rect 2372 26936 2378 26988
rect 2409 26979 2467 26985
rect 2409 26945 2421 26979
rect 2455 26945 2467 26979
rect 2409 26939 2467 26945
rect 3329 26979 3387 26985
rect 3329 26945 3341 26979
rect 3375 26976 3387 26979
rect 3786 26976 3792 26988
rect 3375 26948 3792 26976
rect 3375 26945 3387 26948
rect 3329 26939 3387 26945
rect 2222 26732 2228 26784
rect 2280 26732 2286 26784
rect 2424 26772 2452 26939
rect 3786 26936 3792 26948
rect 3844 26936 3850 26988
rect 4908 26985 4936 27072
rect 4893 26979 4951 26985
rect 4893 26945 4905 26979
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 5077 26979 5135 26985
rect 5077 26945 5089 26979
rect 5123 26976 5135 26979
rect 5460 26976 5488 27072
rect 5123 26948 5488 26976
rect 5736 26976 5764 27072
rect 6638 27004 6644 27056
rect 6696 27044 6702 27056
rect 7006 27044 7012 27056
rect 6696 27016 7012 27044
rect 6696 27004 6702 27016
rect 7006 27004 7012 27016
rect 7064 27044 7070 27056
rect 8312 27044 8340 27072
rect 7064 27016 8248 27044
rect 8312 27016 8984 27044
rect 7064 27004 7070 27016
rect 8220 26988 8248 27016
rect 5905 26979 5963 26985
rect 5905 26976 5917 26979
rect 5736 26948 5917 26976
rect 5123 26945 5135 26948
rect 5077 26939 5135 26945
rect 5905 26945 5917 26948
rect 5951 26945 5963 26979
rect 5905 26939 5963 26945
rect 5994 26936 6000 26988
rect 6052 26936 6058 26988
rect 6089 26979 6147 26985
rect 6089 26945 6101 26979
rect 6135 26976 6147 26979
rect 7469 26979 7527 26985
rect 7469 26976 7481 26979
rect 6135 26948 7481 26976
rect 6135 26945 6147 26948
rect 6089 26939 6147 26945
rect 7469 26945 7481 26948
rect 7515 26945 7527 26979
rect 7469 26939 7527 26945
rect 8202 26936 8208 26988
rect 8260 26936 8266 26988
rect 8956 26985 8984 27016
rect 9030 27004 9036 27056
rect 9088 27044 9094 27056
rect 9088 27016 9996 27044
rect 9088 27004 9094 27016
rect 8297 26979 8355 26985
rect 8297 26945 8309 26979
rect 8343 26945 8355 26979
rect 8297 26939 8355 26945
rect 8941 26979 8999 26985
rect 8941 26945 8953 26979
rect 8987 26945 8999 26979
rect 8941 26939 8999 26945
rect 3510 26868 3516 26920
rect 3568 26868 3574 26920
rect 4157 26911 4215 26917
rect 4157 26908 4169 26911
rect 3712 26880 4169 26908
rect 3712 26849 3740 26880
rect 4157 26877 4169 26880
rect 4203 26877 4215 26911
rect 6270 26908 6276 26920
rect 4157 26871 4215 26877
rect 5736 26880 6276 26908
rect 3145 26843 3203 26849
rect 3145 26809 3157 26843
rect 3191 26840 3203 26843
rect 3697 26843 3755 26849
rect 3697 26840 3709 26843
rect 3191 26812 3709 26840
rect 3191 26809 3203 26812
rect 3145 26803 3203 26809
rect 3697 26809 3709 26812
rect 3743 26809 3755 26843
rect 3697 26803 3755 26809
rect 4709 26843 4767 26849
rect 4709 26809 4721 26843
rect 4755 26840 4767 26843
rect 5258 26840 5264 26852
rect 4755 26812 5264 26840
rect 4755 26809 4767 26812
rect 4709 26803 4767 26809
rect 5258 26800 5264 26812
rect 5316 26800 5322 26852
rect 5736 26849 5764 26880
rect 6270 26868 6276 26880
rect 6328 26868 6334 26920
rect 6362 26868 6368 26920
rect 6420 26868 6426 26920
rect 6549 26911 6607 26917
rect 6549 26877 6561 26911
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 7285 26911 7343 26917
rect 7285 26877 7297 26911
rect 7331 26908 7343 26911
rect 8312 26908 8340 26939
rect 9858 26936 9864 26988
rect 9916 26936 9922 26988
rect 9968 26976 9996 27016
rect 10152 26985 10180 27084
rect 10597 27081 10609 27115
rect 10643 27112 10655 27115
rect 10962 27112 10968 27124
rect 10643 27084 10968 27112
rect 10643 27081 10655 27084
rect 10597 27075 10655 27081
rect 10704 26985 10732 27084
rect 10962 27072 10968 27084
rect 11020 27072 11026 27124
rect 11054 27072 11060 27124
rect 11112 27072 11118 27124
rect 11517 27115 11575 27121
rect 11517 27081 11529 27115
rect 11563 27081 11575 27115
rect 11517 27075 11575 27081
rect 10137 26979 10195 26985
rect 9968 26948 10088 26976
rect 7331 26880 8156 26908
rect 7331 26877 7343 26880
rect 7285 26871 7343 26877
rect 5721 26843 5779 26849
rect 5721 26809 5733 26843
rect 5767 26809 5779 26843
rect 5721 26803 5779 26809
rect 5902 26800 5908 26852
rect 5960 26840 5966 26852
rect 6564 26840 6592 26871
rect 7653 26843 7711 26849
rect 7653 26840 7665 26843
rect 5960 26812 6592 26840
rect 6932 26812 7665 26840
rect 5960 26800 5966 26812
rect 6932 26784 6960 26812
rect 7653 26809 7665 26812
rect 7699 26809 7711 26843
rect 7653 26803 7711 26809
rect 3234 26772 3240 26784
rect 2424 26744 3240 26772
rect 3234 26732 3240 26744
rect 3292 26732 3298 26784
rect 6178 26732 6184 26784
rect 6236 26772 6242 26784
rect 6733 26775 6791 26781
rect 6733 26772 6745 26775
rect 6236 26744 6745 26772
rect 6236 26732 6242 26744
rect 6733 26741 6745 26744
rect 6779 26741 6791 26775
rect 6733 26735 6791 26741
rect 6914 26732 6920 26784
rect 6972 26732 6978 26784
rect 8128 26772 8156 26880
rect 8220 26880 8340 26908
rect 8757 26911 8815 26917
rect 8220 26852 8248 26880
rect 8757 26877 8769 26911
rect 8803 26908 8815 26911
rect 9953 26911 10011 26917
rect 8803 26880 9674 26908
rect 8803 26877 8815 26880
rect 8757 26871 8815 26877
rect 8202 26800 8208 26852
rect 8260 26800 8266 26852
rect 8772 26840 8800 26871
rect 8312 26812 8800 26840
rect 9646 26840 9674 26880
rect 9953 26877 9965 26911
rect 9999 26877 10011 26911
rect 10060 26908 10088 26948
rect 10137 26945 10149 26979
rect 10183 26945 10195 26979
rect 10137 26939 10195 26945
rect 10689 26979 10747 26985
rect 10689 26945 10701 26979
rect 10735 26945 10747 26979
rect 11072 26976 11100 27072
rect 11532 27044 11560 27075
rect 12894 27072 12900 27124
rect 12952 27072 12958 27124
rect 12986 27072 12992 27124
rect 13044 27072 13050 27124
rect 13722 27072 13728 27124
rect 13780 27072 13786 27124
rect 14642 27072 14648 27124
rect 14700 27072 14706 27124
rect 16485 27115 16543 27121
rect 16485 27081 16497 27115
rect 16531 27112 16543 27115
rect 16850 27112 16856 27124
rect 16531 27084 16856 27112
rect 16531 27081 16543 27084
rect 16485 27075 16543 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 18049 27115 18107 27121
rect 18049 27081 18061 27115
rect 18095 27112 18107 27115
rect 18322 27112 18328 27124
rect 18095 27084 18328 27112
rect 18095 27081 18107 27084
rect 18049 27075 18107 27081
rect 18322 27072 18328 27084
rect 18380 27072 18386 27124
rect 18874 27072 18880 27124
rect 18932 27072 18938 27124
rect 19518 27072 19524 27124
rect 19576 27072 19582 27124
rect 20993 27115 21051 27121
rect 20993 27112 21005 27115
rect 19628 27084 21005 27112
rect 11977 27047 12035 27053
rect 11977 27044 11989 27047
rect 11532 27016 11989 27044
rect 11977 27013 11989 27016
rect 12023 27013 12035 27047
rect 13004 27044 13032 27072
rect 11977 27007 12035 27013
rect 12728 27016 13032 27044
rect 13532 27047 13590 27053
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11072 26948 11713 26976
rect 10689 26939 10747 26945
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 10873 26911 10931 26917
rect 10873 26908 10885 26911
rect 10060 26880 10885 26908
rect 9953 26871 10011 26877
rect 10873 26877 10885 26880
rect 10919 26877 10931 26911
rect 10873 26871 10931 26877
rect 11333 26911 11391 26917
rect 11333 26877 11345 26911
rect 11379 26908 11391 26911
rect 11885 26911 11943 26917
rect 11885 26908 11897 26911
rect 11379 26880 11897 26908
rect 11379 26877 11391 26880
rect 11333 26871 11391 26877
rect 11885 26877 11897 26880
rect 11931 26908 11943 26911
rect 12728 26908 12756 27016
rect 13532 27013 13544 27047
rect 13578 27044 13590 27047
rect 13740 27044 13768 27072
rect 18408 27047 18466 27053
rect 13578 27016 13768 27044
rect 15120 27016 18184 27044
rect 13578 27013 13590 27016
rect 13532 27007 13590 27013
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 13081 26979 13139 26985
rect 13081 26976 13093 26979
rect 12860 26948 13093 26976
rect 12860 26936 12866 26948
rect 13081 26945 13093 26948
rect 13127 26945 13139 26979
rect 14274 26976 14280 26988
rect 13081 26939 13139 26945
rect 13188 26948 14280 26976
rect 11931 26880 12756 26908
rect 11931 26877 11943 26880
rect 11885 26871 11943 26877
rect 9858 26840 9864 26852
rect 9646 26812 9864 26840
rect 8312 26772 8340 26812
rect 9858 26800 9864 26812
rect 9916 26800 9922 26852
rect 9968 26840 9996 26871
rect 10042 26840 10048 26852
rect 9968 26812 10048 26840
rect 10042 26800 10048 26812
rect 10100 26840 10106 26852
rect 10778 26840 10784 26852
rect 10100 26812 10784 26840
rect 10100 26800 10106 26812
rect 10778 26800 10784 26812
rect 10836 26800 10842 26852
rect 12434 26800 12440 26852
rect 12492 26800 12498 26852
rect 12621 26843 12679 26849
rect 12621 26809 12633 26843
rect 12667 26840 12679 26843
rect 13188 26840 13216 26948
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 15120 26985 15148 27016
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15372 26979 15430 26985
rect 15372 26945 15384 26979
rect 15418 26976 15430 26979
rect 16298 26976 16304 26988
rect 15418 26948 16304 26976
rect 15418 26945 15430 26948
rect 15372 26939 15430 26945
rect 13262 26868 13268 26920
rect 13320 26868 13326 26920
rect 14752 26908 14780 26939
rect 16298 26936 16304 26948
rect 16356 26936 16362 26988
rect 16592 26908 16620 27016
rect 16936 26979 16994 26985
rect 16936 26945 16948 26979
rect 16982 26976 16994 26979
rect 17402 26976 17408 26988
rect 16982 26948 17408 26976
rect 16982 26945 16994 26948
rect 16936 26939 16994 26945
rect 17402 26936 17408 26948
rect 17460 26936 17466 26988
rect 18156 26985 18184 27016
rect 18408 27013 18420 27047
rect 18454 27044 18466 27047
rect 18892 27044 18920 27072
rect 19628 27044 19656 27084
rect 20993 27081 21005 27084
rect 21039 27081 21051 27115
rect 20993 27075 21051 27081
rect 21269 27115 21327 27121
rect 21269 27081 21281 27115
rect 21315 27112 21327 27115
rect 21358 27112 21364 27124
rect 21315 27084 21364 27112
rect 21315 27081 21327 27084
rect 21269 27075 21327 27081
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 21821 27115 21879 27121
rect 21821 27081 21833 27115
rect 21867 27112 21879 27115
rect 22370 27112 22376 27124
rect 21867 27084 22376 27112
rect 21867 27081 21879 27084
rect 21821 27075 21879 27081
rect 22370 27072 22376 27084
rect 22428 27072 22434 27124
rect 22738 27072 22744 27124
rect 22796 27072 22802 27124
rect 25409 27115 25467 27121
rect 25409 27081 25421 27115
rect 25455 27112 25467 27115
rect 26050 27112 26056 27124
rect 25455 27084 26056 27112
rect 25455 27081 25467 27084
rect 25409 27075 25467 27081
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 18454 27016 18920 27044
rect 18984 27016 19656 27044
rect 19880 27047 19938 27053
rect 18454 27013 18466 27016
rect 18408 27007 18466 27013
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18984 26976 19012 27016
rect 19880 27013 19892 27047
rect 19926 27044 19938 27047
rect 20806 27044 20812 27056
rect 19926 27016 20812 27044
rect 19926 27013 19938 27016
rect 19880 27007 19938 27013
rect 20806 27004 20812 27016
rect 20864 27004 20870 27056
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 18141 26939 18199 26945
rect 18248 26948 19012 26976
rect 19260 26948 21097 26976
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 14752 26880 15148 26908
rect 15120 26852 15148 26880
rect 16592 26880 16681 26908
rect 12667 26812 13216 26840
rect 12667 26809 12679 26812
rect 12621 26803 12679 26809
rect 15102 26800 15108 26852
rect 15160 26800 15166 26852
rect 16592 26784 16620 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 17770 26868 17776 26920
rect 17828 26908 17834 26920
rect 18248 26908 18276 26948
rect 17828 26880 18276 26908
rect 17828 26868 17834 26880
rect 19260 26784 19288 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26877 19671 26911
rect 21100 26908 21128 26939
rect 21450 26936 21456 26988
rect 21508 26976 21514 26988
rect 21981 26979 22039 26985
rect 21981 26976 21993 26979
rect 21508 26948 21993 26976
rect 21508 26936 21514 26948
rect 21981 26945 21993 26948
rect 22027 26976 22039 26979
rect 22089 26979 22147 26985
rect 22089 26976 22101 26979
rect 22027 26948 22101 26976
rect 22027 26945 22039 26948
rect 21981 26939 22039 26945
rect 22089 26945 22101 26948
rect 22135 26945 22147 26979
rect 22089 26939 22147 26945
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26976 22247 26979
rect 22649 26979 22707 26985
rect 22649 26976 22661 26979
rect 22235 26948 22661 26976
rect 22235 26945 22247 26948
rect 22189 26939 22247 26945
rect 22649 26945 22661 26948
rect 22695 26945 22707 26979
rect 22756 26976 22784 27072
rect 27246 27044 27252 27056
rect 23492 27016 27252 27044
rect 23385 26979 23443 26985
rect 23385 26976 23397 26979
rect 22756 26948 23397 26976
rect 22649 26939 22707 26945
rect 23385 26945 23397 26948
rect 23431 26945 23443 26979
rect 23385 26939 23443 26945
rect 22465 26911 22523 26917
rect 21100 26880 21680 26908
rect 19613 26871 19671 26877
rect 8128 26744 8340 26772
rect 8386 26732 8392 26784
rect 8444 26732 8450 26784
rect 9398 26732 9404 26784
rect 9456 26732 9462 26784
rect 9674 26732 9680 26784
rect 9732 26732 9738 26784
rect 10134 26732 10140 26784
rect 10192 26772 10198 26784
rect 13170 26772 13176 26784
rect 10192 26744 13176 26772
rect 10192 26732 10198 26744
rect 13170 26732 13176 26744
rect 13228 26732 13234 26784
rect 14829 26775 14887 26781
rect 14829 26741 14841 26775
rect 14875 26772 14887 26775
rect 15286 26772 15292 26784
rect 14875 26744 15292 26772
rect 14875 26741 14887 26744
rect 14829 26735 14887 26741
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 16574 26732 16580 26784
rect 16632 26732 16638 26784
rect 19242 26732 19248 26784
rect 19300 26732 19306 26784
rect 19628 26772 19656 26871
rect 20622 26772 20628 26784
rect 19628 26744 20628 26772
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 21542 26732 21548 26784
rect 21600 26732 21606 26784
rect 21652 26772 21680 26880
rect 22465 26877 22477 26911
rect 22511 26908 22523 26911
rect 22738 26908 22744 26920
rect 22511 26880 22744 26908
rect 22511 26877 22523 26880
rect 22465 26871 22523 26877
rect 22738 26868 22744 26880
rect 22796 26868 22802 26920
rect 23201 26911 23259 26917
rect 23201 26877 23213 26911
rect 23247 26908 23259 26911
rect 23492 26908 23520 27016
rect 27246 27004 27252 27016
rect 27304 27004 27310 27056
rect 24210 26936 24216 26988
rect 24268 26976 24274 26988
rect 24673 26979 24731 26985
rect 24673 26976 24685 26979
rect 24268 26948 24685 26976
rect 24268 26936 24274 26948
rect 24673 26945 24685 26948
rect 24719 26945 24731 26979
rect 24673 26939 24731 26945
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26976 25651 26979
rect 25774 26976 25780 26988
rect 25639 26948 25780 26976
rect 25639 26945 25651 26948
rect 25593 26939 25651 26945
rect 25774 26936 25780 26948
rect 25832 26976 25838 26988
rect 25869 26979 25927 26985
rect 25869 26976 25881 26979
rect 25832 26948 25881 26976
rect 25832 26936 25838 26948
rect 25869 26945 25881 26948
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26976 26019 26979
rect 26329 26979 26387 26985
rect 26329 26976 26341 26979
rect 26007 26948 26341 26976
rect 26007 26945 26019 26948
rect 25961 26939 26019 26945
rect 26329 26945 26341 26948
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 26510 26936 26516 26988
rect 26568 26976 26574 26988
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26568 26948 27169 26976
rect 26568 26936 26574 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27890 26936 27896 26988
rect 27948 26936 27954 26988
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 28537 26979 28595 26985
rect 28537 26976 28549 26979
rect 28316 26948 28549 26976
rect 28316 26936 28322 26948
rect 28537 26945 28549 26948
rect 28583 26945 28595 26979
rect 28537 26939 28595 26945
rect 23937 26911 23995 26917
rect 23937 26908 23949 26911
rect 23247 26880 23520 26908
rect 23584 26880 23949 26908
rect 23247 26877 23259 26880
rect 23201 26871 23259 26877
rect 23584 26849 23612 26880
rect 23937 26877 23949 26880
rect 23983 26877 23995 26911
rect 23937 26871 23995 26877
rect 24026 26868 24032 26920
rect 24084 26908 24090 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 24084 26880 24133 26908
rect 24084 26868 24090 26880
rect 24121 26877 24133 26880
rect 24167 26877 24179 26911
rect 24121 26871 24179 26877
rect 24854 26868 24860 26920
rect 24912 26868 24918 26920
rect 25682 26868 25688 26920
rect 25740 26908 25746 26920
rect 26142 26908 26148 26920
rect 25740 26880 26148 26908
rect 25740 26868 25746 26880
rect 26142 26868 26148 26880
rect 26200 26868 26206 26920
rect 26418 26868 26424 26920
rect 26476 26908 26482 26920
rect 26973 26911 27031 26917
rect 26973 26908 26985 26911
rect 26476 26880 26985 26908
rect 26476 26868 26482 26880
rect 26973 26877 26985 26880
rect 27019 26877 27031 26911
rect 26973 26871 27031 26877
rect 27614 26868 27620 26920
rect 27672 26908 27678 26920
rect 27985 26911 28043 26917
rect 27985 26908 27997 26911
rect 27672 26880 27997 26908
rect 27672 26868 27678 26880
rect 27985 26877 27997 26880
rect 28031 26877 28043 26911
rect 27985 26871 28043 26877
rect 23109 26843 23167 26849
rect 23109 26809 23121 26843
rect 23155 26840 23167 26843
rect 23569 26843 23627 26849
rect 23569 26840 23581 26843
rect 23155 26812 23581 26840
rect 23155 26809 23167 26812
rect 23109 26803 23167 26809
rect 23569 26809 23581 26812
rect 23615 26809 23627 26843
rect 23569 26803 23627 26809
rect 23676 26812 26372 26840
rect 23676 26772 23704 26812
rect 26344 26784 26372 26812
rect 21652 26744 23704 26772
rect 24302 26732 24308 26784
rect 24360 26772 24366 26784
rect 25041 26775 25099 26781
rect 25041 26772 25053 26775
rect 24360 26744 25053 26772
rect 24360 26732 24366 26744
rect 25041 26741 25053 26744
rect 25087 26741 25099 26775
rect 25041 26735 25099 26741
rect 26326 26732 26332 26784
rect 26384 26732 26390 26784
rect 26694 26732 26700 26784
rect 26752 26772 26758 26784
rect 26789 26775 26847 26781
rect 26789 26772 26801 26775
rect 26752 26744 26801 26772
rect 26752 26732 26758 26744
rect 26789 26741 26801 26744
rect 26835 26772 26847 26775
rect 27341 26775 27399 26781
rect 27341 26772 27353 26775
rect 26835 26744 27353 26772
rect 26835 26741 26847 26744
rect 26789 26735 26847 26741
rect 27341 26741 27353 26744
rect 27387 26741 27399 26775
rect 27341 26735 27399 26741
rect 27706 26732 27712 26784
rect 27764 26732 27770 26784
rect 28350 26732 28356 26784
rect 28408 26732 28414 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 2222 26528 2228 26580
rect 2280 26528 2286 26580
rect 2682 26528 2688 26580
rect 2740 26568 2746 26580
rect 2869 26571 2927 26577
rect 2869 26568 2881 26571
rect 2740 26540 2881 26568
rect 2740 26528 2746 26540
rect 2869 26537 2881 26540
rect 2915 26537 2927 26571
rect 2869 26531 2927 26537
rect 3329 26571 3387 26577
rect 3329 26537 3341 26571
rect 3375 26568 3387 26571
rect 3510 26568 3516 26580
rect 3375 26540 3516 26568
rect 3375 26537 3387 26540
rect 3329 26531 3387 26537
rect 3510 26528 3516 26540
rect 3568 26528 3574 26580
rect 4617 26571 4675 26577
rect 4617 26537 4629 26571
rect 4663 26568 4675 26571
rect 5074 26568 5080 26580
rect 4663 26540 5080 26568
rect 4663 26537 4675 26540
rect 4617 26531 4675 26537
rect 5074 26528 5080 26540
rect 5132 26528 5138 26580
rect 6822 26528 6828 26580
rect 6880 26568 6886 26580
rect 7653 26571 7711 26577
rect 7653 26568 7665 26571
rect 6880 26540 7665 26568
rect 6880 26528 6886 26540
rect 7653 26537 7665 26540
rect 7699 26537 7711 26571
rect 7653 26531 7711 26537
rect 8386 26528 8392 26580
rect 8444 26528 8450 26580
rect 8478 26528 8484 26580
rect 8536 26528 8542 26580
rect 9398 26528 9404 26580
rect 9456 26528 9462 26580
rect 9766 26528 9772 26580
rect 9824 26528 9830 26580
rect 11425 26571 11483 26577
rect 11425 26537 11437 26571
rect 11471 26568 11483 26571
rect 12710 26568 12716 26580
rect 11471 26540 12716 26568
rect 11471 26537 11483 26540
rect 11425 26531 11483 26537
rect 12710 26528 12716 26540
rect 12768 26528 12774 26580
rect 13170 26528 13176 26580
rect 13228 26568 13234 26580
rect 13228 26540 13492 26568
rect 13228 26528 13234 26540
rect 2240 26364 2268 26528
rect 5169 26503 5227 26509
rect 5169 26469 5181 26503
rect 5215 26500 5227 26503
rect 5215 26472 6592 26500
rect 5215 26469 5227 26472
rect 5169 26463 5227 26469
rect 5258 26392 5264 26444
rect 5316 26432 5322 26444
rect 5537 26435 5595 26441
rect 5537 26432 5549 26435
rect 5316 26404 5549 26432
rect 5316 26392 5322 26404
rect 5537 26401 5549 26404
rect 5583 26401 5595 26435
rect 5537 26395 5595 26401
rect 6178 26392 6184 26444
rect 6236 26392 6242 26444
rect 3053 26367 3111 26373
rect 3053 26364 3065 26367
rect 2240 26336 3065 26364
rect 3053 26333 3065 26336
rect 3099 26333 3111 26367
rect 3053 26327 3111 26333
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26333 3295 26367
rect 3237 26327 3295 26333
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26364 4583 26367
rect 4798 26364 4804 26376
rect 4571 26336 4804 26364
rect 4571 26333 4583 26336
rect 4525 26327 4583 26333
rect 3252 26240 3280 26327
rect 4798 26324 4804 26336
rect 4856 26364 4862 26376
rect 6564 26373 6592 26472
rect 6730 26460 6736 26512
rect 6788 26500 6794 26512
rect 7929 26503 7987 26509
rect 7929 26500 7941 26503
rect 6788 26472 7941 26500
rect 6788 26460 6794 26472
rect 7929 26469 7941 26472
rect 7975 26469 7987 26503
rect 7929 26463 7987 26469
rect 6914 26392 6920 26444
rect 6972 26392 6978 26444
rect 7006 26392 7012 26444
rect 7064 26392 7070 26444
rect 7101 26435 7159 26441
rect 7101 26401 7113 26435
rect 7147 26432 7159 26435
rect 8404 26432 8432 26528
rect 7147 26404 8432 26432
rect 8496 26432 8524 26528
rect 9125 26435 9183 26441
rect 9125 26432 9137 26435
rect 8496 26404 9137 26432
rect 7147 26401 7159 26404
rect 7101 26395 7159 26401
rect 9125 26401 9137 26404
rect 9171 26401 9183 26435
rect 9416 26432 9444 26528
rect 9784 26500 9812 26528
rect 12161 26503 12219 26509
rect 9784 26472 9996 26500
rect 9968 26441 9996 26472
rect 12161 26469 12173 26503
rect 12207 26500 12219 26503
rect 12434 26500 12440 26512
rect 12207 26472 12440 26500
rect 12207 26469 12219 26472
rect 12161 26463 12219 26469
rect 12434 26460 12440 26472
rect 12492 26460 12498 26512
rect 13464 26500 13492 26540
rect 13906 26528 13912 26580
rect 13964 26528 13970 26580
rect 14016 26540 15424 26568
rect 14016 26500 14044 26540
rect 13464 26472 14044 26500
rect 15396 26500 15424 26540
rect 15838 26528 15844 26580
rect 15896 26528 15902 26580
rect 18874 26568 18880 26580
rect 15948 26540 17632 26568
rect 15470 26500 15476 26512
rect 15396 26472 15476 26500
rect 15470 26460 15476 26472
rect 15528 26500 15534 26512
rect 15948 26500 15976 26540
rect 15528 26472 15976 26500
rect 16117 26503 16175 26509
rect 15528 26460 15534 26472
rect 16117 26469 16129 26503
rect 16163 26500 16175 26503
rect 17037 26503 17095 26509
rect 16163 26472 16620 26500
rect 16163 26469 16175 26472
rect 16117 26463 16175 26469
rect 9769 26435 9827 26441
rect 9769 26432 9781 26435
rect 9416 26404 9781 26432
rect 9125 26395 9183 26401
rect 9769 26401 9781 26404
rect 9815 26401 9827 26435
rect 9769 26395 9827 26401
rect 9953 26435 10011 26441
rect 9953 26401 9965 26435
rect 9999 26401 10011 26435
rect 12342 26432 12348 26444
rect 9953 26395 10011 26401
rect 10060 26404 12348 26432
rect 5353 26367 5411 26373
rect 5353 26364 5365 26367
rect 4856 26336 4936 26364
rect 4856 26324 4862 26336
rect 4908 26240 4936 26336
rect 5184 26336 5365 26364
rect 5184 26240 5212 26336
rect 5353 26333 5365 26336
rect 5399 26333 5411 26367
rect 5353 26327 5411 26333
rect 6549 26367 6607 26373
rect 6549 26333 6561 26367
rect 6595 26333 6607 26367
rect 6549 26327 6607 26333
rect 6825 26367 6883 26373
rect 6825 26333 6837 26367
rect 6871 26358 6883 26367
rect 7024 26364 7052 26392
rect 6932 26358 7052 26364
rect 6871 26336 7052 26358
rect 6871 26333 6960 26336
rect 6825 26330 6960 26333
rect 6825 26327 6883 26330
rect 7282 26324 7288 26376
rect 7340 26364 7346 26376
rect 7561 26367 7619 26373
rect 7561 26364 7573 26367
rect 7340 26336 7573 26364
rect 7340 26324 7346 26336
rect 7561 26333 7573 26336
rect 7607 26333 7619 26367
rect 7561 26327 7619 26333
rect 7650 26324 7656 26376
rect 7708 26364 7714 26376
rect 7837 26367 7895 26373
rect 7837 26364 7849 26367
rect 7708 26336 7849 26364
rect 7708 26324 7714 26336
rect 7837 26333 7849 26336
rect 7883 26333 7895 26367
rect 7837 26327 7895 26333
rect 7926 26324 7932 26376
rect 7984 26364 7990 26376
rect 8113 26367 8171 26373
rect 8113 26364 8125 26367
rect 7984 26336 8125 26364
rect 7984 26324 7990 26336
rect 8113 26333 8125 26336
rect 8159 26364 8171 26367
rect 8202 26364 8208 26376
rect 8159 26336 8208 26364
rect 8159 26333 8171 26336
rect 8113 26327 8171 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 8481 26367 8539 26373
rect 8481 26364 8493 26367
rect 8352 26336 8493 26364
rect 8352 26324 8358 26336
rect 8481 26333 8493 26336
rect 8527 26333 8539 26367
rect 8481 26327 8539 26333
rect 8757 26367 8815 26373
rect 8757 26333 8769 26367
rect 8803 26333 8815 26367
rect 8757 26327 8815 26333
rect 5629 26299 5687 26305
rect 5629 26265 5641 26299
rect 5675 26296 5687 26299
rect 8772 26296 8800 26327
rect 8846 26324 8852 26376
rect 8904 26324 8910 26376
rect 8938 26324 8944 26376
rect 8996 26364 9002 26376
rect 10060 26364 10088 26404
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 14461 26435 14519 26441
rect 14461 26432 14473 26435
rect 13547 26404 14473 26432
rect 10505 26367 10563 26373
rect 10505 26364 10517 26367
rect 8996 26336 10088 26364
rect 10152 26336 10517 26364
rect 8996 26324 9002 26336
rect 5675 26268 6132 26296
rect 5675 26265 5687 26268
rect 5629 26259 5687 26265
rect 3234 26188 3240 26240
rect 3292 26188 3298 26240
rect 4338 26188 4344 26240
rect 4396 26188 4402 26240
rect 4890 26188 4896 26240
rect 4948 26188 4954 26240
rect 5166 26188 5172 26240
rect 5224 26188 5230 26240
rect 6104 26228 6132 26268
rect 6748 26268 8800 26296
rect 8864 26296 8892 26324
rect 9582 26296 9588 26308
rect 8864 26268 9588 26296
rect 6365 26231 6423 26237
rect 6365 26228 6377 26231
rect 6104 26200 6377 26228
rect 6365 26197 6377 26200
rect 6411 26197 6423 26231
rect 6365 26191 6423 26197
rect 6641 26231 6699 26237
rect 6641 26197 6653 26231
rect 6687 26228 6699 26231
rect 6748 26228 6776 26268
rect 9582 26256 9588 26268
rect 9640 26296 9646 26308
rect 10152 26296 10180 26336
rect 10505 26333 10517 26336
rect 10551 26333 10563 26367
rect 10505 26327 10563 26333
rect 11238 26324 11244 26376
rect 11296 26324 11302 26376
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 13262 26364 13268 26376
rect 12584 26336 13268 26364
rect 12584 26324 12590 26336
rect 13262 26324 13268 26336
rect 13320 26364 13326 26376
rect 13547 26364 13575 26404
rect 14461 26401 14473 26404
rect 14507 26401 14519 26435
rect 14461 26395 14519 26401
rect 16393 26435 16451 26441
rect 16393 26401 16405 26435
rect 16439 26432 16451 26435
rect 16482 26432 16488 26444
rect 16439 26404 16488 26432
rect 16439 26401 16451 26404
rect 16393 26395 16451 26401
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 16592 26441 16620 26472
rect 17037 26469 17049 26503
rect 17083 26500 17095 26503
rect 17494 26500 17500 26512
rect 17083 26472 17500 26500
rect 17083 26469 17095 26472
rect 17037 26463 17095 26469
rect 17494 26460 17500 26472
rect 17552 26460 17558 26512
rect 17604 26500 17632 26540
rect 17972 26540 18880 26568
rect 17972 26500 18000 26540
rect 18874 26528 18880 26540
rect 18932 26528 18938 26580
rect 18969 26571 19027 26577
rect 18969 26537 18981 26571
rect 19015 26568 19027 26571
rect 19242 26568 19248 26580
rect 19015 26540 19248 26568
rect 19015 26537 19027 26540
rect 18969 26531 19027 26537
rect 19242 26528 19248 26540
rect 19300 26528 19306 26580
rect 19334 26528 19340 26580
rect 19392 26528 19398 26580
rect 19610 26528 19616 26580
rect 19668 26528 19674 26580
rect 20257 26571 20315 26577
rect 20257 26537 20269 26571
rect 20303 26568 20315 26571
rect 21082 26568 21088 26580
rect 20303 26540 21088 26568
rect 20303 26537 20315 26540
rect 20257 26531 20315 26537
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21266 26528 21272 26580
rect 21324 26528 21330 26580
rect 21358 26528 21364 26580
rect 21416 26528 21422 26580
rect 21542 26528 21548 26580
rect 21600 26528 21606 26580
rect 23658 26528 23664 26580
rect 23716 26528 23722 26580
rect 23845 26571 23903 26577
rect 23845 26537 23857 26571
rect 23891 26568 23903 26571
rect 24854 26568 24860 26580
rect 23891 26540 24860 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 26970 26568 26976 26580
rect 25424 26540 26976 26568
rect 19352 26500 19380 26528
rect 17604 26472 18000 26500
rect 18616 26472 19380 26500
rect 16577 26435 16635 26441
rect 16577 26401 16589 26435
rect 16623 26401 16635 26435
rect 16577 26395 16635 26401
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26432 17187 26435
rect 17678 26432 17684 26444
rect 17175 26404 17684 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 17678 26392 17684 26404
rect 17736 26392 17742 26444
rect 18616 26432 18644 26472
rect 17972 26404 18644 26432
rect 18693 26435 18751 26441
rect 13320 26336 13575 26364
rect 14185 26367 14243 26373
rect 13320 26324 13326 26336
rect 14185 26333 14197 26367
rect 14231 26333 14243 26367
rect 14185 26327 14243 26333
rect 14728 26367 14786 26373
rect 14728 26333 14740 26367
rect 14774 26364 14786 26367
rect 15194 26364 15200 26376
rect 14774 26336 15200 26364
rect 14774 26333 14786 26336
rect 14728 26327 14786 26333
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 9640 26268 10180 26296
rect 10428 26268 11621 26296
rect 9640 26256 9646 26268
rect 10428 26240 10456 26268
rect 11609 26265 11621 26268
rect 11655 26265 11667 26299
rect 11609 26259 11667 26265
rect 11698 26256 11704 26308
rect 11756 26256 11762 26308
rect 12618 26256 12624 26308
rect 12676 26296 12682 26308
rect 12774 26299 12832 26305
rect 12774 26296 12786 26299
rect 12676 26268 12786 26296
rect 12676 26256 12682 26268
rect 12774 26265 12786 26268
rect 12820 26265 12832 26299
rect 12774 26259 12832 26265
rect 14200 26240 14228 26327
rect 15194 26324 15200 26336
rect 15252 26324 15258 26376
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26364 16359 26367
rect 16666 26364 16672 26376
rect 16347 26336 16672 26364
rect 16347 26333 16359 26336
rect 16301 26327 16359 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17313 26367 17371 26373
rect 17313 26364 17325 26367
rect 17092 26336 17325 26364
rect 17092 26324 17098 26336
rect 17313 26333 17325 26336
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 17865 26367 17923 26373
rect 17865 26333 17877 26367
rect 17911 26364 17923 26367
rect 17972 26364 18000 26404
rect 18693 26401 18705 26435
rect 18739 26432 18751 26435
rect 19429 26435 19487 26441
rect 19429 26432 19441 26435
rect 18739 26404 19441 26432
rect 18739 26401 18751 26404
rect 18693 26395 18751 26401
rect 19429 26401 19441 26404
rect 19475 26401 19487 26435
rect 19429 26395 19487 26401
rect 17911 26336 18000 26364
rect 18049 26367 18107 26373
rect 17911 26333 17923 26336
rect 17865 26327 17923 26333
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 18601 26367 18659 26373
rect 18601 26364 18613 26367
rect 18049 26327 18107 26333
rect 18156 26336 18613 26364
rect 14277 26299 14335 26305
rect 14277 26265 14289 26299
rect 14323 26296 14335 26299
rect 14642 26296 14648 26308
rect 14323 26268 14648 26296
rect 14323 26265 14335 26268
rect 14277 26259 14335 26265
rect 14642 26256 14648 26268
rect 14700 26256 14706 26308
rect 17586 26256 17592 26308
rect 17644 26296 17650 26308
rect 18064 26296 18092 26327
rect 17644 26268 18092 26296
rect 17644 26256 17650 26268
rect 6687 26200 6776 26228
rect 8297 26231 8355 26237
rect 6687 26197 6699 26200
rect 6641 26191 6699 26197
rect 8297 26197 8309 26231
rect 8343 26228 8355 26231
rect 8386 26228 8392 26240
rect 8343 26200 8392 26228
rect 8343 26197 8355 26200
rect 8297 26191 8355 26197
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 8570 26188 8576 26240
rect 8628 26188 8634 26240
rect 10410 26188 10416 26240
rect 10468 26188 10474 26240
rect 11146 26188 11152 26240
rect 11204 26188 11210 26240
rect 14182 26188 14188 26240
rect 14240 26188 14246 26240
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 18156 26228 18184 26336
rect 18601 26333 18613 26336
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18877 26367 18935 26373
rect 18877 26333 18889 26367
rect 18923 26364 18935 26367
rect 19150 26364 19156 26376
rect 18923 26336 19156 26364
rect 18923 26333 18935 26336
rect 18877 26327 18935 26333
rect 19150 26324 19156 26336
rect 19208 26324 19214 26376
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 19628 26364 19656 26528
rect 19981 26503 20039 26509
rect 19981 26469 19993 26503
rect 20027 26469 20039 26503
rect 21376 26500 21404 26528
rect 19981 26463 20039 26469
rect 20640 26472 21404 26500
rect 19996 26432 20024 26463
rect 20640 26441 20668 26472
rect 20625 26435 20683 26441
rect 19996 26404 20484 26432
rect 19291 26336 19656 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 20162 26324 20168 26376
rect 20220 26324 20226 26376
rect 20456 26373 20484 26404
rect 20625 26401 20637 26435
rect 20671 26401 20683 26435
rect 20625 26395 20683 26401
rect 20809 26435 20867 26441
rect 20809 26401 20821 26435
rect 20855 26432 20867 26435
rect 21560 26432 21588 26528
rect 23293 26503 23351 26509
rect 23293 26469 23305 26503
rect 23339 26469 23351 26503
rect 23676 26500 23704 26528
rect 24673 26503 24731 26509
rect 23676 26472 24072 26500
rect 23293 26463 23351 26469
rect 20855 26404 21588 26432
rect 21821 26435 21879 26441
rect 20855 26401 20867 26404
rect 20809 26395 20867 26401
rect 21821 26401 21833 26435
rect 21867 26432 21879 26435
rect 22465 26435 22523 26441
rect 22465 26432 22477 26435
rect 21867 26404 22477 26432
rect 21867 26401 21879 26404
rect 21821 26395 21879 26401
rect 22465 26401 22477 26404
rect 22511 26401 22523 26435
rect 22465 26395 22523 26401
rect 22830 26392 22836 26444
rect 22888 26392 22894 26444
rect 23308 26432 23336 26463
rect 23308 26404 23796 26432
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26333 20499 26367
rect 20441 26327 20499 26333
rect 21266 26324 21272 26376
rect 21324 26364 21330 26376
rect 21637 26367 21695 26373
rect 21637 26364 21649 26367
rect 21324 26336 21649 26364
rect 21324 26324 21330 26336
rect 21637 26333 21649 26336
rect 21683 26333 21695 26367
rect 21637 26327 21695 26333
rect 22373 26367 22431 26373
rect 22373 26333 22385 26367
rect 22419 26364 22431 26367
rect 22848 26364 22876 26392
rect 22419 26336 22876 26364
rect 22419 26333 22431 26336
rect 22373 26327 22431 26333
rect 23382 26324 23388 26376
rect 23440 26364 23446 26376
rect 23768 26373 23796 26404
rect 24044 26373 24072 26472
rect 24673 26469 24685 26503
rect 24719 26500 24731 26503
rect 24946 26500 24952 26512
rect 24719 26472 24952 26500
rect 24719 26469 24731 26472
rect 24673 26463 24731 26469
rect 24946 26460 24952 26472
rect 25004 26460 25010 26512
rect 25038 26392 25044 26444
rect 25096 26432 25102 26444
rect 25424 26441 25452 26540
rect 26970 26528 26976 26540
rect 27028 26528 27034 26580
rect 27614 26528 27620 26580
rect 27672 26528 27678 26580
rect 27706 26528 27712 26580
rect 27764 26528 27770 26580
rect 27798 26528 27804 26580
rect 27856 26568 27862 26580
rect 28169 26571 28227 26577
rect 28169 26568 28181 26571
rect 27856 26540 28181 26568
rect 27856 26528 27862 26540
rect 28169 26537 28181 26540
rect 28215 26537 28227 26571
rect 28169 26531 28227 26537
rect 27632 26500 27660 26528
rect 26160 26472 26556 26500
rect 26160 26444 26188 26472
rect 25409 26435 25467 26441
rect 25409 26432 25421 26435
rect 25096 26404 25421 26432
rect 25096 26392 25102 26404
rect 25409 26401 25421 26404
rect 25455 26401 25467 26435
rect 25409 26395 25467 26401
rect 26142 26392 26148 26444
rect 26200 26392 26206 26444
rect 26418 26392 26424 26444
rect 26476 26392 26482 26444
rect 23477 26367 23535 26373
rect 23477 26364 23489 26367
rect 23440 26336 23489 26364
rect 23440 26324 23446 26336
rect 23477 26333 23489 26336
rect 23523 26333 23535 26367
rect 23477 26327 23535 26333
rect 23753 26367 23811 26373
rect 23753 26333 23765 26367
rect 23799 26333 23811 26367
rect 23753 26327 23811 26333
rect 24029 26367 24087 26373
rect 24029 26333 24041 26367
rect 24075 26333 24087 26367
rect 24029 26327 24087 26333
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 25130 26364 25136 26376
rect 24903 26336 25136 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 25130 26324 25136 26336
rect 25188 26324 25194 26376
rect 25590 26324 25596 26376
rect 25648 26324 25654 26376
rect 25774 26324 25780 26376
rect 25832 26364 25838 26376
rect 26237 26367 26295 26373
rect 26237 26364 26249 26367
rect 25832 26336 26249 26364
rect 25832 26324 25838 26336
rect 26237 26333 26249 26336
rect 26283 26333 26295 26367
rect 26237 26327 26295 26333
rect 18506 26256 18512 26308
rect 18564 26296 18570 26308
rect 19889 26299 19947 26305
rect 19889 26296 19901 26299
rect 18564 26268 19901 26296
rect 18564 26256 18570 26268
rect 19889 26265 19901 26268
rect 19935 26265 19947 26299
rect 26436 26296 26464 26392
rect 19889 26259 19947 26265
rect 19996 26268 26464 26296
rect 26528 26296 26556 26472
rect 27356 26472 27660 26500
rect 26605 26435 26663 26441
rect 26605 26401 26617 26435
rect 26651 26432 26663 26435
rect 26694 26432 26700 26444
rect 26651 26404 26700 26432
rect 26651 26401 26663 26404
rect 26605 26395 26663 26401
rect 26694 26392 26700 26404
rect 26752 26392 26758 26444
rect 27356 26441 27384 26472
rect 27341 26435 27399 26441
rect 27341 26401 27353 26435
rect 27387 26401 27399 26435
rect 27341 26395 27399 26401
rect 27525 26435 27583 26441
rect 27525 26401 27537 26435
rect 27571 26432 27583 26435
rect 27724 26432 27752 26528
rect 28074 26460 28080 26512
rect 28132 26500 28138 26512
rect 28353 26503 28411 26509
rect 28353 26500 28365 26503
rect 28132 26472 28365 26500
rect 28132 26460 28138 26472
rect 28353 26469 28365 26472
rect 28399 26469 28411 26503
rect 28353 26463 28411 26469
rect 27571 26404 27752 26432
rect 27571 26401 27583 26404
rect 27525 26395 27583 26401
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26364 26847 26367
rect 27062 26364 27068 26376
rect 26835 26336 27068 26364
rect 26835 26333 26847 26336
rect 26789 26327 26847 26333
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 28077 26367 28135 26373
rect 28077 26364 28089 26367
rect 27172 26336 28089 26364
rect 27172 26296 27200 26336
rect 28077 26333 28089 26336
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 28534 26324 28540 26376
rect 28592 26324 28598 26376
rect 26528 26268 27200 26296
rect 27249 26299 27307 26305
rect 17000 26200 18184 26228
rect 17000 26188 17006 26200
rect 18874 26188 18880 26240
rect 18932 26228 18938 26240
rect 19996 26228 20024 26268
rect 27249 26265 27261 26299
rect 27295 26296 27307 26299
rect 27706 26296 27712 26308
rect 27295 26268 27712 26296
rect 27295 26265 27307 26268
rect 27249 26259 27307 26265
rect 27706 26256 27712 26268
rect 27764 26296 27770 26308
rect 27985 26299 28043 26305
rect 27985 26296 27997 26299
rect 27764 26268 27997 26296
rect 27764 26256 27770 26268
rect 27985 26265 27997 26268
rect 28031 26265 28043 26299
rect 27985 26259 28043 26265
rect 18932 26200 20024 26228
rect 18932 26188 18938 26200
rect 22278 26188 22284 26240
rect 22336 26188 22342 26240
rect 23566 26188 23572 26240
rect 23624 26188 23630 26240
rect 25130 26188 25136 26240
rect 25188 26228 25194 26240
rect 25774 26228 25780 26240
rect 25188 26200 25780 26228
rect 25188 26188 25194 26200
rect 25774 26188 25780 26200
rect 25832 26188 25838 26240
rect 26050 26188 26056 26240
rect 26108 26188 26114 26240
rect 26234 26188 26240 26240
rect 26292 26228 26298 26240
rect 26329 26231 26387 26237
rect 26329 26228 26341 26231
rect 26292 26200 26341 26228
rect 26292 26188 26298 26200
rect 26329 26197 26341 26200
rect 26375 26197 26387 26231
rect 26329 26191 26387 26197
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 1765 26027 1823 26033
rect 1765 25993 1777 26027
rect 1811 25993 1823 26027
rect 1765 25987 1823 25993
rect 1780 25956 1808 25987
rect 2314 25984 2320 26036
rect 2372 26024 2378 26036
rect 5261 26027 5319 26033
rect 2372 25996 2728 26024
rect 2372 25984 2378 25996
rect 2700 25956 2728 25996
rect 5261 25993 5273 26027
rect 5307 26024 5319 26027
rect 5902 26024 5908 26036
rect 5307 25996 5908 26024
rect 5307 25993 5319 25996
rect 5261 25987 5319 25993
rect 5902 25984 5908 25996
rect 5960 25984 5966 26036
rect 6362 26024 6368 26036
rect 6104 25996 6368 26024
rect 4985 25959 5043 25965
rect 1780 25928 2636 25956
rect 1578 25848 1584 25900
rect 1636 25848 1642 25900
rect 2608 25897 2636 25928
rect 2700 25928 4936 25956
rect 2700 25897 2728 25928
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25888 2007 25891
rect 2225 25891 2283 25897
rect 1995 25860 2176 25888
rect 1995 25857 2007 25860
rect 1949 25851 2007 25857
rect 1394 25644 1400 25696
rect 1452 25644 1458 25696
rect 2038 25644 2044 25696
rect 2096 25644 2102 25696
rect 2148 25684 2176 25860
rect 2225 25857 2237 25891
rect 2271 25857 2283 25891
rect 2225 25851 2283 25857
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25857 2651 25891
rect 2593 25851 2651 25857
rect 2685 25891 2743 25897
rect 2685 25857 2697 25891
rect 2731 25857 2743 25891
rect 2685 25851 2743 25857
rect 2240 25820 2268 25851
rect 2498 25820 2504 25832
rect 2240 25792 2504 25820
rect 2498 25780 2504 25792
rect 2556 25780 2562 25832
rect 2869 25823 2927 25829
rect 2869 25820 2881 25823
rect 2746 25792 2881 25820
rect 2409 25755 2467 25761
rect 2409 25721 2421 25755
rect 2455 25752 2467 25755
rect 2746 25752 2774 25792
rect 2869 25789 2881 25792
rect 2915 25789 2927 25823
rect 2869 25783 2927 25789
rect 3418 25780 3424 25832
rect 3476 25780 3482 25832
rect 3602 25780 3608 25832
rect 3660 25780 3666 25832
rect 4341 25823 4399 25829
rect 4341 25820 4353 25823
rect 3804 25792 4353 25820
rect 3804 25761 3832 25792
rect 4341 25789 4353 25792
rect 4387 25789 4399 25823
rect 4341 25783 4399 25789
rect 4525 25823 4583 25829
rect 4525 25789 4537 25823
rect 4571 25789 4583 25823
rect 4525 25783 4583 25789
rect 2455 25724 2774 25752
rect 3329 25755 3387 25761
rect 2455 25721 2467 25724
rect 2409 25715 2467 25721
rect 3329 25721 3341 25755
rect 3375 25752 3387 25755
rect 3789 25755 3847 25761
rect 3789 25752 3801 25755
rect 3375 25724 3801 25752
rect 3375 25721 3387 25724
rect 3329 25715 3387 25721
rect 3789 25721 3801 25724
rect 3835 25721 3847 25755
rect 3789 25715 3847 25721
rect 3970 25712 3976 25764
rect 4028 25752 4034 25764
rect 4540 25752 4568 25783
rect 4028 25724 4568 25752
rect 4908 25752 4936 25928
rect 4985 25925 4997 25959
rect 5031 25956 5043 25959
rect 6104 25956 6132 25996
rect 6362 25984 6368 25996
rect 6420 25984 6426 26036
rect 7282 25984 7288 26036
rect 7340 26024 7346 26036
rect 8021 26027 8079 26033
rect 8021 26024 8033 26027
rect 7340 25996 8033 26024
rect 7340 25984 7346 25996
rect 8021 25993 8033 25996
rect 8067 25993 8079 26027
rect 8021 25987 8079 25993
rect 10410 25984 10416 26036
rect 10468 25984 10474 26036
rect 11333 26027 11391 26033
rect 11333 25993 11345 26027
rect 11379 26024 11391 26027
rect 12618 26024 12624 26036
rect 11379 25996 12624 26024
rect 11379 25993 11391 25996
rect 11333 25987 11391 25993
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 14366 25984 14372 26036
rect 14424 26024 14430 26036
rect 14550 26024 14556 26036
rect 14424 25996 14556 26024
rect 14424 25984 14430 25996
rect 14550 25984 14556 25996
rect 14608 26024 14614 26036
rect 21542 26024 21548 26036
rect 14608 25996 21548 26024
rect 14608 25984 14614 25996
rect 21542 25984 21548 25996
rect 21600 25984 21606 26036
rect 22278 25984 22284 26036
rect 22336 26024 22342 26036
rect 22465 26027 22523 26033
rect 22465 26024 22477 26027
rect 22336 25996 22477 26024
rect 22336 25984 22342 25996
rect 22465 25993 22477 25996
rect 22511 25993 22523 26027
rect 22465 25987 22523 25993
rect 5031 25928 6132 25956
rect 5031 25925 5043 25928
rect 4985 25919 5043 25925
rect 6178 25916 6184 25968
rect 6236 25956 6242 25968
rect 6457 25959 6515 25965
rect 6457 25956 6469 25959
rect 6236 25928 6469 25956
rect 6236 25916 6242 25928
rect 6457 25925 6469 25928
rect 6503 25925 6515 25959
rect 6457 25919 6515 25925
rect 6546 25916 6552 25968
rect 6604 25916 6610 25968
rect 8294 25956 8300 25968
rect 7944 25928 8300 25956
rect 5166 25888 5172 25900
rect 5224 25897 5230 25900
rect 7944 25897 7972 25928
rect 8294 25916 8300 25928
rect 8352 25916 8358 25968
rect 14182 25956 14188 25968
rect 11808 25928 14188 25956
rect 5135 25860 5172 25888
rect 5166 25848 5172 25860
rect 5224 25888 5235 25897
rect 5537 25891 5595 25897
rect 5537 25888 5549 25891
rect 5224 25860 5549 25888
rect 5224 25851 5235 25860
rect 5537 25857 5549 25860
rect 5583 25857 5595 25891
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 5537 25851 5595 25857
rect 7208 25860 7941 25888
rect 5224 25848 5230 25851
rect 6454 25780 6460 25832
rect 6512 25820 6518 25832
rect 7208 25829 7236 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25888 8539 25891
rect 8570 25888 8576 25900
rect 8527 25860 8576 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 9582 25888 9588 25900
rect 9048 25860 9588 25888
rect 9048 25829 9076 25860
rect 9582 25848 9588 25860
rect 9640 25848 9646 25900
rect 9674 25848 9680 25900
rect 9732 25888 9738 25900
rect 11808 25897 11836 25928
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 14274 25916 14280 25968
rect 14332 25956 14338 25968
rect 20162 25956 20168 25968
rect 14332 25928 14596 25956
rect 14332 25916 14338 25928
rect 9953 25891 10011 25897
rect 9953 25888 9965 25891
rect 9732 25860 9965 25888
rect 9732 25848 9738 25860
rect 9953 25857 9965 25860
rect 9999 25857 10011 25891
rect 9953 25851 10011 25857
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25857 11851 25891
rect 11793 25851 11851 25857
rect 12342 25848 12348 25900
rect 12400 25848 12406 25900
rect 14568 25897 14596 25928
rect 14660 25928 16896 25956
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25857 14611 25891
rect 14553 25851 14611 25857
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6512 25792 7205 25820
rect 6512 25780 6518 25792
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 8297 25823 8355 25829
rect 8297 25820 8309 25823
rect 7193 25783 7251 25789
rect 7760 25792 8309 25820
rect 4908 25724 6960 25752
rect 4028 25712 4034 25724
rect 3234 25684 3240 25696
rect 2148 25656 3240 25684
rect 3234 25644 3240 25656
rect 3292 25644 3298 25696
rect 6086 25644 6092 25696
rect 6144 25644 6150 25696
rect 6932 25684 6960 25724
rect 7006 25712 7012 25764
rect 7064 25712 7070 25764
rect 7760 25684 7788 25792
rect 8297 25789 8309 25792
rect 8343 25789 8355 25823
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 8297 25783 8355 25789
rect 8496 25792 9045 25820
rect 6932 25656 7788 25684
rect 7834 25644 7840 25696
rect 7892 25644 7898 25696
rect 8312 25684 8340 25783
rect 8496 25764 8524 25792
rect 9033 25789 9045 25792
rect 9079 25789 9091 25823
rect 9033 25783 9091 25789
rect 9214 25780 9220 25832
rect 9272 25780 9278 25832
rect 9769 25823 9827 25829
rect 9769 25820 9781 25823
rect 9416 25792 9781 25820
rect 8478 25712 8484 25764
rect 8536 25712 8542 25764
rect 9416 25761 9444 25792
rect 9769 25789 9781 25792
rect 9815 25789 9827 25823
rect 9769 25783 9827 25789
rect 10781 25823 10839 25829
rect 10781 25789 10793 25823
rect 10827 25789 10839 25823
rect 10781 25783 10839 25789
rect 8941 25755 8999 25761
rect 8941 25721 8953 25755
rect 8987 25752 8999 25755
rect 9401 25755 9459 25761
rect 9401 25752 9413 25755
rect 8987 25724 9413 25752
rect 8987 25721 8999 25724
rect 8941 25715 8999 25721
rect 9401 25721 9413 25724
rect 9447 25721 9459 25755
rect 10796 25752 10824 25783
rect 12434 25780 12440 25832
rect 12492 25780 12498 25832
rect 12621 25823 12679 25829
rect 12621 25789 12633 25823
rect 12667 25820 12679 25823
rect 12710 25820 12716 25832
rect 12667 25792 12716 25820
rect 12667 25789 12679 25792
rect 12621 25783 12679 25789
rect 12710 25780 12716 25792
rect 12768 25780 12774 25832
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 12897 25823 12955 25829
rect 12897 25820 12909 25823
rect 12860 25792 12909 25820
rect 12860 25780 12866 25792
rect 12897 25789 12909 25792
rect 12943 25820 12955 25823
rect 14660 25820 14688 25928
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 15286 25888 15292 25900
rect 15243 25860 15292 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15378 25848 15384 25900
rect 15436 25888 15442 25900
rect 16868 25897 16896 25928
rect 19996 25928 20168 25956
rect 15933 25891 15991 25897
rect 15933 25888 15945 25891
rect 15436 25860 15945 25888
rect 15436 25848 15442 25860
rect 15933 25857 15945 25860
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 16899 25860 17141 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 17129 25857 17141 25860
rect 17175 25857 17187 25891
rect 17129 25851 17187 25857
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25888 17279 25891
rect 17267 25860 17448 25888
rect 17267 25857 17279 25860
rect 17221 25851 17279 25857
rect 17420 25832 17448 25860
rect 17494 25848 17500 25900
rect 17552 25888 17558 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17552 25860 17601 25888
rect 17552 25848 17558 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 18506 25848 18512 25900
rect 18564 25848 18570 25900
rect 19996 25897 20024 25928
rect 20162 25916 20168 25928
rect 20220 25956 20226 25968
rect 21450 25956 21456 25968
rect 20220 25928 21456 25956
rect 20220 25916 20226 25928
rect 21284 25900 21312 25928
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 22480 25956 22508 25987
rect 24946 25984 24952 26036
rect 25004 25984 25010 26036
rect 25041 26027 25099 26033
rect 25041 25993 25053 26027
rect 25087 26024 25099 26027
rect 25590 26024 25596 26036
rect 25087 25996 25596 26024
rect 25087 25993 25099 25996
rect 25041 25987 25099 25993
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 26050 25984 26056 26036
rect 26108 26024 26114 26036
rect 26145 26027 26203 26033
rect 26145 26024 26157 26027
rect 26108 25996 26157 26024
rect 26108 25984 26114 25996
rect 26145 25993 26157 25996
rect 26191 25993 26203 26027
rect 26145 25987 26203 25993
rect 22480 25928 22968 25956
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25857 20039 25891
rect 19981 25851 20039 25857
rect 20257 25891 20315 25897
rect 20257 25857 20269 25891
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 12943 25792 14688 25820
rect 12943 25789 12955 25792
rect 12897 25783 12955 25789
rect 14734 25780 14740 25832
rect 14792 25820 14798 25832
rect 15013 25823 15071 25829
rect 15013 25820 15025 25823
rect 14792 25792 15025 25820
rect 14792 25780 14798 25792
rect 15013 25789 15025 25792
rect 15059 25789 15071 25823
rect 15013 25783 15071 25789
rect 15746 25780 15752 25832
rect 15804 25780 15810 25832
rect 17402 25780 17408 25832
rect 17460 25780 17466 25832
rect 17770 25780 17776 25832
rect 17828 25780 17834 25832
rect 18690 25780 18696 25832
rect 18748 25780 18754 25832
rect 20272 25820 20300 25851
rect 21266 25848 21272 25900
rect 21324 25848 21330 25900
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22741 25891 22799 25897
rect 22741 25888 22753 25891
rect 21968 25860 22753 25888
rect 21968 25848 21974 25860
rect 22741 25857 22753 25860
rect 22787 25888 22799 25891
rect 22830 25888 22836 25900
rect 22787 25860 22836 25888
rect 22787 25857 22799 25860
rect 22741 25851 22799 25857
rect 22830 25848 22836 25860
rect 22888 25848 22894 25900
rect 22940 25897 22968 25928
rect 22925 25891 22983 25897
rect 22925 25857 22937 25891
rect 22971 25857 22983 25891
rect 22925 25851 22983 25857
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 23845 25891 23903 25897
rect 23845 25888 23857 25891
rect 23624 25860 23857 25888
rect 23624 25848 23630 25860
rect 23845 25857 23857 25860
rect 23891 25857 23903 25891
rect 23845 25851 23903 25857
rect 24394 25848 24400 25900
rect 24452 25848 24458 25900
rect 24964 25888 24992 25984
rect 26160 25956 26188 25987
rect 26160 25928 27016 25956
rect 25225 25891 25283 25897
rect 25225 25888 25237 25891
rect 24964 25860 25237 25888
rect 25225 25857 25237 25860
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 26326 25848 26332 25900
rect 26384 25848 26390 25900
rect 26988 25897 27016 25928
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27706 25848 27712 25900
rect 27764 25848 27770 25900
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25888 27951 25891
rect 28350 25888 28356 25900
rect 27939 25860 28356 25888
rect 27939 25857 27951 25860
rect 27893 25851 27951 25857
rect 28350 25848 28356 25860
rect 28408 25848 28414 25900
rect 19812 25792 20300 25820
rect 13906 25752 13912 25764
rect 10796 25724 13912 25752
rect 9401 25715 9459 25721
rect 13906 25712 13912 25724
rect 13964 25712 13970 25764
rect 19812 25761 19840 25792
rect 20530 25780 20536 25832
rect 20588 25780 20594 25832
rect 20717 25823 20775 25829
rect 20717 25789 20729 25823
rect 20763 25789 20775 25823
rect 20717 25783 20775 25789
rect 19797 25755 19855 25761
rect 14292 25724 19334 25752
rect 13170 25684 13176 25696
rect 8312 25656 13176 25684
rect 13170 25644 13176 25656
rect 13228 25684 13234 25696
rect 14292 25684 14320 25724
rect 13228 25656 14320 25684
rect 14369 25687 14427 25693
rect 13228 25644 13234 25656
rect 14369 25653 14381 25687
rect 14415 25684 14427 25687
rect 15286 25684 15292 25696
rect 14415 25656 15292 25684
rect 14415 25653 14427 25656
rect 14369 25647 14427 25653
rect 15286 25644 15292 25656
rect 15344 25644 15350 25696
rect 15657 25687 15715 25693
rect 15657 25653 15669 25687
rect 15703 25684 15715 25687
rect 16114 25684 16120 25696
rect 15703 25656 16120 25684
rect 15703 25653 15715 25656
rect 15657 25647 15715 25653
rect 16114 25644 16120 25656
rect 16172 25644 16178 25696
rect 16666 25644 16672 25696
rect 16724 25644 16730 25696
rect 16945 25687 17003 25693
rect 16945 25653 16957 25687
rect 16991 25684 17003 25687
rect 17218 25684 17224 25696
rect 16991 25656 17224 25684
rect 16991 25653 17003 25656
rect 16945 25647 17003 25653
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 17310 25644 17316 25696
rect 17368 25644 17374 25696
rect 18233 25687 18291 25693
rect 18233 25653 18245 25687
rect 18279 25684 18291 25687
rect 18782 25684 18788 25696
rect 18279 25656 18788 25684
rect 18279 25653 18291 25656
rect 18233 25647 18291 25653
rect 18782 25644 18788 25656
rect 18840 25684 18846 25696
rect 18877 25687 18935 25693
rect 18877 25684 18889 25687
rect 18840 25656 18889 25684
rect 18840 25644 18846 25656
rect 18877 25653 18889 25656
rect 18923 25653 18935 25687
rect 19306 25684 19334 25724
rect 19797 25721 19809 25755
rect 19843 25721 19855 25755
rect 19797 25715 19855 25721
rect 20073 25755 20131 25761
rect 20073 25721 20085 25755
rect 20119 25752 20131 25755
rect 20732 25752 20760 25783
rect 21174 25780 21180 25832
rect 21232 25820 21238 25832
rect 21821 25823 21879 25829
rect 21821 25820 21833 25823
rect 21232 25792 21833 25820
rect 21232 25780 21238 25792
rect 21821 25789 21833 25792
rect 21867 25789 21879 25823
rect 21821 25783 21879 25789
rect 22002 25780 22008 25832
rect 22060 25780 22066 25832
rect 23106 25780 23112 25832
rect 23164 25780 23170 25832
rect 23661 25823 23719 25829
rect 23661 25789 23673 25823
rect 23707 25820 23719 25823
rect 24302 25820 24308 25832
rect 23707 25792 24308 25820
rect 23707 25789 23719 25792
rect 23661 25783 23719 25789
rect 24302 25780 24308 25792
rect 24360 25780 24366 25832
rect 25501 25823 25559 25829
rect 25501 25789 25513 25823
rect 25547 25789 25559 25823
rect 25501 25783 25559 25789
rect 25685 25823 25743 25829
rect 25685 25789 25697 25823
rect 25731 25820 25743 25823
rect 26234 25820 26240 25832
rect 25731 25792 26240 25820
rect 25731 25789 25743 25792
rect 25685 25783 25743 25789
rect 25516 25752 25544 25783
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 26510 25780 26516 25832
rect 26568 25820 26574 25832
rect 27157 25823 27215 25829
rect 27157 25820 27169 25823
rect 26568 25792 27169 25820
rect 26568 25780 26574 25792
rect 27157 25789 27169 25792
rect 27203 25789 27215 25823
rect 27157 25783 27215 25789
rect 26605 25755 26663 25761
rect 26605 25752 26617 25755
rect 20119 25724 20760 25752
rect 22066 25724 26617 25752
rect 20119 25721 20131 25724
rect 20073 25715 20131 25721
rect 20346 25684 20352 25696
rect 19306 25656 20352 25684
rect 18877 25647 18935 25653
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 21358 25644 21364 25696
rect 21416 25644 21422 25696
rect 21542 25644 21548 25696
rect 21600 25684 21606 25696
rect 22066 25684 22094 25724
rect 26605 25721 26617 25724
rect 26651 25721 26663 25755
rect 26605 25715 26663 25721
rect 21600 25656 22094 25684
rect 21600 25644 21606 25656
rect 22554 25644 22560 25696
rect 22612 25644 22618 25696
rect 23569 25687 23627 25693
rect 23569 25653 23581 25687
rect 23615 25684 23627 25687
rect 24026 25684 24032 25696
rect 23615 25656 24032 25684
rect 23615 25653 23627 25656
rect 23569 25647 23627 25653
rect 24026 25644 24032 25656
rect 24084 25644 24090 25696
rect 24578 25644 24584 25696
rect 24636 25644 24642 25696
rect 27338 25644 27344 25696
rect 27396 25644 27402 25696
rect 27982 25644 27988 25696
rect 28040 25684 28046 25696
rect 28077 25687 28135 25693
rect 28077 25684 28089 25687
rect 28040 25656 28089 25684
rect 28040 25644 28046 25656
rect 28077 25653 28089 25656
rect 28123 25653 28135 25687
rect 28077 25647 28135 25653
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 1394 25440 1400 25492
rect 1452 25440 1458 25492
rect 2038 25440 2044 25492
rect 2096 25440 2102 25492
rect 3513 25483 3571 25489
rect 3513 25449 3525 25483
rect 3559 25480 3571 25483
rect 3602 25480 3608 25492
rect 3559 25452 3608 25480
rect 3559 25449 3571 25452
rect 3513 25443 3571 25449
rect 3602 25440 3608 25452
rect 3660 25440 3666 25492
rect 3970 25440 3976 25492
rect 4028 25440 4034 25492
rect 4801 25483 4859 25489
rect 4801 25449 4813 25483
rect 4847 25480 4859 25483
rect 6546 25480 6552 25492
rect 4847 25452 6552 25480
rect 4847 25449 4859 25452
rect 4801 25443 4859 25449
rect 6546 25440 6552 25452
rect 6604 25440 6610 25492
rect 7834 25440 7840 25492
rect 7892 25440 7898 25492
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 9214 25480 9220 25492
rect 8435 25452 9220 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 9214 25440 9220 25452
rect 9272 25440 9278 25492
rect 9861 25483 9919 25489
rect 9861 25449 9873 25483
rect 9907 25480 9919 25483
rect 11698 25480 11704 25492
rect 9907 25452 11704 25480
rect 9907 25449 9919 25452
rect 9861 25443 9919 25449
rect 11698 25440 11704 25452
rect 11756 25440 11762 25492
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 15470 25480 15476 25492
rect 13964 25452 15476 25480
rect 13964 25440 13970 25452
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 16114 25440 16120 25492
rect 16172 25440 16178 25492
rect 17034 25440 17040 25492
rect 17092 25440 17098 25492
rect 17589 25483 17647 25489
rect 17589 25449 17601 25483
rect 17635 25480 17647 25483
rect 17770 25480 17776 25492
rect 17635 25452 17776 25480
rect 17635 25449 17647 25452
rect 17589 25443 17647 25449
rect 17770 25440 17776 25452
rect 17828 25440 17834 25492
rect 18509 25483 18567 25489
rect 18509 25449 18521 25483
rect 18555 25449 18567 25483
rect 18509 25443 18567 25449
rect 1412 25276 1440 25440
rect 2056 25344 2084 25440
rect 2498 25372 2504 25424
rect 2556 25412 2562 25424
rect 2556 25384 3188 25412
rect 2556 25372 2562 25384
rect 2056 25316 2544 25344
rect 1581 25279 1639 25285
rect 1581 25276 1593 25279
rect 1412 25248 1593 25276
rect 1581 25245 1593 25248
rect 1627 25245 1639 25279
rect 1581 25239 1639 25245
rect 1670 25236 1676 25288
rect 1728 25276 1734 25288
rect 2516 25285 2544 25316
rect 2041 25279 2099 25285
rect 2041 25276 2053 25279
rect 1728 25248 2053 25276
rect 1728 25236 1734 25248
rect 2041 25245 2053 25248
rect 2087 25245 2099 25279
rect 2041 25239 2099 25245
rect 2501 25279 2559 25285
rect 2501 25245 2513 25279
rect 2547 25245 2559 25279
rect 2501 25239 2559 25245
rect 2590 25236 2596 25288
rect 2648 25236 2654 25288
rect 2866 25236 2872 25288
rect 2924 25236 2930 25288
rect 3160 25285 3188 25384
rect 6454 25372 6460 25424
rect 6512 25372 6518 25424
rect 3878 25304 3884 25356
rect 3936 25344 3942 25356
rect 5077 25347 5135 25353
rect 5077 25344 5089 25347
rect 3936 25316 5089 25344
rect 3936 25304 3942 25316
rect 5077 25313 5089 25316
rect 5123 25313 5135 25347
rect 6825 25347 6883 25353
rect 6825 25344 6837 25347
rect 5077 25307 5135 25313
rect 6104 25316 6837 25344
rect 3145 25279 3203 25285
rect 3145 25245 3157 25279
rect 3191 25245 3203 25279
rect 3421 25279 3479 25285
rect 3421 25276 3433 25279
rect 3145 25239 3203 25245
rect 3344 25248 3433 25276
rect 2685 25211 2743 25217
rect 2685 25177 2697 25211
rect 2731 25208 2743 25211
rect 3050 25208 3056 25220
rect 2731 25180 3056 25208
rect 2731 25177 2743 25180
rect 2685 25171 2743 25177
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 3344 25152 3372 25248
rect 3421 25245 3433 25248
rect 3467 25245 3479 25279
rect 3421 25239 3479 25245
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25276 4215 25279
rect 4338 25276 4344 25288
rect 4203 25248 4344 25276
rect 4203 25245 4215 25248
rect 4157 25239 4215 25245
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 4433 25279 4491 25285
rect 4433 25245 4445 25279
rect 4479 25245 4491 25279
rect 4433 25239 4491 25245
rect 4709 25279 4767 25285
rect 4709 25245 4721 25279
rect 4755 25276 4767 25279
rect 4798 25276 4804 25288
rect 4755 25248 4804 25276
rect 4755 25245 4767 25248
rect 4709 25239 4767 25245
rect 4448 25208 4476 25239
rect 4798 25236 4804 25248
rect 4856 25236 4862 25288
rect 4890 25236 4896 25288
rect 4948 25236 4954 25288
rect 4985 25279 5043 25285
rect 4985 25245 4997 25279
rect 5031 25245 5043 25279
rect 5092 25276 5120 25307
rect 6104 25276 6132 25316
rect 6825 25313 6837 25316
rect 6871 25313 6883 25347
rect 6825 25307 6883 25313
rect 5092 25248 6132 25276
rect 4985 25239 5043 25245
rect 4908 25208 4936 25236
rect 4448 25180 4936 25208
rect 1673 25143 1731 25149
rect 1673 25109 1685 25143
rect 1719 25140 1731 25143
rect 1946 25140 1952 25152
rect 1719 25112 1952 25140
rect 1719 25109 1731 25112
rect 1673 25103 1731 25109
rect 1946 25100 1952 25112
rect 2004 25100 2010 25152
rect 2038 25100 2044 25152
rect 2096 25140 2102 25152
rect 2133 25143 2191 25149
rect 2133 25140 2145 25143
rect 2096 25112 2145 25140
rect 2096 25100 2102 25112
rect 2133 25109 2145 25112
rect 2179 25109 2191 25143
rect 2133 25103 2191 25109
rect 2317 25143 2375 25149
rect 2317 25109 2329 25143
rect 2363 25140 2375 25143
rect 2774 25140 2780 25152
rect 2363 25112 2780 25140
rect 2363 25109 2375 25112
rect 2317 25103 2375 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 2958 25100 2964 25152
rect 3016 25100 3022 25152
rect 3234 25100 3240 25152
rect 3292 25100 3298 25152
rect 3326 25100 3332 25152
rect 3384 25100 3390 25152
rect 4246 25100 4252 25152
rect 4304 25100 4310 25152
rect 4522 25100 4528 25152
rect 4580 25100 4586 25152
rect 5000 25140 5028 25239
rect 6730 25236 6736 25288
rect 6788 25236 6794 25288
rect 7092 25279 7150 25285
rect 7092 25245 7104 25279
rect 7138 25276 7150 25279
rect 7852 25276 7880 25440
rect 8573 25415 8631 25421
rect 8573 25381 8585 25415
rect 8619 25412 8631 25415
rect 9950 25412 9956 25424
rect 8619 25384 9956 25412
rect 8619 25381 8631 25384
rect 8573 25375 8631 25381
rect 9950 25372 9956 25384
rect 10008 25372 10014 25424
rect 14829 25415 14887 25421
rect 14829 25381 14841 25415
rect 14875 25412 14887 25415
rect 14875 25384 15608 25412
rect 14875 25381 14887 25384
rect 14829 25375 14887 25381
rect 8386 25304 8392 25356
rect 8444 25304 8450 25356
rect 12526 25304 12532 25356
rect 12584 25304 12590 25356
rect 15378 25304 15384 25356
rect 15436 25304 15442 25356
rect 15580 25353 15608 25384
rect 16132 25353 16160 25440
rect 16482 25372 16488 25424
rect 16540 25412 16546 25424
rect 18524 25412 18552 25443
rect 18690 25440 18696 25492
rect 18748 25440 18754 25492
rect 18782 25440 18788 25492
rect 18840 25440 18846 25492
rect 21174 25440 21180 25492
rect 21232 25440 21238 25492
rect 21358 25440 21364 25492
rect 21416 25440 21422 25492
rect 22554 25440 22560 25492
rect 22612 25440 22618 25492
rect 23106 25440 23112 25492
rect 23164 25440 23170 25492
rect 24026 25440 24032 25492
rect 24084 25440 24090 25492
rect 27249 25483 27307 25489
rect 27249 25449 27261 25483
rect 27295 25480 27307 25483
rect 27338 25480 27344 25492
rect 27295 25452 27344 25480
rect 27295 25449 27307 25452
rect 27249 25443 27307 25449
rect 27338 25440 27344 25452
rect 27396 25440 27402 25492
rect 27890 25440 27896 25492
rect 27948 25480 27954 25492
rect 28077 25483 28135 25489
rect 28077 25480 28089 25483
rect 27948 25452 28089 25480
rect 27948 25440 27954 25452
rect 28077 25449 28089 25452
rect 28123 25449 28135 25483
rect 28077 25443 28135 25449
rect 28353 25483 28411 25489
rect 28353 25449 28365 25483
rect 28399 25480 28411 25483
rect 28534 25480 28540 25492
rect 28399 25452 28540 25480
rect 28399 25449 28411 25452
rect 28353 25443 28411 25449
rect 28534 25440 28540 25452
rect 28592 25440 28598 25492
rect 16540 25384 18552 25412
rect 16540 25372 16546 25384
rect 15565 25347 15623 25353
rect 15565 25313 15577 25347
rect 15611 25313 15623 25347
rect 15565 25307 15623 25313
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25313 16175 25347
rect 16117 25307 16175 25313
rect 16301 25347 16359 25353
rect 16301 25313 16313 25347
rect 16347 25344 16359 25347
rect 17310 25344 17316 25356
rect 16347 25316 17316 25344
rect 16347 25313 16359 25316
rect 16301 25307 16359 25313
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 18800 25344 18828 25440
rect 18877 25415 18935 25421
rect 18877 25381 18889 25415
rect 18923 25412 18935 25415
rect 18923 25384 19472 25412
rect 18923 25381 18935 25384
rect 18877 25375 18935 25381
rect 19444 25353 19472 25384
rect 19245 25347 19303 25353
rect 19245 25344 19257 25347
rect 17512 25316 18644 25344
rect 18800 25316 19257 25344
rect 7138 25248 7880 25276
rect 7138 25245 7150 25248
rect 7092 25239 7150 25245
rect 8294 25236 8300 25288
rect 8352 25236 8358 25288
rect 5344 25211 5402 25217
rect 5344 25177 5356 25211
rect 5390 25208 5402 25211
rect 6086 25208 6092 25220
rect 5390 25180 6092 25208
rect 5390 25177 5402 25180
rect 5344 25171 5402 25177
rect 6086 25168 6092 25180
rect 6144 25168 6150 25220
rect 8404 25208 8432 25304
rect 17512 25288 17540 25316
rect 8757 25279 8815 25285
rect 8757 25245 8769 25279
rect 8803 25276 8815 25279
rect 8941 25279 8999 25285
rect 8803 25248 8892 25276
rect 8803 25245 8815 25248
rect 8757 25239 8815 25245
rect 8864 25220 8892 25248
rect 8941 25245 8953 25279
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25276 9827 25279
rect 10229 25279 10287 25285
rect 10229 25276 10241 25279
rect 9815 25248 10241 25276
rect 9815 25245 9827 25248
rect 9769 25239 9827 25245
rect 10229 25245 10241 25248
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 6196 25180 8432 25208
rect 6196 25140 6224 25180
rect 8846 25168 8852 25220
rect 8904 25168 8910 25220
rect 5000 25112 6224 25140
rect 6549 25143 6607 25149
rect 6549 25109 6561 25143
rect 6595 25140 6607 25143
rect 7190 25140 7196 25152
rect 6595 25112 7196 25140
rect 6595 25109 6607 25112
rect 6549 25103 6607 25109
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 8205 25143 8263 25149
rect 8205 25109 8217 25143
rect 8251 25140 8263 25143
rect 8294 25140 8300 25152
rect 8251 25112 8300 25140
rect 8251 25109 8263 25112
rect 8205 25103 8263 25109
rect 8294 25100 8300 25112
rect 8352 25140 8358 25152
rect 8956 25140 8984 25239
rect 10244 25208 10272 25239
rect 10318 25236 10324 25288
rect 10376 25236 10382 25288
rect 10588 25279 10646 25285
rect 10588 25245 10600 25279
rect 10634 25276 10646 25279
rect 11146 25276 11152 25288
rect 10634 25248 11152 25276
rect 10634 25245 10646 25248
rect 10588 25239 10646 25245
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 11793 25279 11851 25285
rect 11793 25276 11805 25279
rect 11716 25248 11805 25276
rect 11054 25208 11060 25220
rect 10244 25180 11060 25208
rect 11054 25168 11060 25180
rect 11112 25208 11118 25220
rect 11716 25208 11744 25248
rect 11793 25245 11805 25248
rect 11839 25245 11851 25279
rect 11793 25239 11851 25245
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 12785 25279 12843 25285
rect 12785 25276 12797 25279
rect 12400 25248 12797 25276
rect 12400 25236 12406 25248
rect 12785 25245 12797 25248
rect 12831 25245 12843 25279
rect 12785 25239 12843 25245
rect 14090 25236 14096 25288
rect 14148 25236 14154 25288
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25245 15071 25279
rect 15013 25239 15071 25245
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25276 15163 25279
rect 15194 25276 15200 25288
rect 15151 25248 15200 25276
rect 15151 25245 15163 25248
rect 15105 25239 15163 25245
rect 11112 25180 11744 25208
rect 15028 25208 15056 25239
rect 15194 25236 15200 25248
rect 15252 25276 15258 25288
rect 15252 25248 16344 25276
rect 15252 25236 15258 25248
rect 16316 25220 16344 25248
rect 16942 25236 16948 25288
rect 17000 25236 17006 25288
rect 17494 25236 17500 25288
rect 17552 25272 17558 25288
rect 17552 25244 17593 25272
rect 17552 25236 17558 25244
rect 17678 25236 17684 25288
rect 17736 25276 17742 25288
rect 17773 25279 17831 25285
rect 17773 25276 17785 25279
rect 17736 25248 17785 25276
rect 17736 25236 17742 25248
rect 17773 25245 17785 25248
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 17862 25236 17868 25288
rect 17920 25236 17926 25288
rect 18616 25285 18644 25316
rect 19245 25313 19257 25316
rect 19291 25313 19303 25347
rect 19245 25307 19303 25313
rect 19429 25347 19487 25353
rect 19429 25313 19441 25347
rect 19475 25313 19487 25347
rect 19429 25307 19487 25313
rect 20901 25347 20959 25353
rect 20901 25313 20913 25347
rect 20947 25344 20959 25347
rect 21376 25344 21404 25440
rect 20947 25316 21404 25344
rect 20947 25313 20959 25316
rect 20901 25307 20959 25313
rect 21450 25304 21456 25356
rect 21508 25344 21514 25356
rect 21910 25344 21916 25356
rect 21508 25316 21916 25344
rect 21508 25304 21514 25316
rect 21910 25304 21916 25316
rect 21968 25304 21974 25356
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 19058 25236 19064 25288
rect 19116 25236 19122 25288
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 22002 25236 22008 25288
rect 22060 25236 22066 25288
rect 22572 25276 22600 25440
rect 24044 25344 24072 25440
rect 24489 25347 24547 25353
rect 24489 25344 24501 25347
rect 24044 25316 24501 25344
rect 24489 25313 24501 25316
rect 24535 25313 24547 25347
rect 24489 25307 24547 25313
rect 25866 25304 25872 25356
rect 25924 25304 25930 25356
rect 27356 25353 27384 25440
rect 27982 25372 27988 25424
rect 28040 25372 28046 25424
rect 27341 25347 27399 25353
rect 27341 25313 27353 25347
rect 27387 25313 27399 25347
rect 27341 25307 27399 25313
rect 28166 25304 28172 25356
rect 28224 25344 28230 25356
rect 28224 25316 28580 25344
rect 28224 25304 28230 25316
rect 22741 25279 22799 25285
rect 22741 25276 22753 25279
rect 22572 25248 22753 25276
rect 22741 25245 22753 25248
rect 22787 25245 22799 25279
rect 22741 25239 22799 25245
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25276 23075 25279
rect 23106 25276 23112 25288
rect 23063 25248 23112 25276
rect 23063 25245 23075 25248
rect 23017 25239 23075 25245
rect 23106 25236 23112 25248
rect 23164 25276 23170 25288
rect 23382 25276 23388 25288
rect 23164 25248 23388 25276
rect 23164 25236 23170 25248
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 15028 25180 15332 25208
rect 11112 25168 11118 25180
rect 8352 25112 8984 25140
rect 8352 25100 8358 25112
rect 9582 25100 9588 25152
rect 9640 25100 9646 25152
rect 10042 25100 10048 25152
rect 10100 25100 10106 25152
rect 11716 25149 11744 25180
rect 11701 25143 11759 25149
rect 11701 25109 11713 25143
rect 11747 25109 11759 25143
rect 11701 25103 11759 25109
rect 12434 25100 12440 25152
rect 12492 25100 12498 25152
rect 14734 25100 14740 25152
rect 14792 25100 14798 25152
rect 15194 25100 15200 25152
rect 15252 25100 15258 25152
rect 15304 25140 15332 25180
rect 16298 25168 16304 25220
rect 16356 25208 16362 25220
rect 16960 25208 16988 25236
rect 17497 25235 17555 25236
rect 16356 25180 16988 25208
rect 22020 25208 22048 25236
rect 22020 25180 22600 25208
rect 16356 25168 16362 25180
rect 15654 25140 15660 25152
rect 15304 25112 15660 25140
rect 15654 25100 15660 25112
rect 15712 25100 15718 25152
rect 16025 25143 16083 25149
rect 16025 25109 16037 25143
rect 16071 25140 16083 25143
rect 16758 25140 16764 25152
rect 16071 25112 16764 25140
rect 16071 25109 16083 25112
rect 16025 25103 16083 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17313 25143 17371 25149
rect 17313 25109 17325 25143
rect 17359 25140 17371 25143
rect 17678 25140 17684 25152
rect 17359 25112 17684 25140
rect 17359 25109 17371 25112
rect 17313 25103 17371 25109
rect 17678 25100 17684 25112
rect 17736 25100 17742 25152
rect 19702 25100 19708 25152
rect 19760 25140 19766 25152
rect 19889 25143 19947 25149
rect 19889 25140 19901 25143
rect 19760 25112 19901 25140
rect 19760 25100 19766 25112
rect 19889 25109 19901 25112
rect 19935 25109 19947 25143
rect 19889 25103 19947 25109
rect 22186 25100 22192 25152
rect 22244 25140 22250 25152
rect 22572 25149 22600 25180
rect 24578 25168 24584 25220
rect 24636 25168 24642 25220
rect 24854 25168 24860 25220
rect 24912 25208 24918 25220
rect 25501 25211 25559 25217
rect 25501 25208 25513 25211
rect 24912 25180 25513 25208
rect 24912 25168 24918 25180
rect 25501 25177 25513 25180
rect 25547 25177 25559 25211
rect 25501 25171 25559 25177
rect 25792 25152 25820 25239
rect 25958 25236 25964 25288
rect 26016 25276 26022 25288
rect 26053 25279 26111 25285
rect 26053 25276 26065 25279
rect 26016 25248 26065 25276
rect 26016 25236 26022 25248
rect 26053 25245 26065 25248
rect 26099 25245 26111 25279
rect 26605 25279 26663 25285
rect 26605 25276 26617 25279
rect 26053 25239 26111 25245
rect 26528 25248 26617 25276
rect 22465 25143 22523 25149
rect 22465 25140 22477 25143
rect 22244 25112 22477 25140
rect 22244 25100 22250 25112
rect 22465 25109 22477 25112
rect 22511 25109 22523 25143
rect 22465 25103 22523 25109
rect 22557 25143 22615 25149
rect 22557 25109 22569 25143
rect 22603 25109 22615 25143
rect 22557 25103 22615 25109
rect 24026 25100 24032 25152
rect 24084 25100 24090 25152
rect 25590 25100 25596 25152
rect 25648 25100 25654 25152
rect 25774 25100 25780 25152
rect 25832 25100 25838 25152
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26528 25149 26556 25248
rect 26605 25245 26617 25248
rect 26651 25245 26663 25279
rect 26605 25239 26663 25245
rect 26786 25236 26792 25288
rect 26844 25236 26850 25288
rect 27522 25236 27528 25288
rect 27580 25236 27586 25288
rect 28552 25285 28580 25316
rect 28261 25279 28319 25285
rect 28261 25245 28273 25279
rect 28307 25245 28319 25279
rect 28261 25239 28319 25245
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25245 28595 25279
rect 28537 25239 28595 25245
rect 27154 25168 27160 25220
rect 27212 25208 27218 25220
rect 28276 25208 28304 25239
rect 27212 25180 28304 25208
rect 27212 25168 27218 25180
rect 26513 25143 26571 25149
rect 26513 25140 26525 25143
rect 26292 25112 26525 25140
rect 26292 25100 26298 25112
rect 26513 25109 26525 25112
rect 26559 25109 26571 25143
rect 26513 25103 26571 25109
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 4522 24896 4528 24948
rect 4580 24936 4586 24948
rect 7650 24936 7656 24948
rect 4580 24908 7656 24936
rect 4580 24896 4586 24908
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 7742 24896 7748 24948
rect 7800 24896 7806 24948
rect 10042 24896 10048 24948
rect 10100 24936 10106 24948
rect 10100 24908 10824 24936
rect 10100 24896 10106 24908
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 6641 24871 6699 24877
rect 2832 24840 3280 24868
rect 2832 24828 2838 24840
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 2041 24803 2099 24809
rect 1627 24772 1900 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 1872 24673 1900 24772
rect 2041 24769 2053 24803
rect 2087 24769 2099 24803
rect 2041 24763 2099 24769
rect 1857 24667 1915 24673
rect 1857 24633 1869 24667
rect 1903 24633 1915 24667
rect 1857 24627 1915 24633
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24596 1731 24599
rect 1762 24596 1768 24608
rect 1719 24568 1768 24596
rect 1719 24565 1731 24568
rect 1673 24559 1731 24565
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 2056 24596 2084 24763
rect 2498 24760 2504 24812
rect 2556 24760 2562 24812
rect 2961 24803 3019 24809
rect 2961 24800 2973 24803
rect 2746 24772 2973 24800
rect 2746 24732 2774 24772
rect 2961 24769 2973 24772
rect 3007 24769 3019 24803
rect 2961 24763 3019 24769
rect 3050 24760 3056 24812
rect 3108 24760 3114 24812
rect 3252 24809 3280 24840
rect 6641 24837 6653 24871
rect 6687 24868 6699 24871
rect 7282 24868 7288 24880
rect 6687 24840 7288 24868
rect 6687 24837 6699 24840
rect 6641 24831 6699 24837
rect 7282 24828 7288 24840
rect 7340 24828 7346 24880
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24769 3295 24803
rect 3237 24763 3295 24769
rect 3786 24760 3792 24812
rect 3844 24760 3850 24812
rect 4332 24803 4390 24809
rect 4332 24769 4344 24803
rect 4378 24800 4390 24803
rect 5810 24800 5816 24812
rect 4378 24772 5816 24800
rect 4378 24769 4390 24772
rect 4332 24763 4390 24769
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24800 7435 24803
rect 7760 24800 7788 24896
rect 10318 24868 10324 24880
rect 9232 24840 10324 24868
rect 7423 24772 7788 24800
rect 7837 24803 7895 24809
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 7837 24769 7849 24803
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 2332 24704 2774 24732
rect 2332 24673 2360 24704
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 4065 24735 4123 24741
rect 4065 24732 4077 24735
rect 3936 24704 4077 24732
rect 3936 24692 3942 24704
rect 4065 24701 4077 24704
rect 4111 24701 4123 24735
rect 4065 24695 4123 24701
rect 5534 24692 5540 24744
rect 5592 24692 5598 24744
rect 5718 24692 5724 24744
rect 5776 24692 5782 24744
rect 6546 24692 6552 24744
rect 6604 24692 6610 24744
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7392 24732 7420 24763
rect 7340 24704 7420 24732
rect 7340 24692 7346 24704
rect 7558 24692 7564 24744
rect 7616 24732 7622 24744
rect 7852 24732 7880 24763
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8754 24800 8760 24812
rect 8352 24772 8760 24800
rect 8352 24760 8358 24772
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 9033 24803 9091 24809
rect 9033 24769 9045 24803
rect 9079 24800 9091 24803
rect 9232 24800 9260 24840
rect 10318 24828 10324 24840
rect 10376 24868 10382 24880
rect 10686 24868 10692 24880
rect 10376 24840 10692 24868
rect 10376 24828 10382 24840
rect 10686 24828 10692 24840
rect 10744 24828 10750 24880
rect 9079 24772 9260 24800
rect 9300 24803 9358 24809
rect 9079 24769 9091 24772
rect 9033 24763 9091 24769
rect 9300 24769 9312 24803
rect 9346 24800 9358 24803
rect 9582 24800 9588 24812
rect 9346 24772 9588 24800
rect 9346 24769 9358 24772
rect 9300 24763 9358 24769
rect 9582 24760 9588 24772
rect 9640 24760 9646 24812
rect 10796 24809 10824 24908
rect 11054 24896 11060 24948
rect 11112 24896 11118 24948
rect 14182 24896 14188 24948
rect 14240 24936 14246 24948
rect 14277 24939 14335 24945
rect 14277 24936 14289 24939
rect 14240 24908 14289 24936
rect 14240 24896 14246 24908
rect 14277 24905 14289 24908
rect 14323 24905 14335 24939
rect 14277 24899 14335 24905
rect 14734 24896 14740 24948
rect 14792 24896 14798 24948
rect 15470 24896 15476 24948
rect 15528 24896 15534 24948
rect 15654 24896 15660 24948
rect 15712 24936 15718 24948
rect 16117 24939 16175 24945
rect 16117 24936 16129 24939
rect 15712 24908 16129 24936
rect 15712 24896 15718 24908
rect 16117 24905 16129 24908
rect 16163 24905 16175 24939
rect 17862 24936 17868 24948
rect 16117 24899 16175 24905
rect 17052 24908 17868 24936
rect 11072 24868 11100 24896
rect 12710 24868 12716 24880
rect 10888 24840 11100 24868
rect 12452 24840 12716 24868
rect 10888 24809 10916 24840
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10873 24803 10931 24809
rect 10873 24769 10885 24803
rect 10919 24769 10931 24803
rect 10873 24763 10931 24769
rect 11333 24803 11391 24809
rect 11333 24769 11345 24803
rect 11379 24800 11391 24803
rect 11609 24803 11667 24809
rect 11609 24800 11621 24803
rect 11379 24772 11621 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 11609 24769 11621 24772
rect 11655 24800 11667 24803
rect 11882 24800 11888 24812
rect 11655 24772 11888 24800
rect 11655 24769 11667 24772
rect 11609 24763 11667 24769
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 12069 24803 12127 24809
rect 12069 24769 12081 24803
rect 12115 24800 12127 24803
rect 12452 24800 12480 24840
rect 12710 24828 12716 24840
rect 12768 24828 12774 24880
rect 12115 24772 12480 24800
rect 13164 24803 13222 24809
rect 12115 24769 12127 24772
rect 12069 24763 12127 24769
rect 13164 24769 13176 24803
rect 13210 24800 13222 24803
rect 14752 24800 14780 24896
rect 15194 24800 15200 24812
rect 13210 24772 14780 24800
rect 14844 24772 15200 24800
rect 13210 24769 13222 24772
rect 13164 24763 13222 24769
rect 7616 24704 7880 24732
rect 7616 24692 7622 24704
rect 8570 24692 8576 24744
rect 8628 24692 8634 24744
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11698 24732 11704 24744
rect 11011 24704 11704 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 11698 24692 11704 24704
rect 11756 24692 11762 24744
rect 12158 24692 12164 24744
rect 12216 24692 12222 24744
rect 12250 24692 12256 24744
rect 12308 24732 12314 24744
rect 12526 24732 12532 24744
rect 12308 24704 12532 24732
rect 12308 24692 12314 24704
rect 12526 24692 12532 24704
rect 12584 24732 12590 24744
rect 12897 24735 12955 24741
rect 12897 24732 12909 24735
rect 12584 24704 12909 24732
rect 12584 24692 12590 24704
rect 12897 24701 12909 24704
rect 12943 24701 12955 24735
rect 12897 24695 12955 24701
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 14844 24732 14872 24772
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15488 24800 15516 24896
rect 17052 24868 17080 24908
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 18693 24939 18751 24945
rect 18693 24905 18705 24939
rect 18739 24936 18751 24939
rect 19058 24936 19064 24948
rect 18739 24908 19064 24936
rect 18739 24905 18751 24908
rect 18693 24899 18751 24905
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 20714 24896 20720 24948
rect 20772 24936 20778 24948
rect 24210 24936 24216 24948
rect 20772 24908 24216 24936
rect 20772 24896 20778 24908
rect 24210 24896 24216 24908
rect 24268 24936 24274 24948
rect 26329 24939 26387 24945
rect 24268 24908 24808 24936
rect 24268 24896 24274 24908
rect 16868 24840 17080 24868
rect 15841 24803 15899 24809
rect 15841 24800 15853 24803
rect 15488 24772 15853 24800
rect 15841 24769 15853 24772
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 16022 24760 16028 24812
rect 16080 24800 16086 24812
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 16080 24772 16313 24800
rect 16080 24760 16086 24772
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 16758 24760 16764 24812
rect 16816 24760 16822 24812
rect 16868 24809 16896 24840
rect 17218 24828 17224 24880
rect 17276 24828 17282 24880
rect 21082 24868 21088 24880
rect 20548 24840 21088 24868
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 17236 24800 17264 24828
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 17236 24772 17509 24800
rect 16853 24763 16911 24769
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24800 18475 24803
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 18463 24772 18889 24800
rect 18463 24769 18475 24772
rect 18417 24763 18475 24769
rect 18877 24769 18889 24772
rect 18923 24800 18935 24803
rect 19705 24803 19763 24809
rect 18923 24772 19656 24800
rect 18923 24769 18935 24772
rect 18877 24763 18935 24769
rect 14599 24704 14872 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 2317 24667 2375 24673
rect 2317 24633 2329 24667
rect 2363 24633 2375 24667
rect 3050 24664 3056 24676
rect 2317 24627 2375 24633
rect 2700 24636 3056 24664
rect 2700 24596 2728 24636
rect 3050 24624 3056 24636
rect 3108 24624 3114 24676
rect 7006 24624 7012 24676
rect 7064 24664 7070 24676
rect 7101 24667 7159 24673
rect 7101 24664 7113 24667
rect 7064 24636 7113 24664
rect 7064 24624 7070 24636
rect 7101 24633 7113 24636
rect 7147 24633 7159 24667
rect 7101 24627 7159 24633
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 14384 24664 14412 24695
rect 14918 24692 14924 24744
rect 14976 24732 14982 24744
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 14976 24704 15117 24732
rect 14976 24692 14982 24704
rect 15105 24701 15117 24704
rect 15151 24701 15163 24735
rect 16776 24732 16804 24760
rect 17681 24735 17739 24741
rect 17681 24732 17693 24735
rect 16776 24704 17693 24732
rect 15105 24695 15163 24701
rect 17681 24701 17693 24704
rect 17727 24701 17739 24735
rect 17681 24695 17739 24701
rect 17865 24735 17923 24741
rect 17865 24701 17877 24735
rect 17911 24732 17923 24735
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 17911 24704 18521 24732
rect 17911 24701 17923 24704
rect 17865 24695 17923 24701
rect 18509 24701 18521 24704
rect 18555 24701 18567 24735
rect 18509 24695 18567 24701
rect 15933 24667 15991 24673
rect 15933 24664 15945 24667
rect 11931 24636 12940 24664
rect 14384 24636 15945 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 2056 24568 2728 24596
rect 2774 24556 2780 24608
rect 2832 24556 2838 24608
rect 3694 24556 3700 24608
rect 3752 24556 3758 24608
rect 3881 24599 3939 24605
rect 3881 24565 3893 24599
rect 3927 24596 3939 24599
rect 3970 24596 3976 24608
rect 3927 24568 3976 24596
rect 3927 24565 3939 24568
rect 3881 24559 3939 24565
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4798 24556 4804 24608
rect 4856 24596 4862 24608
rect 5166 24596 5172 24608
rect 4856 24568 5172 24596
rect 4856 24556 4862 24568
rect 5166 24556 5172 24568
rect 5224 24596 5230 24608
rect 5445 24599 5503 24605
rect 5445 24596 5457 24599
rect 5224 24568 5457 24596
rect 5224 24556 5230 24568
rect 5445 24565 5457 24568
rect 5491 24565 5503 24599
rect 5445 24559 5503 24565
rect 6086 24556 6092 24608
rect 6144 24556 6150 24608
rect 7466 24556 7472 24608
rect 7524 24556 7530 24608
rect 7929 24599 7987 24605
rect 7929 24565 7941 24599
rect 7975 24596 7987 24599
rect 8294 24596 8300 24608
rect 7975 24568 8300 24596
rect 7975 24565 7987 24568
rect 7929 24559 7987 24565
rect 8294 24556 8300 24568
rect 8352 24556 8358 24608
rect 10410 24556 10416 24608
rect 10468 24556 10474 24608
rect 10597 24599 10655 24605
rect 10597 24565 10609 24599
rect 10643 24596 10655 24599
rect 10870 24596 10876 24608
rect 10643 24568 10876 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 11238 24596 11244 24608
rect 11195 24568 11244 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 11790 24596 11796 24608
rect 11747 24568 11796 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 12802 24556 12808 24608
rect 12860 24556 12866 24608
rect 12912 24596 12940 24636
rect 15933 24633 15945 24636
rect 15979 24633 15991 24667
rect 15933 24627 15991 24633
rect 17313 24667 17371 24673
rect 17313 24633 17325 24667
rect 17359 24664 17371 24667
rect 17586 24664 17592 24676
rect 17359 24636 17592 24664
rect 17359 24633 17371 24636
rect 17313 24627 17371 24633
rect 17586 24624 17592 24636
rect 17644 24624 17650 24676
rect 19628 24608 19656 24772
rect 19705 24769 19717 24803
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 20340 24803 20398 24809
rect 20340 24769 20352 24803
rect 20386 24800 20398 24803
rect 20548 24800 20576 24840
rect 21082 24828 21088 24840
rect 21140 24828 21146 24880
rect 23560 24871 23618 24877
rect 22020 24840 22324 24868
rect 20386 24772 20576 24800
rect 20386 24769 20398 24772
rect 20340 24763 20398 24769
rect 19720 24664 19748 24763
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 20680 24772 21833 24800
rect 20680 24760 20686 24772
rect 21821 24769 21833 24772
rect 21867 24800 21879 24803
rect 22020 24800 22048 24840
rect 22094 24809 22100 24812
rect 21867 24772 22048 24800
rect 21867 24769 21879 24772
rect 21821 24763 21879 24769
rect 22088 24763 22100 24809
rect 22152 24800 22158 24812
rect 22296 24800 22324 24840
rect 23560 24837 23572 24871
rect 23606 24868 23618 24871
rect 24026 24868 24032 24880
rect 23606 24840 24032 24868
rect 23606 24837 23618 24840
rect 23560 24831 23618 24837
rect 24026 24828 24032 24840
rect 24084 24828 24090 24880
rect 24780 24868 24808 24908
rect 26329 24905 26341 24939
rect 26375 24936 26387 24939
rect 26510 24936 26516 24948
rect 26375 24908 26516 24936
rect 26375 24905 26387 24908
rect 26329 24899 26387 24905
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 26605 24939 26663 24945
rect 26605 24905 26617 24939
rect 26651 24936 26663 24939
rect 26786 24936 26792 24948
rect 26651 24908 26792 24936
rect 26651 24905 26663 24908
rect 26605 24899 26663 24905
rect 26786 24896 26792 24908
rect 26844 24896 26850 24948
rect 28166 24896 28172 24948
rect 28224 24896 28230 24948
rect 27154 24868 27160 24880
rect 24780 24840 25268 24868
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 22152 24772 22188 24800
rect 22296 24772 23305 24800
rect 22094 24760 22100 24763
rect 22152 24760 22158 24772
rect 23293 24769 23305 24772
rect 23339 24769 23351 24803
rect 24854 24800 24860 24812
rect 23293 24763 23351 24769
rect 24504 24772 24860 24800
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 20073 24735 20131 24741
rect 20073 24732 20085 24735
rect 19852 24704 20085 24732
rect 19852 24692 19858 24704
rect 20073 24701 20085 24704
rect 20119 24701 20131 24735
rect 20073 24695 20131 24701
rect 21450 24692 21456 24744
rect 21508 24692 21514 24744
rect 19720 24636 20116 24664
rect 20088 24608 20116 24636
rect 13538 24596 13544 24608
rect 12912 24568 13544 24596
rect 13538 24556 13544 24568
rect 13596 24556 13602 24608
rect 15013 24599 15071 24605
rect 15013 24565 15025 24599
rect 15059 24596 15071 24599
rect 15378 24596 15384 24608
rect 15059 24568 15384 24596
rect 15059 24565 15071 24568
rect 15013 24559 15071 24565
rect 15378 24556 15384 24568
rect 15436 24596 15442 24608
rect 15473 24599 15531 24605
rect 15473 24596 15485 24599
rect 15436 24568 15485 24596
rect 15436 24556 15442 24568
rect 15473 24565 15485 24568
rect 15519 24565 15531 24599
rect 15473 24559 15531 24565
rect 16942 24556 16948 24608
rect 17000 24556 17006 24608
rect 18230 24556 18236 24608
rect 18288 24556 18294 24608
rect 19518 24556 19524 24608
rect 19576 24556 19582 24608
rect 19610 24556 19616 24608
rect 19668 24556 19674 24608
rect 20070 24556 20076 24608
rect 20128 24556 20134 24608
rect 21468 24605 21496 24692
rect 21453 24599 21511 24605
rect 21453 24565 21465 24599
rect 21499 24596 21511 24599
rect 22462 24596 22468 24608
rect 21499 24568 22468 24596
rect 21499 24565 21511 24568
rect 21453 24559 21511 24565
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 23164 24568 23213 24596
rect 23164 24556 23170 24568
rect 23201 24565 23213 24568
rect 23247 24565 23259 24599
rect 23308 24596 23336 24763
rect 23474 24596 23480 24608
rect 23308 24568 23480 24596
rect 23201 24559 23259 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 24504 24596 24532 24772
rect 24854 24760 24860 24772
rect 24912 24800 24918 24812
rect 25130 24800 25136 24812
rect 24912 24772 25136 24800
rect 24912 24760 24918 24772
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 25240 24800 25268 24840
rect 26252 24840 27160 24868
rect 25501 24803 25559 24809
rect 25501 24800 25513 24803
rect 25240 24772 25513 24800
rect 25501 24769 25513 24772
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 26050 24760 26056 24812
rect 26108 24800 26114 24812
rect 26252 24809 26280 24840
rect 26237 24803 26295 24809
rect 26237 24800 26249 24803
rect 26108 24772 26249 24800
rect 26108 24760 26114 24772
rect 26237 24769 26249 24772
rect 26283 24769 26295 24803
rect 26237 24763 26295 24769
rect 26510 24760 26516 24812
rect 26568 24800 26574 24812
rect 26988 24809 27016 24840
rect 27154 24828 27160 24840
rect 27212 24828 27218 24880
rect 26789 24803 26847 24809
rect 26789 24800 26801 24803
rect 26568 24772 26801 24800
rect 26568 24760 26574 24772
rect 26789 24769 26801 24772
rect 26835 24769 26847 24803
rect 26789 24763 26847 24769
rect 26973 24803 27031 24809
rect 26973 24769 26985 24803
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27062 24760 27068 24812
rect 27120 24760 27126 24812
rect 28077 24803 28135 24809
rect 28077 24769 28089 24803
rect 28123 24800 28135 24803
rect 28184 24800 28212 24896
rect 28350 24800 28356 24812
rect 28123 24772 28356 24800
rect 28123 24769 28135 24772
rect 28077 24763 28135 24769
rect 28350 24760 28356 24772
rect 28408 24760 28414 24812
rect 28537 24803 28595 24809
rect 28537 24769 28549 24803
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 24765 24735 24823 24741
rect 24765 24732 24777 24735
rect 24688 24704 24777 24732
rect 24688 24676 24716 24704
rect 24765 24701 24777 24704
rect 24811 24701 24823 24735
rect 24765 24695 24823 24701
rect 25682 24692 25688 24744
rect 25740 24692 25746 24744
rect 27154 24692 27160 24744
rect 27212 24732 27218 24744
rect 27341 24735 27399 24741
rect 27341 24732 27353 24735
rect 27212 24704 27353 24732
rect 27212 24692 27218 24704
rect 27341 24701 27353 24704
rect 27387 24732 27399 24735
rect 28552 24732 28580 24763
rect 27387 24704 28580 24732
rect 27387 24701 27399 24704
rect 27341 24695 27399 24701
rect 24670 24624 24676 24676
rect 24728 24624 24734 24676
rect 26145 24667 26203 24673
rect 26145 24633 26157 24667
rect 26191 24664 26203 24667
rect 26234 24664 26240 24676
rect 26191 24636 26240 24664
rect 26191 24633 26203 24636
rect 26145 24627 26203 24633
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 28258 24624 28264 24676
rect 28316 24624 28322 24676
rect 23624 24568 24532 24596
rect 23624 24556 23630 24568
rect 24578 24556 24584 24608
rect 24636 24596 24642 24608
rect 25409 24599 25467 24605
rect 25409 24596 25421 24599
rect 24636 24568 25421 24596
rect 24636 24556 24642 24568
rect 25409 24565 25421 24568
rect 25455 24565 25467 24599
rect 25409 24559 25467 24565
rect 27982 24556 27988 24608
rect 28040 24556 28046 24608
rect 28166 24556 28172 24608
rect 28224 24556 28230 24608
rect 28276 24596 28304 24624
rect 28353 24599 28411 24605
rect 28353 24596 28365 24599
rect 28276 24568 28365 24596
rect 28353 24565 28365 24568
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 1762 24352 1768 24404
rect 1820 24392 1826 24404
rect 2777 24395 2835 24401
rect 1820 24364 2728 24392
rect 1820 24352 1826 24364
rect 1394 24148 1400 24200
rect 1452 24148 1458 24200
rect 1664 24123 1722 24129
rect 1664 24089 1676 24123
rect 1710 24120 1722 24123
rect 2130 24120 2136 24132
rect 1710 24092 2136 24120
rect 1710 24089 1722 24092
rect 1664 24083 1722 24089
rect 2130 24080 2136 24092
rect 2188 24080 2194 24132
rect 2700 24120 2728 24364
rect 2777 24361 2789 24395
rect 2823 24392 2835 24395
rect 2866 24392 2872 24404
rect 2823 24364 2872 24392
rect 2823 24361 2835 24364
rect 2777 24355 2835 24361
rect 2866 24352 2872 24364
rect 2924 24352 2930 24404
rect 4525 24395 4583 24401
rect 4525 24361 4537 24395
rect 4571 24392 4583 24395
rect 5718 24392 5724 24404
rect 4571 24364 5724 24392
rect 4571 24361 4583 24364
rect 4525 24355 4583 24361
rect 5718 24352 5724 24364
rect 5776 24352 5782 24404
rect 5810 24352 5816 24404
rect 5868 24392 5874 24404
rect 6089 24395 6147 24401
rect 6089 24392 6101 24395
rect 5868 24364 6101 24392
rect 5868 24352 5874 24364
rect 6089 24361 6101 24364
rect 6135 24361 6147 24395
rect 6089 24355 6147 24361
rect 6546 24352 6552 24404
rect 6604 24352 6610 24404
rect 6638 24352 6644 24404
rect 6696 24392 6702 24404
rect 6696 24364 8248 24392
rect 6696 24352 6702 24364
rect 2884 24265 2912 24352
rect 3694 24284 3700 24336
rect 3752 24324 3758 24336
rect 4157 24327 4215 24333
rect 4157 24324 4169 24327
rect 3752 24296 4169 24324
rect 3752 24284 3758 24296
rect 4157 24293 4169 24296
rect 4203 24293 4215 24327
rect 7282 24324 7288 24336
rect 4157 24287 4215 24293
rect 5552 24296 7288 24324
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24225 2927 24259
rect 2869 24219 2927 24225
rect 2958 24216 2964 24268
rect 3016 24216 3022 24268
rect 3234 24216 3240 24268
rect 3292 24256 3298 24268
rect 3973 24259 4031 24265
rect 3973 24256 3985 24259
rect 3292 24228 3985 24256
rect 3292 24216 3298 24228
rect 3973 24225 3985 24228
rect 4019 24225 4031 24259
rect 4890 24256 4896 24268
rect 3973 24219 4031 24225
rect 4816 24228 4896 24256
rect 2976 24188 3004 24216
rect 3789 24191 3847 24197
rect 3789 24188 3801 24191
rect 2976 24160 3801 24188
rect 3789 24157 3801 24160
rect 3835 24157 3847 24191
rect 3789 24151 3847 24157
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 4816 24197 4844 24228
rect 4890 24216 4896 24228
rect 4948 24256 4954 24268
rect 5552 24265 5580 24296
rect 7282 24284 7288 24296
rect 7340 24284 7346 24336
rect 8021 24327 8079 24333
rect 8021 24293 8033 24327
rect 8067 24293 8079 24327
rect 8021 24287 8079 24293
rect 5537 24259 5595 24265
rect 5537 24256 5549 24259
rect 4948 24228 5549 24256
rect 4948 24216 4954 24228
rect 5537 24225 5549 24228
rect 5583 24225 5595 24259
rect 5537 24219 5595 24225
rect 6365 24259 6423 24265
rect 6365 24225 6377 24259
rect 6411 24256 6423 24259
rect 6822 24256 6828 24268
rect 6411 24228 6828 24256
rect 6411 24225 6423 24228
rect 6365 24219 6423 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 8036 24256 8064 24287
rect 7668 24228 8064 24256
rect 4709 24191 4767 24197
rect 4709 24188 4721 24191
rect 4304 24160 4721 24188
rect 4304 24148 4310 24160
rect 4709 24157 4721 24160
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 5166 24148 5172 24200
rect 5224 24148 5230 24200
rect 6181 24191 6239 24197
rect 6181 24157 6193 24191
rect 6227 24188 6239 24191
rect 6914 24188 6920 24200
rect 6227 24160 6920 24188
rect 6227 24157 6239 24160
rect 6181 24151 6239 24157
rect 6914 24148 6920 24160
rect 6972 24148 6978 24200
rect 7668 24197 7696 24228
rect 8220 24197 8248 24364
rect 10686 24352 10692 24404
rect 10744 24392 10750 24404
rect 11514 24392 11520 24404
rect 10744 24364 11520 24392
rect 10744 24352 10750 24364
rect 8846 24324 8852 24336
rect 8312 24296 8852 24324
rect 8312 24197 8340 24296
rect 8846 24284 8852 24296
rect 8904 24324 8910 24336
rect 9214 24324 9220 24336
rect 8904 24296 9220 24324
rect 8904 24284 8910 24296
rect 9214 24284 9220 24296
rect 9272 24284 9278 24336
rect 11164 24265 11192 24364
rect 11514 24352 11520 24364
rect 11572 24352 11578 24404
rect 11882 24352 11888 24404
rect 11940 24392 11946 24404
rect 11940 24364 12112 24392
rect 11940 24352 11946 24364
rect 12084 24324 12112 24364
rect 12158 24352 12164 24404
rect 12216 24392 12222 24404
rect 13998 24392 14004 24404
rect 12216 24364 14004 24392
rect 12216 24352 12222 24364
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 16942 24352 16948 24404
rect 17000 24352 17006 24404
rect 18230 24352 18236 24404
rect 18288 24352 18294 24404
rect 19518 24352 19524 24404
rect 19576 24352 19582 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 23566 24392 23572 24404
rect 19668 24364 23572 24392
rect 19668 24352 19674 24364
rect 23566 24352 23572 24364
rect 23624 24352 23630 24404
rect 23937 24395 23995 24401
rect 23937 24361 23949 24395
rect 23983 24392 23995 24395
rect 24394 24392 24400 24404
rect 23983 24364 24400 24392
rect 23983 24361 23995 24364
rect 23937 24355 23995 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 24670 24352 24676 24404
rect 24728 24352 24734 24404
rect 25501 24395 25559 24401
rect 25501 24361 25513 24395
rect 25547 24392 25559 24395
rect 25682 24392 25688 24404
rect 25547 24364 25688 24392
rect 25547 24361 25559 24364
rect 25501 24355 25559 24361
rect 25682 24352 25688 24364
rect 25740 24352 25746 24404
rect 25958 24352 25964 24404
rect 26016 24352 26022 24404
rect 27522 24352 27528 24404
rect 27580 24352 27586 24404
rect 12529 24327 12587 24333
rect 12529 24324 12541 24327
rect 12084 24296 12541 24324
rect 12529 24293 12541 24296
rect 12575 24324 12587 24327
rect 12575 24296 12664 24324
rect 12575 24293 12587 24296
rect 12529 24287 12587 24293
rect 12636 24265 12664 24296
rect 14734 24284 14740 24336
rect 14792 24324 14798 24336
rect 15010 24324 15016 24336
rect 14792 24296 15016 24324
rect 14792 24284 14798 24296
rect 15010 24284 15016 24296
rect 15068 24284 15074 24336
rect 16117 24327 16175 24333
rect 16117 24293 16129 24327
rect 16163 24293 16175 24327
rect 16117 24287 16175 24293
rect 16485 24327 16543 24333
rect 16485 24293 16497 24327
rect 16531 24324 16543 24327
rect 16531 24296 16887 24324
rect 16531 24293 16543 24296
rect 16485 24287 16543 24293
rect 8665 24259 8723 24265
rect 8665 24225 8677 24259
rect 8711 24256 8723 24259
rect 9769 24259 9827 24265
rect 9769 24256 9781 24259
rect 8711 24228 9781 24256
rect 8711 24225 8723 24228
rect 8665 24219 8723 24225
rect 9769 24225 9781 24228
rect 9815 24225 9827 24259
rect 9769 24219 9827 24225
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24225 11207 24259
rect 11149 24219 11207 24225
rect 12621 24259 12679 24265
rect 12621 24225 12633 24259
rect 12667 24225 12679 24259
rect 16132 24256 16160 24287
rect 12621 24219 12679 24225
rect 13280 24228 15332 24256
rect 16132 24228 16712 24256
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24157 7711 24191
rect 7653 24151 7711 24157
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 8205 24191 8263 24197
rect 8205 24157 8217 24191
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 8297 24191 8355 24197
rect 8297 24157 8309 24191
rect 8343 24157 8355 24191
rect 8297 24151 8355 24157
rect 5261 24123 5319 24129
rect 2700 24092 4844 24120
rect 4816 24064 4844 24092
rect 5261 24089 5273 24123
rect 5307 24120 5319 24123
rect 6270 24120 6276 24132
rect 5307 24092 6276 24120
rect 5307 24089 5319 24092
rect 5261 24083 5319 24089
rect 6270 24080 6276 24092
rect 6328 24080 6334 24132
rect 7300 24120 7328 24151
rect 6380 24092 7328 24120
rect 3510 24012 3516 24064
rect 3568 24012 3574 24064
rect 4798 24012 4804 24064
rect 4856 24012 4862 24064
rect 4890 24012 4896 24064
rect 4948 24012 4954 24064
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 6380 24052 6408 24092
rect 5132 24024 6408 24052
rect 5132 24012 5138 24024
rect 7098 24012 7104 24064
rect 7156 24012 7162 24064
rect 7469 24055 7527 24061
rect 7469 24021 7481 24055
rect 7515 24052 7527 24055
rect 7650 24052 7656 24064
rect 7515 24024 7656 24052
rect 7515 24021 7527 24024
rect 7469 24015 7527 24021
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 7742 24012 7748 24064
rect 7800 24012 7806 24064
rect 7944 24052 7972 24151
rect 8570 24148 8576 24200
rect 8628 24148 8634 24200
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 8812 24160 9321 24188
rect 8812 24148 8818 24160
rect 9309 24157 9321 24160
rect 9355 24157 9367 24191
rect 9582 24188 9588 24200
rect 9543 24160 9588 24188
rect 9309 24151 9367 24157
rect 9582 24148 9588 24160
rect 9640 24188 9646 24200
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 9640 24160 10793 24188
rect 9640 24148 9646 24160
rect 10781 24157 10793 24160
rect 10827 24157 10839 24191
rect 10781 24151 10839 24157
rect 11057 24191 11115 24197
rect 11057 24157 11069 24191
rect 11103 24157 11115 24191
rect 11057 24151 11115 24157
rect 8389 24123 8447 24129
rect 8389 24089 8401 24123
rect 8435 24120 8447 24123
rect 10318 24120 10324 24132
rect 8435 24092 10324 24120
rect 8435 24089 8447 24092
rect 8389 24083 8447 24089
rect 10318 24080 10324 24092
rect 10376 24080 10382 24132
rect 10413 24123 10471 24129
rect 10413 24089 10425 24123
rect 10459 24120 10471 24123
rect 10502 24120 10508 24132
rect 10459 24092 10508 24120
rect 10459 24089 10471 24092
rect 10413 24083 10471 24089
rect 10502 24080 10508 24092
rect 10560 24120 10566 24132
rect 11072 24120 11100 24151
rect 11238 24148 11244 24200
rect 11296 24188 11302 24200
rect 11974 24188 11980 24200
rect 11296 24160 11980 24188
rect 11296 24148 11302 24160
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 13280 24188 13308 24228
rect 12800 24160 13308 24188
rect 11146 24120 11152 24132
rect 10560 24092 11008 24120
rect 11072 24092 11152 24120
rect 10560 24080 10566 24092
rect 8754 24052 8760 24064
rect 7944 24024 8760 24052
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 9125 24055 9183 24061
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 9306 24052 9312 24064
rect 9171 24024 9312 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 10226 24012 10232 24064
rect 10284 24012 10290 24064
rect 10870 24012 10876 24064
rect 10928 24012 10934 24064
rect 10980 24052 11008 24092
rect 11146 24080 11152 24092
rect 11204 24080 11210 24132
rect 11416 24123 11474 24129
rect 11416 24089 11428 24123
rect 11462 24120 11474 24123
rect 12434 24120 12440 24132
rect 11462 24092 12440 24120
rect 11462 24089 11474 24092
rect 11416 24083 11474 24089
rect 12434 24080 12440 24092
rect 12492 24080 12498 24132
rect 12800 24052 12828 24160
rect 13538 24148 13544 24200
rect 13596 24148 13602 24200
rect 13906 24148 13912 24200
rect 13964 24148 13970 24200
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 14056 24160 14105 24188
rect 14056 24148 14062 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 13541 24133 13553 24148
rect 13587 24133 13599 24148
rect 13541 24127 13599 24133
rect 14108 24120 14136 24151
rect 14366 24148 14372 24200
rect 14424 24148 14430 24200
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 14599 24160 14964 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 14458 24120 14464 24132
rect 14108 24092 14464 24120
rect 14458 24080 14464 24092
rect 14516 24080 14522 24132
rect 10980 24024 12828 24052
rect 12894 24012 12900 24064
rect 12952 24052 12958 24064
rect 13265 24055 13323 24061
rect 13265 24052 13277 24055
rect 12952 24024 13277 24052
rect 12952 24012 12958 24024
rect 13265 24021 13277 24024
rect 13311 24021 13323 24055
rect 13265 24015 13323 24021
rect 13354 24012 13360 24064
rect 13412 24012 13418 24064
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24052 13783 24055
rect 13998 24052 14004 24064
rect 13771 24024 14004 24052
rect 13771 24021 13783 24024
rect 13725 24015 13783 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 14182 24012 14188 24064
rect 14240 24012 14246 24064
rect 14936 24052 14964 24160
rect 15010 24148 15016 24200
rect 15068 24188 15074 24200
rect 15185 24191 15243 24197
rect 15185 24188 15197 24191
rect 15068 24160 15197 24188
rect 15068 24148 15074 24160
rect 15185 24157 15197 24160
rect 15231 24157 15243 24191
rect 15185 24151 15243 24157
rect 15304 24120 15332 24228
rect 15378 24148 15384 24200
rect 15436 24148 15442 24200
rect 16298 24148 16304 24200
rect 16356 24148 16362 24200
rect 16684 24197 16712 24228
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24157 16727 24191
rect 16859 24188 16887 24296
rect 16960 24265 16988 24352
rect 18509 24327 18567 24333
rect 18509 24324 18521 24327
rect 17972 24296 18521 24324
rect 17972 24265 18000 24296
rect 18509 24293 18521 24296
rect 18555 24293 18567 24327
rect 18509 24287 18567 24293
rect 19245 24327 19303 24333
rect 19245 24293 19257 24327
rect 19291 24293 19303 24327
rect 19245 24287 19303 24293
rect 16945 24259 17003 24265
rect 16945 24225 16957 24259
rect 16991 24225 17003 24259
rect 17957 24259 18015 24265
rect 16945 24219 17003 24225
rect 17236 24228 17908 24256
rect 17129 24191 17187 24197
rect 17129 24188 17141 24191
rect 16859 24160 17141 24188
rect 16669 24151 16727 24157
rect 17129 24157 17141 24160
rect 17175 24157 17187 24191
rect 17129 24151 17187 24157
rect 17236 24120 17264 24228
rect 17773 24191 17831 24197
rect 17773 24188 17785 24191
rect 15304 24092 17264 24120
rect 17420 24160 17785 24188
rect 15470 24052 15476 24064
rect 14936 24024 15476 24052
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 15746 24012 15752 24064
rect 15804 24052 15810 24064
rect 15841 24055 15899 24061
rect 15841 24052 15853 24055
rect 15804 24024 15853 24052
rect 15804 24012 15810 24024
rect 15841 24021 15853 24024
rect 15887 24052 15899 24055
rect 17420 24052 17448 24160
rect 17773 24157 17785 24160
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 17880 24120 17908 24228
rect 17957 24225 17969 24259
rect 18003 24225 18015 24259
rect 19260 24256 19288 24287
rect 19536 24256 19564 24352
rect 17957 24219 18015 24225
rect 18708 24228 19288 24256
rect 19352 24228 19564 24256
rect 18708 24197 18736 24228
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 19061 24191 19119 24197
rect 19061 24157 19073 24191
rect 19107 24188 19119 24191
rect 19352 24188 19380 24228
rect 19107 24160 19380 24188
rect 19429 24191 19487 24197
rect 19107 24157 19119 24160
rect 19061 24151 19119 24157
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19521 24191 19579 24197
rect 19521 24188 19533 24191
rect 19475 24160 19533 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19521 24157 19533 24160
rect 19567 24188 19579 24191
rect 19628 24188 19656 24352
rect 21913 24327 21971 24333
rect 21913 24293 21925 24327
rect 21959 24324 21971 24327
rect 23658 24324 23664 24336
rect 21959 24296 23664 24324
rect 21959 24293 21971 24296
rect 21913 24287 21971 24293
rect 23658 24284 23664 24296
rect 23716 24284 23722 24336
rect 24688 24324 24716 24352
rect 24320 24296 24716 24324
rect 25133 24327 25191 24333
rect 22278 24256 22284 24268
rect 19567 24160 19656 24188
rect 19720 24228 21680 24256
rect 19567 24157 19579 24160
rect 19521 24151 19579 24157
rect 19720 24120 19748 24228
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 20714 24188 20720 24200
rect 19935 24160 20720 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 17880 24092 19748 24120
rect 20441 24123 20499 24129
rect 20441 24089 20453 24123
rect 20487 24120 20499 24123
rect 20622 24120 20628 24132
rect 20487 24092 20628 24120
rect 20487 24089 20499 24092
rect 20441 24083 20499 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 20824 24120 20852 24151
rect 20990 24148 20996 24200
rect 21048 24148 21054 24200
rect 21358 24120 21364 24132
rect 20824 24092 21364 24120
rect 21358 24080 21364 24092
rect 21416 24080 21422 24132
rect 21652 24129 21680 24228
rect 22112 24228 22284 24256
rect 22112 24197 22140 24228
rect 22278 24216 22284 24228
rect 22336 24216 22342 24268
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22235 24160 22416 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 22388 24132 22416 24160
rect 22462 24148 22468 24200
rect 22520 24148 22526 24200
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24157 23075 24191
rect 23017 24151 23075 24157
rect 21637 24123 21695 24129
rect 21637 24089 21649 24123
rect 21683 24089 21695 24123
rect 21637 24083 21695 24089
rect 22370 24080 22376 24132
rect 22428 24080 22434 24132
rect 23032 24120 23060 24151
rect 23106 24148 23112 24200
rect 23164 24148 23170 24200
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24188 23719 24191
rect 24121 24191 24179 24197
rect 24121 24188 24133 24191
rect 23707 24160 24133 24188
rect 23707 24157 23719 24160
rect 23661 24151 23719 24157
rect 24121 24157 24133 24160
rect 24167 24188 24179 24191
rect 24320 24188 24348 24296
rect 25133 24293 25145 24327
rect 25179 24324 25191 24327
rect 25976 24324 26004 24352
rect 25179 24296 26004 24324
rect 25179 24293 25191 24296
rect 25133 24287 25191 24293
rect 25961 24259 26019 24265
rect 25961 24256 25973 24259
rect 24688 24228 25973 24256
rect 24688 24200 24716 24228
rect 25961 24225 25973 24228
rect 26007 24225 26019 24259
rect 25961 24219 26019 24225
rect 24167 24160 24348 24188
rect 24489 24191 24547 24197
rect 24167 24157 24179 24160
rect 24121 24151 24179 24157
rect 24489 24157 24501 24191
rect 24535 24157 24547 24191
rect 24489 24151 24547 24157
rect 23842 24120 23848 24132
rect 23032 24092 23848 24120
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 24504 24120 24532 24151
rect 24670 24148 24676 24200
rect 24728 24148 24734 24200
rect 25317 24191 25375 24197
rect 25317 24157 25329 24191
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 25498 24188 25504 24200
rect 25455 24160 25504 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 24854 24120 24860 24132
rect 24504 24092 24860 24120
rect 24854 24080 24860 24092
rect 24912 24080 24918 24132
rect 25332 24120 25360 24151
rect 25498 24148 25504 24160
rect 25556 24148 25562 24200
rect 25590 24148 25596 24200
rect 25648 24148 25654 24200
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24188 25927 24191
rect 26050 24188 26056 24200
rect 25915 24160 26056 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 26510 24188 26516 24200
rect 26160 24160 26516 24188
rect 25608 24120 25636 24148
rect 25332 24092 25636 24120
rect 15887 24024 17448 24052
rect 15887 24021 15899 24024
rect 15841 24015 15899 24021
rect 17586 24012 17592 24064
rect 17644 24012 17650 24064
rect 18874 24012 18880 24064
rect 18932 24012 18938 24064
rect 19610 24012 19616 24064
rect 19668 24012 19674 24064
rect 21450 24012 21456 24064
rect 21508 24012 21514 24064
rect 21542 24012 21548 24064
rect 21600 24052 21606 24064
rect 21729 24055 21787 24061
rect 21729 24052 21741 24055
rect 21600 24024 21741 24052
rect 21600 24012 21606 24024
rect 21729 24021 21741 24024
rect 21775 24021 21787 24055
rect 21729 24015 21787 24021
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 22281 24055 22339 24061
rect 22281 24052 22293 24055
rect 22244 24024 22293 24052
rect 22244 24012 22250 24024
rect 22281 24021 22293 24024
rect 22327 24021 22339 24055
rect 22281 24015 22339 24021
rect 22554 24012 22560 24064
rect 22612 24012 22618 24064
rect 22830 24012 22836 24064
rect 22888 24012 22894 24064
rect 23198 24012 23204 24064
rect 23256 24012 23262 24064
rect 23750 24012 23756 24064
rect 23808 24012 23814 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 25004 24024 25053 24052
rect 25004 24012 25010 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25041 24015 25099 24021
rect 25685 24055 25743 24061
rect 25685 24021 25697 24055
rect 25731 24052 25743 24055
rect 26160 24052 26188 24160
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 27433 24191 27491 24197
rect 27433 24188 27445 24191
rect 27356 24160 27445 24188
rect 26228 24123 26286 24129
rect 26228 24089 26240 24123
rect 26274 24120 26286 24123
rect 26786 24120 26792 24132
rect 26274 24092 26792 24120
rect 26274 24089 26286 24092
rect 26228 24083 26286 24089
rect 26786 24080 26792 24092
rect 26844 24080 26850 24132
rect 25731 24024 26188 24052
rect 25731 24021 25743 24024
rect 25685 24015 25743 24021
rect 27154 24012 27160 24064
rect 27212 24052 27218 24064
rect 27356 24061 27384 24160
rect 27433 24157 27445 24160
rect 27479 24157 27491 24191
rect 27433 24151 27491 24157
rect 27890 24080 27896 24132
rect 27948 24080 27954 24132
rect 27985 24123 28043 24129
rect 27985 24089 27997 24123
rect 28031 24120 28043 24123
rect 28074 24120 28080 24132
rect 28031 24092 28080 24120
rect 28031 24089 28043 24092
rect 27985 24083 28043 24089
rect 28074 24080 28080 24092
rect 28132 24080 28138 24132
rect 28258 24080 28264 24132
rect 28316 24120 28322 24132
rect 28537 24123 28595 24129
rect 28537 24120 28549 24123
rect 28316 24092 28549 24120
rect 28316 24080 28322 24092
rect 28537 24089 28549 24092
rect 28583 24089 28595 24123
rect 28537 24083 28595 24089
rect 27341 24055 27399 24061
rect 27341 24052 27353 24055
rect 27212 24024 27353 24052
rect 27212 24012 27218 24024
rect 27341 24021 27353 24024
rect 27387 24021 27399 24055
rect 27341 24015 27399 24021
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 2130 23808 2136 23860
rect 2188 23808 2194 23860
rect 3605 23851 3663 23857
rect 3605 23817 3617 23851
rect 3651 23848 3663 23851
rect 3786 23848 3792 23860
rect 3651 23820 3792 23848
rect 3651 23817 3663 23820
rect 3605 23811 3663 23817
rect 3786 23808 3792 23820
rect 3844 23848 3850 23860
rect 3844 23820 4016 23848
rect 3844 23808 3850 23820
rect 3878 23780 3884 23792
rect 2240 23752 3884 23780
rect 2240 23724 2268 23752
rect 3878 23740 3884 23752
rect 3936 23740 3942 23792
rect 2222 23672 2228 23724
rect 2280 23672 2286 23724
rect 2492 23715 2550 23721
rect 2492 23681 2504 23715
rect 2538 23712 2550 23715
rect 3510 23712 3516 23724
rect 2538 23684 3516 23712
rect 2538 23681 2550 23684
rect 2492 23675 2550 23681
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 3988 23721 4016 23820
rect 4890 23808 4896 23860
rect 4948 23808 4954 23860
rect 6086 23808 6092 23860
rect 6144 23808 6150 23860
rect 6270 23808 6276 23860
rect 6328 23808 6334 23860
rect 6546 23808 6552 23860
rect 6604 23848 6610 23860
rect 7009 23851 7067 23857
rect 7009 23848 7021 23851
rect 6604 23820 7021 23848
rect 6604 23808 6610 23820
rect 7009 23817 7021 23820
rect 7055 23817 7067 23851
rect 7009 23811 7067 23817
rect 7558 23808 7564 23860
rect 7616 23808 7622 23860
rect 7742 23808 7748 23860
rect 7800 23848 7806 23860
rect 8662 23848 8668 23860
rect 7800 23820 8668 23848
rect 7800 23808 7806 23820
rect 8662 23808 8668 23820
rect 8720 23808 8726 23860
rect 9033 23851 9091 23857
rect 9033 23817 9045 23851
rect 9079 23848 9091 23851
rect 9079 23820 9720 23848
rect 9079 23817 9091 23820
rect 9033 23811 9091 23817
rect 4908 23780 4936 23808
rect 4908 23752 5672 23780
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23681 4031 23715
rect 3973 23675 4031 23681
rect 4617 23715 4675 23721
rect 4617 23681 4629 23715
rect 4663 23712 4675 23715
rect 4982 23712 4988 23724
rect 4663 23684 4988 23712
rect 4663 23681 4675 23684
rect 4617 23675 4675 23681
rect 4982 23672 4988 23684
rect 5040 23672 5046 23724
rect 5644 23721 5672 23752
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5629 23715 5687 23721
rect 5123 23684 5580 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 1581 23647 1639 23653
rect 1581 23613 1593 23647
rect 1627 23613 1639 23647
rect 1581 23607 1639 23613
rect 1596 23508 1624 23607
rect 3234 23604 3240 23656
rect 3292 23644 3298 23656
rect 5092 23644 5120 23675
rect 3292 23616 5120 23644
rect 3292 23604 3298 23616
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 5552 23644 5580 23684
rect 5629 23681 5641 23715
rect 5675 23681 5687 23715
rect 6104 23712 6132 23808
rect 6288 23780 6316 23808
rect 7576 23780 7604 23808
rect 6288 23752 6592 23780
rect 6564 23721 6592 23752
rect 7116 23752 7604 23780
rect 7116 23721 7144 23752
rect 8202 23740 8208 23792
rect 8260 23780 8266 23792
rect 9692 23789 9720 23820
rect 10226 23808 10232 23860
rect 10284 23808 10290 23860
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 10376 23820 10548 23848
rect 10376 23808 10382 23820
rect 9585 23783 9643 23789
rect 9585 23780 9597 23783
rect 8260 23752 9597 23780
rect 8260 23740 8266 23752
rect 9585 23749 9597 23752
rect 9631 23749 9643 23783
rect 9585 23743 9643 23749
rect 9677 23783 9735 23789
rect 9677 23749 9689 23783
rect 9723 23749 9735 23783
rect 9677 23743 9735 23749
rect 10244 23780 10272 23808
rect 10520 23789 10548 23820
rect 11698 23808 11704 23860
rect 11756 23848 11762 23860
rect 11756 23820 11928 23848
rect 11756 23808 11762 23820
rect 11900 23789 11928 23820
rect 12802 23808 12808 23860
rect 12860 23808 12866 23860
rect 13354 23808 13360 23860
rect 13412 23808 13418 23860
rect 14001 23851 14059 23857
rect 14001 23817 14013 23851
rect 14047 23848 14059 23851
rect 14090 23848 14096 23860
rect 14047 23820 14096 23848
rect 14047 23817 14059 23820
rect 14001 23811 14059 23817
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14182 23808 14188 23860
rect 14240 23808 14246 23860
rect 14734 23808 14740 23860
rect 14792 23848 14798 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 14792 23820 14933 23848
rect 14792 23808 14798 23820
rect 14921 23817 14933 23820
rect 14967 23817 14979 23851
rect 14921 23811 14979 23817
rect 15378 23808 15384 23860
rect 15436 23848 15442 23860
rect 16117 23851 16175 23857
rect 16117 23848 16129 23851
rect 15436 23820 16129 23848
rect 15436 23808 15442 23820
rect 16117 23817 16129 23820
rect 16163 23817 16175 23851
rect 16117 23811 16175 23817
rect 18230 23808 18236 23860
rect 18288 23808 18294 23860
rect 18800 23820 20116 23848
rect 10413 23783 10471 23789
rect 10413 23780 10425 23783
rect 10244 23752 10425 23780
rect 6365 23715 6423 23721
rect 6365 23712 6377 23715
rect 6104 23684 6377 23712
rect 5629 23675 5687 23681
rect 6365 23681 6377 23684
rect 6411 23681 6423 23715
rect 6365 23675 6423 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 7101 23715 7159 23721
rect 7101 23681 7113 23715
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 5994 23644 6000 23656
rect 5552 23616 6000 23644
rect 5994 23604 6000 23616
rect 6052 23644 6058 23656
rect 7116 23644 7144 23675
rect 7190 23672 7196 23724
rect 7248 23712 7254 23724
rect 7561 23715 7619 23721
rect 7561 23712 7573 23715
rect 7248 23684 7573 23712
rect 7248 23672 7254 23684
rect 7561 23681 7573 23684
rect 7607 23681 7619 23715
rect 7561 23675 7619 23681
rect 7650 23672 7656 23724
rect 7708 23672 7714 23724
rect 8662 23672 8668 23724
rect 8720 23712 8726 23724
rect 10244 23721 10272 23752
rect 10413 23749 10425 23752
rect 10459 23749 10471 23783
rect 10413 23743 10471 23749
rect 10505 23783 10563 23789
rect 10505 23749 10517 23783
rect 10551 23749 10563 23783
rect 10505 23743 10563 23749
rect 11885 23783 11943 23789
rect 11885 23749 11897 23783
rect 11931 23749 11943 23783
rect 11885 23743 11943 23749
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 8720 23684 9229 23712
rect 8720 23672 8726 23684
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23681 10287 23715
rect 11333 23715 11391 23721
rect 11333 23712 11345 23715
rect 10229 23675 10287 23681
rect 11072 23684 11345 23712
rect 6052 23616 7144 23644
rect 6052 23604 6058 23616
rect 7374 23604 7380 23656
rect 7432 23604 7438 23656
rect 4338 23536 4344 23588
rect 4396 23576 4402 23588
rect 4709 23579 4767 23585
rect 4709 23576 4721 23579
rect 4396 23548 4721 23576
rect 4396 23536 4402 23548
rect 4709 23545 4721 23548
rect 4755 23545 4767 23579
rect 4709 23539 4767 23545
rect 6914 23536 6920 23588
rect 6972 23576 6978 23588
rect 7668 23576 7696 23672
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 8297 23647 8355 23653
rect 8297 23644 8309 23647
rect 8260 23616 8309 23644
rect 8260 23604 8266 23616
rect 8297 23613 8309 23616
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 8481 23647 8539 23653
rect 8481 23613 8493 23647
rect 8527 23613 8539 23647
rect 8481 23607 8539 23613
rect 8496 23576 8524 23607
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10410 23644 10416 23656
rect 9916 23616 10416 23644
rect 9916 23604 9922 23616
rect 10410 23604 10416 23616
rect 10468 23644 10474 23656
rect 11072 23644 11100 23684
rect 11333 23681 11345 23684
rect 11379 23681 11391 23715
rect 12820 23712 12848 23808
rect 12877 23715 12935 23721
rect 12877 23712 12889 23715
rect 12820 23684 12889 23712
rect 11333 23675 11391 23681
rect 12877 23681 12889 23684
rect 12923 23681 12935 23715
rect 13372 23712 13400 23808
rect 14200 23712 14228 23808
rect 15841 23783 15899 23789
rect 15841 23749 15853 23783
rect 15887 23780 15899 23783
rect 15887 23752 16344 23780
rect 15887 23749 15899 23752
rect 15841 23743 15899 23749
rect 14277 23715 14335 23721
rect 14277 23712 14289 23715
rect 13372 23684 13952 23712
rect 14200 23684 14289 23712
rect 12877 23675 12935 23681
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 10468 23616 11100 23644
rect 11256 23616 11805 23644
rect 10468 23604 10474 23616
rect 6972 23548 7420 23576
rect 7668 23548 8524 23576
rect 6972 23536 6978 23548
rect 2590 23508 2596 23520
rect 1596 23480 2596 23508
rect 2590 23468 2596 23480
rect 2648 23468 2654 23520
rect 4246 23468 4252 23520
rect 4304 23508 4310 23520
rect 4525 23511 4583 23517
rect 4525 23508 4537 23511
rect 4304 23480 4537 23508
rect 4304 23468 4310 23480
rect 4525 23477 4537 23480
rect 4571 23477 4583 23511
rect 4525 23471 4583 23477
rect 5166 23468 5172 23520
rect 5224 23468 5230 23520
rect 7190 23468 7196 23520
rect 7248 23468 7254 23520
rect 7392 23508 7420 23548
rect 8570 23536 8576 23588
rect 8628 23576 8634 23588
rect 8628 23548 8800 23576
rect 8628 23536 8634 23548
rect 7742 23508 7748 23520
rect 7392 23480 7748 23508
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 8662 23468 8668 23520
rect 8720 23468 8726 23520
rect 8772 23508 8800 23548
rect 9214 23536 9220 23588
rect 9272 23576 9278 23588
rect 9876 23576 9904 23604
rect 11256 23588 11284 23616
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 12250 23644 12256 23656
rect 11793 23607 11851 23613
rect 11900 23616 12256 23644
rect 9272 23548 9904 23576
rect 9272 23536 9278 23548
rect 10962 23536 10968 23588
rect 11020 23536 11026 23588
rect 11238 23536 11244 23588
rect 11296 23536 11302 23588
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 11900 23576 11928 23616
rect 12250 23604 12256 23616
rect 12308 23644 12314 23656
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12308 23616 12633 23644
rect 12308 23604 12314 23616
rect 12621 23613 12633 23616
rect 12667 23613 12679 23647
rect 13924 23644 13952 23684
rect 14277 23681 14289 23684
rect 14323 23681 14335 23715
rect 15289 23715 15347 23721
rect 15289 23712 15301 23715
rect 14277 23675 14335 23681
rect 15212 23684 15301 23712
rect 14461 23647 14519 23653
rect 14461 23644 14473 23647
rect 13924 23616 14473 23644
rect 12621 23607 12679 23613
rect 14461 23613 14473 23616
rect 14507 23613 14519 23647
rect 14461 23607 14519 23613
rect 11572 23548 11928 23576
rect 11572 23536 11578 23548
rect 12066 23536 12072 23588
rect 12124 23576 12130 23588
rect 12345 23579 12403 23585
rect 12345 23576 12357 23579
rect 12124 23548 12357 23576
rect 12124 23536 12130 23548
rect 12345 23545 12357 23548
rect 12391 23545 12403 23579
rect 12345 23539 12403 23545
rect 9490 23508 9496 23520
rect 8772 23480 9496 23508
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 11698 23508 11704 23520
rect 11195 23480 11704 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 15212 23508 15240 23684
rect 15289 23681 15301 23684
rect 15335 23681 15347 23715
rect 15289 23675 15347 23681
rect 16022 23672 16028 23724
rect 16080 23672 16086 23724
rect 16316 23712 16344 23752
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 16316 23684 16957 23712
rect 16316 23656 16344 23684
rect 16945 23681 16957 23684
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17586 23672 17592 23724
rect 17644 23712 17650 23724
rect 17865 23715 17923 23721
rect 17865 23712 17877 23715
rect 17644 23684 17877 23712
rect 17644 23672 17650 23684
rect 17865 23681 17877 23684
rect 17911 23681 17923 23715
rect 17865 23675 17923 23681
rect 16298 23604 16304 23656
rect 16356 23604 16362 23656
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 18248 23644 18276 23808
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23712 18659 23715
rect 18800 23712 18828 23820
rect 20088 23792 20116 23820
rect 20990 23808 20996 23860
rect 21048 23848 21054 23860
rect 23566 23848 23572 23860
rect 21048 23820 23572 23848
rect 21048 23808 21054 23820
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 23750 23808 23756 23860
rect 23808 23848 23814 23860
rect 23808 23820 25176 23848
rect 23808 23808 23814 23820
rect 18874 23740 18880 23792
rect 18932 23780 18938 23792
rect 19153 23783 19211 23789
rect 19153 23780 19165 23783
rect 18932 23752 19165 23780
rect 18932 23740 18938 23752
rect 19153 23749 19165 23752
rect 19199 23749 19211 23783
rect 19153 23743 19211 23749
rect 19702 23740 19708 23792
rect 19760 23740 19766 23792
rect 19978 23740 19984 23792
rect 20036 23740 20042 23792
rect 20070 23740 20076 23792
rect 20128 23780 20134 23792
rect 23198 23780 23204 23792
rect 20128 23752 22784 23780
rect 20128 23740 20134 23752
rect 18647 23684 18828 23712
rect 19720 23712 19748 23740
rect 19797 23715 19855 23721
rect 19797 23712 19809 23715
rect 19720 23684 19809 23712
rect 18647 23681 18659 23684
rect 18601 23675 18659 23681
rect 19797 23681 19809 23684
rect 19843 23681 19855 23715
rect 19797 23675 19855 23681
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21508 23684 21833 23712
rect 21508 23672 21514 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23712 22063 23715
rect 22554 23712 22560 23724
rect 22051 23684 22560 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 22554 23672 22560 23684
rect 22612 23672 22618 23724
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18248 23616 19073 23644
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23644 19763 23647
rect 20254 23644 20260 23656
rect 19751 23616 20260 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 20622 23604 20628 23656
rect 20680 23644 20686 23656
rect 21266 23644 21272 23656
rect 20680 23616 21272 23644
rect 20680 23604 20686 23616
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 22370 23644 22376 23656
rect 21324 23616 22376 23644
rect 21324 23604 21330 23616
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 22646 23604 22652 23656
rect 22704 23604 22710 23656
rect 22756 23644 22784 23752
rect 22848 23752 23204 23780
rect 22848 23721 22876 23752
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 25038 23780 25044 23792
rect 23308 23752 25044 23780
rect 22833 23715 22891 23721
rect 22833 23681 22845 23715
rect 22879 23681 22891 23715
rect 22833 23675 22891 23681
rect 23308 23644 23336 23752
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 25148 23789 25176 23820
rect 26786 23808 26792 23860
rect 26844 23808 26850 23860
rect 27982 23808 27988 23860
rect 28040 23808 28046 23860
rect 28350 23808 28356 23860
rect 28408 23808 28414 23860
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23749 25191 23783
rect 25133 23743 25191 23749
rect 27240 23783 27298 23789
rect 27240 23749 27252 23783
rect 27286 23780 27298 23783
rect 28000 23780 28028 23808
rect 27286 23752 28028 23780
rect 27286 23749 27298 23752
rect 27240 23743 27298 23749
rect 23474 23672 23480 23724
rect 23532 23672 23538 23724
rect 23744 23715 23802 23721
rect 23744 23681 23756 23715
rect 23790 23712 23802 23715
rect 24578 23712 24584 23724
rect 23790 23684 24584 23712
rect 23790 23681 23802 23684
rect 23744 23675 23802 23681
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 26050 23672 26056 23724
rect 26108 23712 26114 23724
rect 26145 23715 26203 23721
rect 26145 23712 26157 23715
rect 26108 23684 26157 23712
rect 26108 23672 26114 23684
rect 26145 23681 26157 23684
rect 26191 23681 26203 23715
rect 26145 23675 26203 23681
rect 25041 23647 25099 23653
rect 25041 23644 25053 23647
rect 22756 23616 23336 23644
rect 24504 23616 25053 23644
rect 18509 23579 18567 23585
rect 18509 23545 18521 23579
rect 18555 23576 18567 23579
rect 19334 23576 19340 23588
rect 18555 23548 19340 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 19334 23536 19340 23548
rect 19392 23536 19398 23588
rect 12860 23480 15240 23508
rect 12860 23468 12866 23480
rect 17034 23468 17040 23520
rect 17092 23468 17098 23520
rect 18693 23511 18751 23517
rect 18693 23477 18705 23511
rect 18739 23508 18751 23511
rect 19978 23508 19984 23520
rect 18739 23480 19984 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 22186 23468 22192 23520
rect 22244 23468 22250 23520
rect 23293 23511 23351 23517
rect 23293 23477 23305 23511
rect 23339 23508 23351 23511
rect 23382 23508 23388 23520
rect 23339 23480 23388 23508
rect 23339 23477 23351 23480
rect 23293 23471 23351 23477
rect 23382 23468 23388 23480
rect 23440 23508 23446 23520
rect 24504 23508 24532 23616
rect 25041 23613 25053 23616
rect 25087 23613 25099 23647
rect 25041 23607 25099 23613
rect 25130 23604 25136 23656
rect 25188 23644 25194 23656
rect 25317 23647 25375 23653
rect 25317 23644 25329 23647
rect 25188 23616 25329 23644
rect 25188 23604 25194 23616
rect 25317 23613 25329 23616
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 26973 23647 27031 23653
rect 26973 23613 26985 23647
rect 27019 23613 27031 23647
rect 26973 23607 27031 23613
rect 24670 23536 24676 23588
rect 24728 23576 24734 23588
rect 26988 23576 27016 23607
rect 24728 23548 27016 23576
rect 24728 23536 24734 23548
rect 23440 23480 24532 23508
rect 23440 23468 23446 23480
rect 24854 23468 24860 23520
rect 24912 23468 24918 23520
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 28258 23508 28264 23520
rect 25096 23480 28264 23508
rect 25096 23468 25102 23480
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 2590 23264 2596 23316
rect 2648 23304 2654 23316
rect 2777 23307 2835 23313
rect 2777 23304 2789 23307
rect 2648 23276 2789 23304
rect 2648 23264 2654 23276
rect 2777 23273 2789 23276
rect 2823 23273 2835 23307
rect 3970 23304 3976 23316
rect 2777 23267 2835 23273
rect 3436 23276 3976 23304
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3145 23171 3203 23177
rect 3145 23168 3157 23171
rect 2832 23140 3157 23168
rect 2832 23128 2838 23140
rect 3145 23137 3157 23140
rect 3191 23137 3203 23171
rect 3145 23131 3203 23137
rect 1394 23060 1400 23112
rect 1452 23100 1458 23112
rect 2222 23100 2228 23112
rect 1452 23072 2228 23100
rect 1452 23060 1458 23072
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 3436 23100 3464 23276
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 5040 23276 5181 23304
rect 5040 23264 5046 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 5169 23267 5227 23273
rect 5629 23307 5687 23313
rect 5629 23273 5641 23307
rect 5675 23304 5687 23307
rect 7193 23307 7251 23313
rect 5675 23276 6868 23304
rect 5675 23273 5687 23276
rect 5629 23267 5687 23273
rect 4890 23196 4896 23248
rect 4948 23236 4954 23248
rect 5644 23236 5672 23267
rect 4948 23208 5672 23236
rect 4948 23196 4954 23208
rect 3007 23072 3464 23100
rect 3789 23103 3847 23109
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 3789 23069 3801 23103
rect 3835 23100 3847 23103
rect 3878 23100 3884 23112
rect 3835 23072 3884 23100
rect 3835 23069 3847 23072
rect 3789 23063 3847 23069
rect 3878 23060 3884 23072
rect 3936 23100 3942 23112
rect 5813 23103 5871 23109
rect 5813 23100 5825 23103
rect 3936 23072 5825 23100
rect 3936 23060 3942 23072
rect 5813 23069 5825 23072
rect 5859 23100 5871 23103
rect 6840 23100 6868 23276
rect 7193 23273 7205 23307
rect 7239 23304 7251 23307
rect 7282 23304 7288 23316
rect 7239 23276 7288 23304
rect 7239 23273 7251 23276
rect 7193 23267 7251 23273
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 7742 23264 7748 23316
rect 7800 23264 7806 23316
rect 8662 23264 8668 23316
rect 8720 23264 8726 23316
rect 8941 23307 8999 23313
rect 8941 23273 8953 23307
rect 8987 23304 8999 23307
rect 11146 23304 11152 23316
rect 8987 23276 11152 23304
rect 8987 23273 8999 23276
rect 8941 23267 8999 23273
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 11900 23276 16804 23304
rect 8680 23236 8708 23264
rect 7392 23208 8708 23236
rect 9217 23239 9275 23245
rect 7392 23177 7420 23208
rect 9217 23205 9229 23239
rect 9263 23236 9275 23239
rect 10318 23236 10324 23248
rect 9263 23208 10324 23236
rect 9263 23205 9275 23208
rect 9217 23199 9275 23205
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 7377 23171 7435 23177
rect 7377 23137 7389 23171
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 7466 23128 7472 23180
rect 7524 23168 7530 23180
rect 7561 23171 7619 23177
rect 7561 23168 7573 23171
rect 7524 23140 7573 23168
rect 7524 23128 7530 23140
rect 7561 23137 7573 23140
rect 7607 23137 7619 23171
rect 7561 23131 7619 23137
rect 7668 23140 8248 23168
rect 7668 23100 7696 23140
rect 5859 23072 6776 23100
rect 6840 23072 7696 23100
rect 8113 23103 8171 23109
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6748 23044 6776 23072
rect 8113 23069 8125 23103
rect 8159 23069 8171 23103
rect 8220 23100 8248 23140
rect 8294 23128 8300 23180
rect 8352 23128 8358 23180
rect 10226 23168 10232 23180
rect 8404 23140 10232 23168
rect 8404 23100 8432 23140
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 10781 23171 10839 23177
rect 10781 23137 10793 23171
rect 10827 23168 10839 23171
rect 11238 23168 11244 23180
rect 10827 23140 11244 23168
rect 10827 23137 10839 23140
rect 10781 23131 10839 23137
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 11900 23112 11928 23276
rect 11977 23171 12035 23177
rect 11977 23137 11989 23171
rect 12023 23168 12035 23171
rect 12066 23168 12072 23180
rect 12023 23140 12072 23168
rect 12023 23137 12035 23140
rect 11977 23131 12035 23137
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 12802 23128 12808 23180
rect 12860 23128 12866 23180
rect 13998 23128 14004 23180
rect 14056 23168 14062 23180
rect 15013 23171 15071 23177
rect 15013 23168 15025 23171
rect 14056 23140 15025 23168
rect 14056 23128 14062 23140
rect 15013 23137 15025 23140
rect 15059 23137 15071 23171
rect 15013 23131 15071 23137
rect 8220 23072 8432 23100
rect 8113 23063 8171 23069
rect 1664 23035 1722 23041
rect 1664 23001 1676 23035
rect 1710 23032 1722 23035
rect 3326 23032 3332 23044
rect 1710 23004 3332 23032
rect 1710 23001 1722 23004
rect 1664 22995 1722 23001
rect 3326 22992 3332 23004
rect 3384 22992 3390 23044
rect 4056 23035 4114 23041
rect 4056 23001 4068 23035
rect 4102 23032 4114 23035
rect 4246 23032 4252 23044
rect 4102 23004 4252 23032
rect 4102 23001 4114 23004
rect 4056 22995 4114 23001
rect 4246 22992 4252 23004
rect 4304 22992 4310 23044
rect 5350 22992 5356 23044
rect 5408 22992 5414 23044
rect 6080 23035 6138 23041
rect 6080 23001 6092 23035
rect 6126 23032 6138 23035
rect 6126 23004 6684 23032
rect 6126 23001 6138 23004
rect 6080 22995 6138 23001
rect 3605 22967 3663 22973
rect 3605 22933 3617 22967
rect 3651 22964 3663 22967
rect 4154 22964 4160 22976
rect 3651 22936 4160 22964
rect 3651 22933 3663 22936
rect 3605 22927 3663 22933
rect 4154 22924 4160 22936
rect 4212 22924 4218 22976
rect 6656 22964 6684 23004
rect 6730 22992 6736 23044
rect 6788 22992 6794 23044
rect 7098 22992 7104 23044
rect 7156 23032 7162 23044
rect 7742 23032 7748 23044
rect 7156 23004 7748 23032
rect 7156 22992 7162 23004
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 8128 23032 8156 23063
rect 8570 23060 8576 23112
rect 8628 23060 8634 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9214 23100 9220 23112
rect 9171 23072 9220 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9364 23072 9413 23100
rect 9364 23060 9370 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9490 23060 9496 23112
rect 9548 23060 9554 23112
rect 9582 23060 9588 23112
rect 9640 23060 9646 23112
rect 9769 23103 9827 23109
rect 9769 23069 9781 23103
rect 9815 23100 9827 23103
rect 9858 23100 9864 23112
rect 9815 23072 9864 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 9858 23060 9864 23072
rect 9916 23060 9922 23112
rect 11882 23060 11888 23112
rect 11940 23060 11946 23112
rect 14090 23060 14096 23112
rect 14148 23060 14154 23112
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 14829 23103 14887 23109
rect 14829 23100 14841 23103
rect 14332 23072 14841 23100
rect 14332 23060 14338 23072
rect 14829 23069 14841 23072
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23100 15807 23103
rect 16574 23100 16580 23112
rect 15795 23072 16580 23100
rect 15795 23069 15807 23072
rect 15749 23063 15807 23069
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 8588 23032 8616 23060
rect 9600 23032 9628 23060
rect 8128 23004 9628 23032
rect 10134 22992 10140 23044
rect 10192 22992 10198 23044
rect 10229 23035 10287 23041
rect 10229 23001 10241 23035
rect 10275 23001 10287 23035
rect 10229 22995 10287 23001
rect 7650 22964 7656 22976
rect 6656 22936 7656 22964
rect 7650 22924 7656 22936
rect 7708 22924 7714 22976
rect 9585 22967 9643 22973
rect 9585 22933 9597 22967
rect 9631 22964 9643 22967
rect 9766 22964 9772 22976
rect 9631 22936 9772 22964
rect 9631 22933 9643 22936
rect 9585 22927 9643 22933
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 9861 22967 9919 22973
rect 9861 22933 9873 22967
rect 9907 22964 9919 22967
rect 10244 22964 10272 22995
rect 10962 22992 10968 23044
rect 11020 22992 11026 23044
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 11790 22992 11796 23044
rect 11848 23032 11854 23044
rect 12253 23035 12311 23041
rect 12253 23032 12265 23035
rect 11848 23004 12265 23032
rect 11848 22992 11854 23004
rect 12253 23001 12265 23004
rect 12299 23001 12311 23035
rect 12253 22995 12311 23001
rect 16016 23035 16074 23041
rect 16016 23001 16028 23035
rect 16062 23032 16074 23035
rect 16482 23032 16488 23044
rect 16062 23004 16488 23032
rect 16062 23001 16074 23004
rect 16016 22995 16074 23001
rect 16482 22992 16488 23004
rect 16540 22992 16546 23044
rect 16776 23032 16804 23276
rect 17586 23264 17592 23316
rect 17644 23264 17650 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 18104 23276 18705 23304
rect 18104 23264 18110 23276
rect 18693 23273 18705 23276
rect 18739 23273 18751 23307
rect 18693 23267 18751 23273
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 21450 23304 21456 23316
rect 21407 23276 21456 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 23201 23307 23259 23313
rect 22244 23276 22784 23304
rect 22244 23264 22250 23276
rect 17957 23239 18015 23245
rect 17957 23205 17969 23239
rect 18003 23205 18015 23239
rect 20990 23236 20996 23248
rect 17957 23199 18015 23205
rect 20732 23208 20996 23236
rect 17034 23128 17040 23180
rect 17092 23168 17098 23180
rect 17405 23171 17463 23177
rect 17405 23168 17417 23171
rect 17092 23140 17417 23168
rect 17092 23128 17098 23140
rect 17405 23137 17417 23140
rect 17451 23137 17463 23171
rect 17972 23168 18000 23199
rect 17972 23140 18920 23168
rect 17405 23131 17463 23137
rect 17218 23060 17224 23112
rect 17276 23060 17282 23112
rect 17586 23060 17592 23112
rect 17644 23100 17650 23112
rect 18892 23109 18920 23140
rect 19702 23128 19708 23180
rect 19760 23128 19766 23180
rect 20732 23177 20760 23208
rect 20990 23196 20996 23208
rect 21048 23236 21054 23248
rect 21542 23236 21548 23248
rect 21048 23208 21548 23236
rect 21048 23196 21054 23208
rect 21542 23196 21548 23208
rect 21600 23196 21606 23248
rect 22388 23208 22600 23236
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23137 20775 23171
rect 20717 23131 20775 23137
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23168 20959 23171
rect 22094 23168 22100 23180
rect 20947 23140 22100 23168
rect 20947 23137 20959 23140
rect 20901 23131 20959 23137
rect 22094 23128 22100 23140
rect 22152 23128 22158 23180
rect 22388 23168 22416 23208
rect 22204 23140 22416 23168
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17644 23072 18153 23100
rect 17644 23060 17650 23072
rect 18141 23069 18153 23072
rect 18187 23100 18199 23103
rect 18417 23103 18475 23109
rect 18417 23100 18429 23103
rect 18187 23072 18429 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18417 23069 18429 23072
rect 18463 23100 18475 23103
rect 18877 23103 18935 23109
rect 18463 23072 18736 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 18708 23032 18736 23072
rect 18877 23069 18889 23103
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 20441 23103 20499 23109
rect 20441 23069 20453 23103
rect 20487 23100 20499 23103
rect 20622 23100 20628 23112
rect 20487 23072 20628 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21545 23103 21603 23109
rect 21545 23100 21557 23103
rect 20864 23072 21557 23100
rect 20864 23060 20870 23072
rect 21545 23069 21557 23072
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22204 23100 22232 23140
rect 21775 23072 22232 23100
rect 22281 23103 22339 23109
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 22281 23069 22293 23103
rect 22327 23100 22339 23103
rect 22462 23100 22468 23112
rect 22327 23072 22468 23100
rect 22327 23069 22339 23072
rect 22281 23063 22339 23069
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 18966 23032 18972 23044
rect 16776 23004 18644 23032
rect 18708 23004 18972 23032
rect 9907 22936 10272 22964
rect 9907 22933 9919 22936
rect 9861 22927 9919 22933
rect 14734 22924 14740 22976
rect 14792 22924 14798 22976
rect 15194 22924 15200 22976
rect 15252 22964 15258 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15252 22936 15485 22964
rect 15252 22924 15258 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 18506 22924 18512 22976
rect 18564 22924 18570 22976
rect 18616 22964 18644 23004
rect 18966 22992 18972 23004
rect 19024 22992 19030 23044
rect 19334 22992 19340 23044
rect 19392 22992 19398 23044
rect 19429 23035 19487 23041
rect 19429 23001 19441 23035
rect 19475 23032 19487 23035
rect 19610 23032 19616 23044
rect 19475 23004 19616 23032
rect 19475 23001 19487 23004
rect 19429 22995 19487 23001
rect 19610 22992 19616 23004
rect 19668 22992 19674 23044
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 21634 23032 21640 23044
rect 20772 23004 21640 23032
rect 20772 22992 20778 23004
rect 21634 22992 21640 23004
rect 21692 22992 21698 23044
rect 22066 23004 22416 23032
rect 19886 22964 19892 22976
rect 18616 22936 19892 22964
rect 19886 22924 19892 22936
rect 19944 22924 19950 22976
rect 20533 22967 20591 22973
rect 20533 22933 20545 22967
rect 20579 22964 20591 22967
rect 20898 22964 20904 22976
rect 20579 22936 20904 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 21542 22924 21548 22976
rect 21600 22964 21606 22976
rect 22066 22964 22094 23004
rect 22388 22973 22416 23004
rect 21600 22936 22094 22964
rect 22373 22967 22431 22973
rect 21600 22924 21606 22936
rect 22373 22933 22385 22967
rect 22419 22933 22431 22967
rect 22572 22964 22600 23208
rect 22649 23171 22707 23177
rect 22649 23137 22661 23171
rect 22695 23168 22707 23171
rect 22756 23168 22784 23276
rect 23201 23273 23213 23307
rect 23247 23304 23259 23307
rect 23382 23304 23388 23316
rect 23247 23276 23388 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 23661 23307 23719 23313
rect 23661 23304 23673 23307
rect 23624 23276 23673 23304
rect 23624 23264 23630 23276
rect 23661 23273 23673 23276
rect 23707 23273 23719 23307
rect 23661 23267 23719 23273
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 23900 23276 24409 23304
rect 23900 23264 23906 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 26050 23264 26056 23316
rect 26108 23264 26114 23316
rect 27154 23304 27160 23316
rect 26252 23276 27160 23304
rect 23290 23196 23296 23248
rect 23348 23236 23354 23248
rect 23937 23239 23995 23245
rect 23937 23236 23949 23239
rect 23348 23208 23949 23236
rect 23348 23196 23354 23208
rect 23937 23205 23949 23208
rect 23983 23205 23995 23239
rect 23937 23199 23995 23205
rect 22695 23140 22784 23168
rect 22695 23137 22707 23140
rect 22649 23131 22707 23137
rect 22830 23128 22836 23180
rect 22888 23128 22894 23180
rect 23474 23128 23480 23180
rect 23532 23168 23538 23180
rect 24670 23168 24676 23180
rect 23532 23140 24676 23168
rect 23532 23128 23538 23140
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 23566 23060 23572 23112
rect 23624 23060 23630 23112
rect 23658 23060 23664 23112
rect 23716 23100 23722 23112
rect 23845 23103 23903 23109
rect 23845 23100 23857 23103
rect 23716 23072 23857 23100
rect 23716 23060 23722 23072
rect 23845 23069 23857 23072
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 24118 23060 24124 23112
rect 24176 23060 24182 23112
rect 24946 23109 24952 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24940 23100 24952 23109
rect 24907 23072 24952 23100
rect 24581 23063 24639 23069
rect 24940 23063 24952 23072
rect 23106 22992 23112 23044
rect 23164 23032 23170 23044
rect 24596 23032 24624 23063
rect 24946 23060 24952 23063
rect 25004 23060 25010 23112
rect 26252 23109 26280 23276
rect 27154 23264 27160 23276
rect 27212 23264 27218 23316
rect 26513 23239 26571 23245
rect 26513 23205 26525 23239
rect 26559 23236 26571 23239
rect 26970 23236 26976 23248
rect 26559 23208 26976 23236
rect 26559 23205 26571 23208
rect 26513 23199 26571 23205
rect 26970 23196 26976 23208
rect 27028 23196 27034 23248
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 28445 23239 28503 23245
rect 28445 23236 28457 23239
rect 28316 23208 28457 23236
rect 28316 23196 28322 23208
rect 28445 23205 28457 23208
rect 28491 23205 28503 23239
rect 28445 23199 28503 23205
rect 27982 23168 27988 23180
rect 26712 23140 27988 23168
rect 26712 23109 26740 23140
rect 27982 23128 27988 23140
rect 28040 23128 28046 23180
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23069 26295 23103
rect 26237 23063 26295 23069
rect 26697 23103 26755 23109
rect 26697 23069 26709 23103
rect 26743 23069 26755 23103
rect 26697 23063 26755 23069
rect 26973 23103 27031 23109
rect 26973 23069 26985 23103
rect 27019 23100 27031 23103
rect 27019 23072 27108 23100
rect 27019 23069 27031 23072
rect 26973 23063 27031 23069
rect 23164 23004 24624 23032
rect 23164 22992 23170 23004
rect 23385 22967 23443 22973
rect 23385 22964 23397 22967
rect 22572 22936 23397 22964
rect 22373 22927 22431 22933
rect 23385 22933 23397 22936
rect 23431 22933 23443 22967
rect 23385 22927 23443 22933
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 26786 22924 26792 22976
rect 26844 22924 26850 22976
rect 27080 22973 27108 23072
rect 27154 23060 27160 23112
rect 27212 23100 27218 23112
rect 27249 23103 27307 23109
rect 27249 23100 27261 23103
rect 27212 23072 27261 23100
rect 27212 23060 27218 23072
rect 27249 23069 27261 23072
rect 27295 23069 27307 23103
rect 27249 23063 27307 23069
rect 27706 23060 27712 23112
rect 27764 23060 27770 23112
rect 27890 22992 27896 23044
rect 27948 22992 27954 23044
rect 27985 23035 28043 23041
rect 27985 23001 27997 23035
rect 28031 23032 28043 23035
rect 28166 23032 28172 23044
rect 28031 23004 28172 23032
rect 28031 23001 28043 23004
rect 27985 22995 28043 23001
rect 28166 22992 28172 23004
rect 28224 22992 28230 23044
rect 27065 22967 27123 22973
rect 27065 22933 27077 22967
rect 27111 22933 27123 22967
rect 27065 22927 27123 22933
rect 27522 22924 27528 22976
rect 27580 22924 27586 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 2133 22763 2191 22769
rect 2133 22729 2145 22763
rect 2179 22729 2191 22763
rect 2133 22723 2191 22729
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22593 1639 22627
rect 1581 22587 1639 22593
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22624 2099 22627
rect 2148 22624 2176 22723
rect 3326 22720 3332 22772
rect 3384 22720 3390 22772
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4433 22763 4491 22769
rect 4433 22760 4445 22763
rect 4212 22732 4445 22760
rect 4212 22720 4218 22732
rect 4433 22729 4445 22732
rect 4479 22729 4491 22763
rect 4433 22723 4491 22729
rect 5169 22763 5227 22769
rect 5169 22729 5181 22763
rect 5215 22760 5227 22763
rect 5442 22760 5448 22772
rect 5215 22732 5448 22760
rect 5215 22729 5227 22732
rect 5169 22723 5227 22729
rect 5442 22720 5448 22732
rect 5500 22760 5506 22772
rect 6178 22760 6184 22772
rect 5500 22732 6184 22760
rect 5500 22720 5506 22732
rect 6178 22720 6184 22732
rect 6236 22720 6242 22772
rect 6638 22720 6644 22772
rect 6696 22720 6702 22772
rect 7190 22720 7196 22772
rect 7248 22720 7254 22772
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7432 22732 7757 22760
rect 7432 22720 7438 22732
rect 7745 22729 7757 22732
rect 7791 22760 7803 22763
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 7791 22732 8493 22760
rect 7791 22729 7803 22732
rect 7745 22723 7803 22729
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 11882 22760 11888 22772
rect 8481 22723 8539 22729
rect 8588 22732 11888 22760
rect 3234 22692 3240 22704
rect 2332 22664 3240 22692
rect 2332 22633 2360 22664
rect 3234 22652 3240 22664
rect 3292 22652 3298 22704
rect 6656 22692 6684 22720
rect 6822 22692 6828 22704
rect 6196 22664 6828 22692
rect 2087 22596 2176 22624
rect 2317 22627 2375 22633
rect 2087 22593 2099 22596
rect 2041 22587 2099 22593
rect 2317 22593 2329 22627
rect 2363 22593 2375 22627
rect 2317 22587 2375 22593
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22624 2467 22627
rect 2498 22624 2504 22636
rect 2455 22596 2504 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 1596 22488 1624 22587
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 2958 22624 2964 22636
rect 2608 22596 2964 22624
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 2608 22556 2636 22596
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 3602 22584 3608 22636
rect 3660 22584 3666 22636
rect 3789 22627 3847 22633
rect 3789 22593 3801 22627
rect 3835 22624 3847 22627
rect 4338 22624 4344 22636
rect 3835 22596 4344 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 4338 22584 4344 22596
rect 4396 22584 4402 22636
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5166 22624 5172 22636
rect 4755 22596 5172 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5994 22584 6000 22636
rect 6052 22624 6058 22636
rect 6196 22633 6224 22664
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 7009 22695 7067 22701
rect 7009 22661 7021 22695
rect 7055 22661 7067 22695
rect 7208 22692 7236 22720
rect 8588 22692 8616 22732
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 14366 22720 14372 22772
rect 14424 22760 14430 22772
rect 14553 22763 14611 22769
rect 14553 22760 14565 22763
rect 14424 22732 14565 22760
rect 14424 22720 14430 22732
rect 14553 22729 14565 22732
rect 14599 22729 14611 22763
rect 14553 22723 14611 22729
rect 14734 22720 14740 22772
rect 14792 22720 14798 22772
rect 15470 22720 15476 22772
rect 15528 22760 15534 22772
rect 16209 22763 16267 22769
rect 16209 22760 16221 22763
rect 15528 22732 16221 22760
rect 15528 22720 15534 22732
rect 16209 22729 16221 22732
rect 16255 22729 16267 22763
rect 16209 22723 16267 22729
rect 17126 22720 17132 22772
rect 17184 22720 17190 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17865 22763 17923 22769
rect 17865 22760 17877 22763
rect 17276 22732 17877 22760
rect 17276 22720 17282 22732
rect 17865 22729 17877 22732
rect 17911 22729 17923 22763
rect 17865 22723 17923 22729
rect 18506 22720 18512 22772
rect 18564 22720 18570 22772
rect 22554 22760 22560 22772
rect 20180 22732 22560 22760
rect 7208 22664 7328 22692
rect 7009 22655 7067 22661
rect 6181 22627 6239 22633
rect 6181 22624 6193 22627
rect 6052 22596 6193 22624
rect 6052 22584 6058 22596
rect 6181 22593 6193 22596
rect 6227 22593 6239 22627
rect 6181 22587 6239 22593
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6420 22596 6653 22624
rect 6420 22584 6426 22596
rect 6641 22593 6653 22596
rect 6687 22593 6699 22627
rect 7024 22624 7052 22655
rect 7300 22633 7328 22664
rect 8496 22664 8616 22692
rect 7285 22627 7343 22633
rect 7024 22596 7236 22624
rect 6641 22587 6699 22593
rect 1719 22528 2636 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2682 22516 2688 22568
rect 2740 22516 2746 22568
rect 3973 22559 4031 22565
rect 3973 22525 3985 22559
rect 4019 22525 4031 22559
rect 3973 22519 4031 22525
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 4890 22556 4896 22568
rect 4571 22528 4896 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 2406 22488 2412 22500
rect 1596 22460 2412 22488
rect 2406 22448 2412 22460
rect 2464 22448 2470 22500
rect 2501 22491 2559 22497
rect 2501 22457 2513 22491
rect 2547 22488 2559 22491
rect 3988 22488 4016 22519
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 4982 22516 4988 22568
rect 5040 22556 5046 22568
rect 5261 22559 5319 22565
rect 5261 22556 5273 22559
rect 5040 22528 5273 22556
rect 5040 22516 5046 22528
rect 5261 22525 5273 22528
rect 5307 22525 5319 22559
rect 5261 22519 5319 22525
rect 2547 22460 4016 22488
rect 2547 22457 2559 22460
rect 2501 22451 2559 22457
rect 5626 22448 5632 22500
rect 5684 22488 5690 22500
rect 5684 22460 6040 22488
rect 5684 22448 5690 22460
rect 1857 22423 1915 22429
rect 1857 22389 1869 22423
rect 1903 22420 1915 22423
rect 2774 22420 2780 22432
rect 1903 22392 2780 22420
rect 1903 22389 1915 22392
rect 1857 22383 1915 22389
rect 2774 22380 2780 22392
rect 2832 22380 2838 22432
rect 3421 22423 3479 22429
rect 3421 22389 3433 22423
rect 3467 22420 3479 22423
rect 5810 22420 5816 22432
rect 3467 22392 5816 22420
rect 3467 22389 3479 22392
rect 3421 22383 3479 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 5902 22380 5908 22432
rect 5960 22380 5966 22432
rect 6012 22429 6040 22460
rect 5997 22423 6055 22429
rect 5997 22389 6009 22423
rect 6043 22389 6055 22423
rect 6656 22420 6684 22587
rect 7101 22559 7159 22565
rect 7101 22525 7113 22559
rect 7147 22525 7159 22559
rect 7208 22556 7236 22596
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7800 22596 8033 22624
rect 7800 22584 7806 22596
rect 8021 22593 8033 22596
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8496 22624 8524 22664
rect 8662 22652 8668 22704
rect 8720 22692 8726 22704
rect 8757 22695 8815 22701
rect 8757 22692 8769 22695
rect 8720 22664 8769 22692
rect 8720 22652 8726 22664
rect 8757 22661 8769 22664
rect 8803 22661 8815 22695
rect 8757 22655 8815 22661
rect 9582 22652 9588 22704
rect 9640 22652 9646 22704
rect 10413 22695 10471 22701
rect 10413 22661 10425 22695
rect 10459 22692 10471 22695
rect 10870 22692 10876 22704
rect 10459 22664 10876 22692
rect 10459 22661 10471 22664
rect 10413 22655 10471 22661
rect 10870 22652 10876 22664
rect 10928 22652 10934 22704
rect 11698 22652 11704 22704
rect 11756 22652 11762 22704
rect 13256 22695 13314 22701
rect 13256 22661 13268 22695
rect 13302 22692 13314 22695
rect 14752 22692 14780 22720
rect 13302 22664 14780 22692
rect 13302 22661 13314 22664
rect 13256 22655 13314 22661
rect 8168 22596 8524 22624
rect 8168 22584 8174 22596
rect 14182 22584 14188 22636
rect 14240 22624 14246 22636
rect 14461 22627 14519 22633
rect 14461 22624 14473 22627
rect 14240 22596 14473 22624
rect 14240 22584 14246 22596
rect 14461 22593 14473 22596
rect 14507 22593 14519 22627
rect 14461 22587 14519 22593
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 15059 22596 15884 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 7837 22559 7895 22565
rect 7837 22556 7849 22559
rect 7208 22528 7849 22556
rect 7101 22519 7159 22525
rect 7837 22525 7849 22528
rect 7883 22556 7895 22559
rect 8294 22556 8300 22568
rect 7883 22528 8300 22556
rect 7883 22525 7895 22528
rect 7837 22519 7895 22525
rect 7116 22488 7144 22519
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 8665 22559 8723 22565
rect 8665 22556 8677 22559
rect 8404 22528 8677 22556
rect 8404 22488 8432 22528
rect 8665 22525 8677 22528
rect 8711 22556 8723 22559
rect 8711 22528 9168 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 7116 22460 8432 22488
rect 9140 22432 9168 22528
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 9769 22559 9827 22565
rect 9769 22525 9781 22559
rect 9815 22556 9827 22559
rect 10321 22559 10379 22565
rect 10321 22556 10333 22559
rect 9815 22528 10333 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 10321 22525 10333 22528
rect 10367 22525 10379 22559
rect 10321 22519 10379 22525
rect 9217 22491 9275 22497
rect 9217 22457 9229 22491
rect 9263 22488 9275 22491
rect 9784 22488 9812 22519
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 11609 22559 11667 22565
rect 11609 22525 11621 22559
rect 11655 22525 11667 22559
rect 11609 22519 11667 22525
rect 11885 22559 11943 22565
rect 11885 22525 11897 22559
rect 11931 22525 11943 22559
rect 11885 22519 11943 22525
rect 9263 22460 9812 22488
rect 9263 22457 9275 22460
rect 9217 22451 9275 22457
rect 11054 22448 11060 22500
rect 11112 22488 11118 22500
rect 11624 22488 11652 22519
rect 11112 22460 11652 22488
rect 11112 22448 11118 22460
rect 8110 22420 8116 22432
rect 6656 22392 8116 22420
rect 5997 22383 6055 22389
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11900 22420 11928 22519
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12308 22528 13001 22556
rect 12308 22516 12314 22528
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 15105 22559 15163 22565
rect 15105 22525 15117 22559
rect 15151 22556 15163 22559
rect 15194 22556 15200 22568
rect 15151 22528 15200 22556
rect 15151 22525 15163 22528
rect 15105 22519 15163 22525
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 15289 22559 15347 22565
rect 15289 22525 15301 22559
rect 15335 22525 15347 22559
rect 15289 22519 15347 22525
rect 14369 22491 14427 22497
rect 14369 22457 14381 22491
rect 14415 22488 14427 22491
rect 14458 22488 14464 22500
rect 14415 22460 14464 22488
rect 14415 22457 14427 22460
rect 14369 22451 14427 22457
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 14829 22491 14887 22497
rect 14829 22457 14841 22491
rect 14875 22488 14887 22491
rect 15304 22488 15332 22519
rect 15746 22516 15752 22568
rect 15804 22516 15810 22568
rect 15856 22497 15884 22596
rect 16022 22584 16028 22636
rect 16080 22584 16086 22636
rect 16117 22627 16175 22633
rect 16117 22593 16129 22627
rect 16163 22624 16175 22627
rect 16298 22624 16304 22636
rect 16163 22596 16304 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 17144 22633 17172 22720
rect 18524 22692 18552 22720
rect 19061 22695 19119 22701
rect 19061 22692 19073 22695
rect 18524 22664 19073 22692
rect 19061 22661 19073 22664
rect 19107 22661 19119 22695
rect 19061 22655 19119 22661
rect 19886 22652 19892 22704
rect 19944 22652 19950 22704
rect 20180 22633 20208 22732
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23624 22732 23765 22760
rect 23624 22720 23630 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 23753 22723 23811 22729
rect 24118 22720 24124 22772
rect 24176 22760 24182 22772
rect 24305 22763 24363 22769
rect 24305 22760 24317 22763
rect 24176 22732 24317 22760
rect 24176 22720 24182 22732
rect 24305 22729 24317 22732
rect 24351 22729 24363 22763
rect 24305 22723 24363 22729
rect 24854 22720 24860 22772
rect 24912 22720 24918 22772
rect 26050 22720 26056 22772
rect 26108 22720 26114 22772
rect 26326 22720 26332 22772
rect 26384 22720 26390 22772
rect 26786 22720 26792 22772
rect 26844 22760 26850 22772
rect 27801 22763 27859 22769
rect 26844 22732 27476 22760
rect 26844 22720 26850 22732
rect 22741 22695 22799 22701
rect 22741 22692 22753 22695
rect 20364 22664 22753 22692
rect 20364 22633 20392 22664
rect 22741 22661 22753 22664
rect 22787 22661 22799 22695
rect 24872 22692 24900 22720
rect 22741 22655 22799 22661
rect 23400 22664 23980 22692
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 17175 22596 17785 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17773 22593 17785 22596
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20772 22596 20913 22624
rect 20772 22584 20778 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 21545 22627 21603 22633
rect 21545 22624 21557 22627
rect 21140 22596 21557 22624
rect 21140 22584 21146 22596
rect 21545 22593 21557 22596
rect 21591 22593 21603 22627
rect 21545 22587 21603 22593
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 16040 22556 16068 22584
rect 17586 22556 17592 22568
rect 16040 22528 17592 22556
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 18138 22516 18144 22568
rect 18196 22516 18202 22568
rect 18322 22516 18328 22568
rect 18380 22516 18386 22568
rect 18969 22559 19027 22565
rect 18969 22556 18981 22559
rect 18892 22528 18981 22556
rect 14875 22460 15332 22488
rect 15841 22491 15899 22497
rect 14875 22457 14887 22460
rect 14829 22451 14887 22457
rect 15841 22457 15853 22491
rect 15887 22457 15899 22491
rect 15841 22451 15899 22457
rect 11296 22392 11928 22420
rect 11296 22380 11302 22392
rect 17678 22380 17684 22432
rect 17736 22380 17742 22432
rect 18785 22423 18843 22429
rect 18785 22389 18797 22423
rect 18831 22420 18843 22423
rect 18892 22420 18920 22528
rect 18969 22525 18981 22528
rect 19015 22525 19027 22559
rect 18969 22519 19027 22525
rect 19334 22516 19340 22568
rect 19392 22516 19398 22568
rect 20806 22516 20812 22568
rect 20864 22516 20870 22568
rect 21836 22556 21864 22587
rect 22002 22584 22008 22636
rect 22060 22624 22066 22636
rect 22278 22624 22284 22636
rect 22060 22596 22284 22624
rect 22060 22584 22066 22596
rect 22278 22584 22284 22596
rect 22336 22624 22342 22636
rect 23400 22633 23428 22664
rect 23952 22633 23980 22664
rect 24872 22664 26004 22692
rect 22557 22627 22615 22633
rect 22557 22624 22569 22627
rect 22336 22596 22569 22624
rect 22336 22584 22342 22596
rect 22557 22593 22569 22596
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 22925 22627 22983 22633
rect 22925 22624 22937 22627
rect 22695 22596 22937 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 22925 22593 22937 22596
rect 22971 22593 22983 22627
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 22925 22587 22983 22593
rect 23023 22596 23397 22624
rect 21008 22528 21864 22556
rect 20073 22491 20131 22497
rect 20073 22457 20085 22491
rect 20119 22488 20131 22491
rect 20438 22488 20444 22500
rect 20119 22460 20444 22488
rect 20119 22457 20131 22460
rect 20073 22451 20131 22457
rect 20438 22448 20444 22460
rect 20496 22448 20502 22500
rect 20530 22448 20536 22500
rect 20588 22488 20594 22500
rect 21008 22488 21036 22528
rect 22370 22516 22376 22568
rect 22428 22556 22434 22568
rect 22664 22556 22692 22587
rect 22428 22528 22692 22556
rect 22428 22516 22434 22528
rect 20588 22460 21036 22488
rect 20588 22448 20594 22460
rect 21910 22448 21916 22500
rect 21968 22448 21974 22500
rect 22002 22448 22008 22500
rect 22060 22488 22066 22500
rect 22097 22491 22155 22497
rect 22097 22488 22109 22491
rect 22060 22460 22109 22488
rect 22060 22448 22066 22460
rect 22097 22457 22109 22460
rect 22143 22457 22155 22491
rect 22097 22451 22155 22457
rect 22462 22448 22468 22500
rect 22520 22488 22526 22500
rect 23023 22488 23051 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 23676 22556 23704 22587
rect 24026 22584 24032 22636
rect 24084 22624 24090 22636
rect 24489 22627 24547 22633
rect 24084 22596 24440 22624
rect 24084 22584 24090 22596
rect 23216 22528 23704 22556
rect 24412 22556 24440 22596
rect 24489 22593 24501 22627
rect 24535 22624 24547 22627
rect 24765 22627 24823 22633
rect 24765 22624 24777 22627
rect 24535 22596 24777 22624
rect 24535 22593 24547 22596
rect 24489 22587 24547 22593
rect 24765 22593 24777 22596
rect 24811 22624 24823 22627
rect 24872 22624 24900 22664
rect 24811 22596 24900 22624
rect 25501 22627 25559 22633
rect 24811 22593 24823 22596
rect 24765 22587 24823 22593
rect 25501 22593 25513 22627
rect 25547 22624 25559 22627
rect 25590 22624 25596 22636
rect 25547 22596 25596 22624
rect 25547 22593 25559 22596
rect 25501 22587 25559 22593
rect 25041 22559 25099 22565
rect 25041 22556 25053 22559
rect 24412 22528 25053 22556
rect 23216 22497 23244 22528
rect 25041 22525 25053 22528
rect 25087 22556 25099 22559
rect 25516 22556 25544 22587
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 25976 22633 26004 22664
rect 25961 22627 26019 22633
rect 25961 22593 25973 22627
rect 26007 22593 26019 22627
rect 26068 22624 26096 22720
rect 26344 22692 26372 22720
rect 26344 22664 27384 22692
rect 26237 22627 26295 22633
rect 26237 22624 26249 22627
rect 26068 22596 26249 22624
rect 25961 22587 26019 22593
rect 26237 22593 26249 22596
rect 26283 22624 26295 22627
rect 26329 22627 26387 22633
rect 26329 22624 26341 22627
rect 26283 22596 26341 22624
rect 26283 22593 26295 22596
rect 26237 22587 26295 22593
rect 26329 22593 26341 22596
rect 26375 22624 26387 22627
rect 26602 22624 26608 22636
rect 26375 22596 26608 22624
rect 26375 22593 26387 22596
rect 26329 22587 26387 22593
rect 26602 22584 26608 22596
rect 26660 22624 26666 22636
rect 27356 22633 27384 22664
rect 26789 22627 26847 22633
rect 26789 22624 26801 22627
rect 26660 22596 26801 22624
rect 26660 22584 26666 22596
rect 26789 22593 26801 22596
rect 26835 22593 26847 22627
rect 26789 22587 26847 22593
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22593 27399 22627
rect 27448 22624 27476 22732
rect 27801 22729 27813 22763
rect 27847 22760 27859 22763
rect 27890 22760 27896 22772
rect 27847 22732 27896 22760
rect 27847 22729 27859 22732
rect 27801 22723 27859 22729
rect 27890 22720 27896 22732
rect 27948 22760 27954 22772
rect 28537 22763 28595 22769
rect 28537 22760 28549 22763
rect 27948 22732 28549 22760
rect 27948 22720 27954 22732
rect 28537 22729 28549 22732
rect 28583 22729 28595 22763
rect 28537 22723 28595 22729
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 27448 22596 28089 22624
rect 27341 22587 27399 22593
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 25087 22528 25544 22556
rect 27157 22559 27215 22565
rect 25087 22525 25099 22528
rect 25041 22519 25099 22525
rect 27157 22525 27169 22559
rect 27203 22525 27215 22559
rect 27157 22519 27215 22525
rect 22520 22460 23051 22488
rect 23201 22491 23259 22497
rect 22520 22448 22526 22460
rect 23201 22457 23213 22491
rect 23247 22457 23259 22491
rect 23201 22451 23259 22457
rect 26234 22448 26240 22500
rect 26292 22488 26298 22500
rect 27172 22488 27200 22519
rect 27706 22516 27712 22568
rect 27764 22516 27770 22568
rect 27890 22516 27896 22568
rect 27948 22516 27954 22568
rect 26292 22460 27200 22488
rect 26292 22448 26298 22460
rect 19610 22420 19616 22432
rect 18831 22392 19616 22420
rect 18831 22389 18843 22392
rect 18785 22383 18843 22389
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 22373 22423 22431 22429
rect 22373 22420 22385 22423
rect 22244 22392 22385 22420
rect 22244 22380 22250 22392
rect 22373 22389 22385 22392
rect 22419 22389 22431 22423
rect 22373 22383 22431 22389
rect 23014 22380 23020 22432
rect 23072 22380 23078 22432
rect 23474 22380 23480 22432
rect 23532 22380 23538 22432
rect 24118 22380 24124 22432
rect 24176 22380 24182 22432
rect 24762 22380 24768 22432
rect 24820 22420 24826 22432
rect 25593 22423 25651 22429
rect 25593 22420 25605 22423
rect 24820 22392 25605 22420
rect 24820 22380 24826 22392
rect 25593 22389 25605 22392
rect 25639 22389 25651 22423
rect 25593 22383 25651 22389
rect 25774 22380 25780 22432
rect 25832 22380 25838 22432
rect 26053 22423 26111 22429
rect 26053 22389 26065 22423
rect 26099 22420 26111 22423
rect 26326 22420 26332 22432
rect 26099 22392 26332 22420
rect 26099 22389 26111 22392
rect 26053 22383 26111 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 26418 22380 26424 22432
rect 26476 22380 26482 22432
rect 26605 22423 26663 22429
rect 26605 22389 26617 22423
rect 26651 22420 26663 22423
rect 27724 22420 27752 22516
rect 26651 22392 27752 22420
rect 26651 22389 26663 22392
rect 26605 22383 26663 22389
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 2682 22176 2688 22228
rect 2740 22216 2746 22228
rect 2777 22219 2835 22225
rect 2777 22216 2789 22219
rect 2740 22188 2789 22216
rect 2740 22176 2746 22188
rect 2777 22185 2789 22188
rect 2823 22185 2835 22219
rect 2777 22179 2835 22185
rect 3421 22219 3479 22225
rect 3421 22185 3433 22219
rect 3467 22216 3479 22219
rect 3602 22216 3608 22228
rect 3467 22188 3608 22216
rect 3467 22185 3479 22188
rect 3421 22179 3479 22185
rect 3602 22176 3608 22188
rect 3660 22176 3666 22228
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 5408 22188 6132 22216
rect 5408 22176 5414 22188
rect 2498 22108 2504 22160
rect 2556 22148 2562 22160
rect 3326 22148 3332 22160
rect 2556 22120 3332 22148
rect 2556 22108 2562 22120
rect 3326 22108 3332 22120
rect 3384 22108 3390 22160
rect 5994 22148 6000 22160
rect 5092 22120 6000 22148
rect 1394 22040 1400 22092
rect 1452 22040 1458 22092
rect 3068 22052 3464 22080
rect 3068 22021 3096 22052
rect 3436 22024 3464 22052
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 3973 22083 4031 22089
rect 3973 22080 3985 22083
rect 3752 22052 3985 22080
rect 3752 22040 3758 22052
rect 3973 22049 3985 22052
rect 4019 22049 4031 22083
rect 5092 22080 5120 22120
rect 5994 22108 6000 22120
rect 6052 22108 6058 22160
rect 6104 22148 6132 22188
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6365 22219 6423 22225
rect 6365 22216 6377 22219
rect 6236 22188 6377 22216
rect 6236 22176 6242 22188
rect 6365 22185 6377 22188
rect 6411 22185 6423 22219
rect 6365 22179 6423 22185
rect 7377 22219 7435 22225
rect 7377 22185 7389 22219
rect 7423 22216 7435 22219
rect 7466 22216 7472 22228
rect 7423 22188 7472 22216
rect 7423 22185 7435 22188
rect 7377 22179 7435 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 7558 22176 7564 22228
rect 7616 22216 7622 22228
rect 9582 22216 9588 22228
rect 7616 22188 9588 22216
rect 7616 22176 7622 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 11698 22176 11704 22228
rect 11756 22176 11762 22228
rect 14090 22176 14096 22228
rect 14148 22176 14154 22228
rect 14737 22219 14795 22225
rect 14737 22185 14749 22219
rect 14783 22216 14795 22219
rect 15102 22216 15108 22228
rect 14783 22188 15108 22216
rect 14783 22185 14795 22188
rect 14737 22179 14795 22185
rect 15102 22176 15108 22188
rect 15160 22176 15166 22228
rect 16298 22176 16304 22228
rect 16356 22216 16362 22228
rect 16356 22188 17540 22216
rect 16356 22176 16362 22188
rect 9858 22148 9864 22160
rect 6104 22120 9864 22148
rect 9858 22108 9864 22120
rect 9916 22108 9922 22160
rect 10134 22108 10140 22160
rect 10192 22108 10198 22160
rect 11517 22151 11575 22157
rect 11517 22148 11529 22151
rect 10428 22120 11529 22148
rect 3973 22043 4031 22049
rect 4080 22052 5120 22080
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 21981 3111 22015
rect 3053 21975 3111 21981
rect 3142 21972 3148 22024
rect 3200 21972 3206 22024
rect 3418 21972 3424 22024
rect 3476 21972 3482 22024
rect 3605 22015 3663 22021
rect 3605 21981 3617 22015
rect 3651 22012 3663 22015
rect 4080 22012 4108 22052
rect 5258 22040 5264 22092
rect 5316 22040 5322 22092
rect 8110 22040 8116 22092
rect 8168 22040 8174 22092
rect 8386 22040 8392 22092
rect 8444 22080 8450 22092
rect 8662 22080 8668 22092
rect 8444 22052 8668 22080
rect 8444 22040 8450 22052
rect 8662 22040 8668 22052
rect 8720 22040 8726 22092
rect 8846 22040 8852 22092
rect 8904 22080 8910 22092
rect 9309 22083 9367 22089
rect 9309 22080 9321 22083
rect 8904 22052 9321 22080
rect 8904 22040 8910 22052
rect 9309 22049 9321 22052
rect 9355 22049 9367 22083
rect 10152 22080 10180 22108
rect 10428 22089 10456 22120
rect 11517 22117 11529 22120
rect 11563 22117 11575 22151
rect 11517 22111 11575 22117
rect 13633 22151 13691 22157
rect 13633 22117 13645 22151
rect 13679 22148 13691 22151
rect 14108 22148 14136 22176
rect 13679 22120 14136 22148
rect 13679 22117 13691 22120
rect 13633 22111 13691 22117
rect 10413 22083 10471 22089
rect 10413 22080 10425 22083
rect 10152 22052 10425 22080
rect 9309 22043 9367 22049
rect 10413 22049 10425 22052
rect 10459 22049 10471 22083
rect 10413 22043 10471 22049
rect 10962 22040 10968 22092
rect 11020 22080 11026 22092
rect 12250 22080 12256 22092
rect 11020 22052 12256 22080
rect 11020 22040 11026 22052
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 13832 22080 13860 22120
rect 13740 22052 13860 22080
rect 14277 22083 14335 22089
rect 3651 21984 4108 22012
rect 4157 22015 4215 22021
rect 3651 21981 3663 21984
rect 3605 21975 3663 21981
rect 4157 21981 4169 22015
rect 4203 22012 4215 22015
rect 4338 22012 4344 22024
rect 4203 21984 4344 22012
rect 4203 21981 4215 21984
rect 4157 21975 4215 21981
rect 4338 21972 4344 21984
rect 4396 21972 4402 22024
rect 4890 21972 4896 22024
rect 4948 21972 4954 22024
rect 5166 21972 5172 22024
rect 5224 21972 5230 22024
rect 5445 22015 5503 22021
rect 5445 22014 5457 22015
rect 5368 22012 5457 22014
rect 5276 21986 5457 22012
rect 5276 21984 5396 21986
rect 1664 21947 1722 21953
rect 1664 21913 1676 21947
rect 1710 21944 1722 21947
rect 2222 21944 2228 21956
rect 1710 21916 2228 21944
rect 1710 21913 1722 21916
rect 1664 21907 1722 21913
rect 2222 21904 2228 21916
rect 2280 21904 2286 21956
rect 3237 21947 3295 21953
rect 3237 21913 3249 21947
rect 3283 21944 3295 21947
rect 5276 21944 5304 21984
rect 5445 21981 5457 21986
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 5905 22015 5963 22021
rect 5905 22012 5917 22015
rect 5592 21984 5917 22012
rect 5592 21972 5598 21984
rect 5905 21981 5917 21984
rect 5951 21981 5963 22015
rect 5905 21975 5963 21981
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 22014 6239 22015
rect 6227 21986 6316 22014
rect 6227 21981 6239 21986
rect 6181 21975 6239 21981
rect 3283 21916 5304 21944
rect 3283 21913 3295 21916
rect 3237 21907 3295 21913
rect 2869 21879 2927 21885
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 4062 21876 4068 21888
rect 2915 21848 4068 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 4062 21836 4068 21848
rect 4120 21836 4126 21888
rect 4614 21836 4620 21888
rect 4672 21836 4678 21888
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 4985 21879 5043 21885
rect 4985 21845 4997 21879
rect 5031 21876 5043 21879
rect 5718 21876 5724 21888
rect 5031 21848 5724 21876
rect 5031 21845 5043 21848
rect 4985 21839 5043 21845
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 5810 21836 5816 21888
rect 5868 21876 5874 21888
rect 6288 21876 6316 21986
rect 6822 21972 6828 22024
rect 6880 21972 6886 22024
rect 7650 21972 7656 22024
rect 7708 21972 7714 22024
rect 8021 22015 8079 22021
rect 8021 21981 8033 22015
rect 8067 22012 8079 22015
rect 8481 22015 8539 22021
rect 8067 21984 8432 22012
rect 8067 21981 8079 21984
rect 8021 21975 8079 21981
rect 8404 21944 8432 21984
rect 8481 21981 8493 22015
rect 8527 22012 8539 22015
rect 8754 22012 8760 22024
rect 8527 21984 8760 22012
rect 8527 21981 8539 21984
rect 8481 21975 8539 21981
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 9140 21944 9168 21975
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12802 22012 12808 22024
rect 12207 21984 12808 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 13740 22021 13768 22052
rect 14277 22049 14289 22083
rect 14323 22080 14335 22083
rect 14921 22083 14979 22089
rect 14921 22080 14933 22083
rect 14323 22052 14933 22080
rect 14323 22049 14335 22052
rect 14277 22043 14335 22049
rect 14921 22049 14933 22052
rect 14967 22049 14979 22083
rect 16500 22080 16528 22188
rect 17512 22148 17540 22188
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18969 22219 19027 22225
rect 18969 22216 18981 22219
rect 18196 22188 18981 22216
rect 18196 22176 18202 22188
rect 18969 22185 18981 22188
rect 19015 22185 19027 22219
rect 18969 22179 19027 22185
rect 19610 22176 19616 22228
rect 19668 22176 19674 22228
rect 20530 22216 20536 22228
rect 20364 22188 20536 22216
rect 20364 22148 20392 22188
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 21269 22219 21327 22225
rect 21269 22216 21281 22219
rect 20864 22188 21281 22216
rect 20864 22176 20870 22188
rect 21269 22185 21281 22188
rect 21315 22185 21327 22219
rect 21269 22179 21327 22185
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 23808 22188 27384 22216
rect 23808 22176 23814 22188
rect 25041 22151 25099 22157
rect 17512 22120 20392 22148
rect 20456 22120 20944 22148
rect 20456 22092 20484 22120
rect 19245 22083 19303 22089
rect 14921 22043 14979 22049
rect 15304 22052 16565 22080
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 13817 22015 13875 22021
rect 13817 21981 13829 22015
rect 13863 22012 13875 22015
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13863 21984 14105 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14829 22015 14887 22021
rect 14829 21981 14841 22015
rect 14875 22012 14887 22015
rect 15304 22012 15332 22052
rect 14875 21984 15332 22012
rect 15381 22015 15439 22021
rect 14875 21981 14887 21984
rect 14829 21975 14887 21981
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 16298 22012 16304 22024
rect 15427 21984 16304 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16500 22021 16528 22052
rect 19245 22049 19257 22083
rect 19291 22080 19303 22083
rect 20073 22083 20131 22089
rect 20073 22080 20085 22083
rect 19291 22052 20085 22080
rect 19291 22049 19303 22052
rect 19245 22043 19303 22049
rect 20073 22049 20085 22052
rect 20119 22049 20131 22083
rect 20073 22043 20131 22049
rect 20438 22040 20444 22092
rect 20496 22040 20502 22092
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16574 21972 16580 22024
rect 16632 21972 16638 22024
rect 16844 22015 16902 22021
rect 16844 21981 16856 22015
rect 16890 22012 16902 22015
rect 17678 22012 17684 22024
rect 16890 21984 17684 22012
rect 16890 21981 16902 21984
rect 16844 21975 16902 21981
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 22012 18199 22015
rect 18877 22015 18935 22021
rect 18877 22012 18889 22015
rect 18187 21984 18889 22012
rect 18187 21981 18199 21984
rect 18141 21975 18199 21981
rect 18877 21981 18889 21984
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 19886 22012 19892 22024
rect 19475 21984 19892 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 6564 21916 8340 21944
rect 8404 21916 8524 21944
rect 6564 21888 6592 21916
rect 5868 21848 6316 21876
rect 5868 21836 5874 21848
rect 6546 21836 6552 21888
rect 6604 21836 6610 21888
rect 7742 21836 7748 21888
rect 7800 21836 7806 21888
rect 8312 21885 8340 21916
rect 8496 21888 8524 21916
rect 8588 21916 9168 21944
rect 9401 21947 9459 21953
rect 8297 21879 8355 21885
rect 8297 21845 8309 21879
rect 8343 21845 8355 21879
rect 8297 21839 8355 21845
rect 8478 21836 8484 21888
rect 8536 21836 8542 21888
rect 8588 21885 8616 21916
rect 9401 21913 9413 21947
rect 9447 21944 9459 21947
rect 9674 21944 9680 21956
rect 9447 21916 9680 21944
rect 9447 21913 9459 21916
rect 9401 21907 9459 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 9950 21904 9956 21956
rect 10008 21904 10014 21956
rect 10134 21904 10140 21956
rect 10192 21904 10198 21956
rect 10229 21947 10287 21953
rect 10229 21913 10241 21947
rect 10275 21913 10287 21947
rect 10229 21907 10287 21913
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 8938 21836 8944 21888
rect 8996 21836 9002 21888
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10244 21876 10272 21907
rect 10410 21904 10416 21956
rect 10468 21944 10474 21956
rect 10965 21947 11023 21953
rect 10965 21944 10977 21947
rect 10468 21916 10977 21944
rect 10468 21904 10474 21916
rect 10965 21913 10977 21916
rect 11011 21913 11023 21947
rect 10965 21907 11023 21913
rect 11057 21947 11115 21953
rect 11057 21913 11069 21947
rect 11103 21913 11115 21947
rect 11057 21907 11115 21913
rect 12520 21947 12578 21953
rect 12520 21913 12532 21947
rect 12566 21944 12578 21947
rect 13262 21944 13268 21956
rect 12566 21916 13268 21944
rect 12566 21913 12578 21916
rect 12520 21907 12578 21913
rect 9824 21848 10272 21876
rect 9824 21836 9830 21848
rect 10318 21836 10324 21888
rect 10376 21876 10382 21888
rect 11072 21876 11100 21907
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 15562 21904 15568 21956
rect 15620 21944 15626 21956
rect 15749 21947 15807 21953
rect 15749 21944 15761 21947
rect 15620 21916 15761 21944
rect 15620 21904 15626 21916
rect 15749 21913 15761 21916
rect 15795 21913 15807 21947
rect 15749 21907 15807 21913
rect 10376 21848 11100 21876
rect 11977 21879 12035 21885
rect 10376 21836 10382 21848
rect 11977 21845 11989 21879
rect 12023 21876 12035 21879
rect 13906 21876 13912 21888
rect 12023 21848 13912 21876
rect 12023 21845 12035 21848
rect 11977 21839 12035 21845
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 16301 21879 16359 21885
rect 16301 21845 16313 21879
rect 16347 21876 16359 21879
rect 17494 21876 17500 21888
rect 16347 21848 17500 21876
rect 16347 21845 16359 21848
rect 16301 21839 16359 21845
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17957 21879 18015 21885
rect 17957 21845 17969 21879
rect 18003 21876 18015 21879
rect 18156 21876 18184 21975
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 19978 21972 19984 22024
rect 20036 21972 20042 22024
rect 20916 22021 20944 22120
rect 25041 22117 25053 22151
rect 25087 22148 25099 22151
rect 25498 22148 25504 22160
rect 25087 22120 25504 22148
rect 25087 22117 25099 22120
rect 25041 22111 25099 22117
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 21542 22040 21548 22092
rect 21600 22080 21606 22092
rect 21821 22083 21879 22089
rect 21821 22080 21833 22083
rect 21600 22052 21833 22080
rect 21600 22040 21606 22052
rect 21821 22049 21833 22052
rect 21867 22049 21879 22083
rect 21821 22043 21879 22049
rect 22557 22083 22615 22089
rect 22557 22049 22569 22083
rect 22603 22080 22615 22083
rect 22603 22052 23244 22080
rect 22603 22049 22615 22052
rect 22557 22043 22615 22049
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 20349 21947 20407 21953
rect 20349 21913 20361 21947
rect 20395 21913 20407 21947
rect 20349 21907 20407 21913
rect 18003 21848 18184 21876
rect 18003 21845 18015 21848
rect 17957 21839 18015 21845
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 20364 21876 20392 21907
rect 18840 21848 20392 21876
rect 20441 21879 20499 21885
rect 18840 21836 18846 21848
rect 20441 21845 20453 21879
rect 20487 21876 20499 21879
rect 20530 21876 20536 21888
rect 20487 21848 20536 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20622 21836 20628 21888
rect 20680 21836 20686 21888
rect 20824 21876 20852 21975
rect 20916 21944 20944 21975
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 21358 21972 21364 22024
rect 21416 22012 21422 22024
rect 21637 22015 21695 22021
rect 21637 22012 21649 22015
rect 21416 21984 21649 22012
rect 21416 21972 21422 21984
rect 21637 21981 21649 21984
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22336 21984 22385 22012
rect 22336 21972 22342 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 21981 23167 22015
rect 23216 22012 23244 22052
rect 23290 22040 23296 22092
rect 23348 22040 23354 22092
rect 24581 22083 24639 22089
rect 24581 22049 24593 22083
rect 24627 22080 24639 22083
rect 24762 22080 24768 22092
rect 24627 22052 24768 22080
rect 24627 22049 24639 22052
rect 24581 22043 24639 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 24946 22040 24952 22092
rect 25004 22080 25010 22092
rect 25869 22083 25927 22089
rect 25869 22080 25881 22083
rect 25004 22052 25881 22080
rect 25004 22040 25010 22052
rect 25869 22049 25881 22052
rect 25915 22049 25927 22083
rect 25869 22043 25927 22049
rect 26053 22083 26111 22089
rect 26053 22049 26065 22083
rect 26099 22080 26111 22083
rect 26418 22080 26424 22092
rect 26099 22052 26424 22080
rect 26099 22049 26111 22052
rect 26053 22043 26111 22049
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 27356 22089 27384 22188
rect 27341 22083 27399 22089
rect 27341 22049 27353 22083
rect 27387 22049 27399 22083
rect 27341 22043 27399 22049
rect 27522 22040 27528 22092
rect 27580 22040 27586 22092
rect 23474 22012 23480 22024
rect 23216 21984 23480 22012
rect 23109 21975 23167 21981
rect 23124 21944 23152 21975
rect 23474 21972 23480 21984
rect 23532 21972 23538 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 22012 23903 22015
rect 24026 22012 24032 22024
rect 23891 21984 24032 22012
rect 23891 21981 23903 21984
rect 23845 21975 23903 21981
rect 24026 21972 24032 21984
rect 24084 21972 24090 22024
rect 24394 21972 24400 22024
rect 24452 21972 24458 22024
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25314 21972 25320 22024
rect 25372 21972 25378 22024
rect 26605 22015 26663 22021
rect 26605 21981 26617 22015
rect 26651 21981 26663 22015
rect 26605 21975 26663 21981
rect 20916 21916 23152 21944
rect 25498 21904 25504 21956
rect 25556 21944 25562 21956
rect 26620 21944 26648 21975
rect 26786 21972 26792 22024
rect 26844 21972 26850 22024
rect 27430 21972 27436 22024
rect 27488 22012 27494 22024
rect 28261 22015 28319 22021
rect 28261 22012 28273 22015
rect 27488 21984 28273 22012
rect 27488 21972 27494 21984
rect 28261 21981 28273 21984
rect 28307 21981 28319 22015
rect 28261 21975 28319 21981
rect 25556 21916 26648 21944
rect 27249 21947 27307 21953
rect 25556 21904 25562 21916
rect 27249 21913 27261 21947
rect 27295 21944 27307 21947
rect 27890 21944 27896 21956
rect 27295 21916 27896 21944
rect 27295 21913 27307 21916
rect 27249 21907 27307 21913
rect 27890 21904 27896 21916
rect 27948 21944 27954 21956
rect 27985 21947 28043 21953
rect 27985 21944 27997 21947
rect 27948 21916 27997 21944
rect 27948 21904 27954 21916
rect 27985 21913 27997 21916
rect 28031 21913 28043 21947
rect 27985 21907 28043 21913
rect 22186 21876 22192 21888
rect 20824 21848 22192 21876
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21876 22339 21879
rect 22646 21876 22652 21888
rect 22327 21848 22652 21876
rect 22327 21845 22339 21848
rect 22281 21839 22339 21845
rect 22646 21836 22652 21848
rect 22704 21876 22710 21888
rect 23017 21879 23075 21885
rect 23017 21876 23029 21879
rect 22704 21848 23029 21876
rect 22704 21836 22710 21848
rect 23017 21845 23029 21848
rect 23063 21845 23075 21879
rect 23017 21839 23075 21845
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 23937 21879 23995 21885
rect 23937 21876 23949 21879
rect 23440 21848 23949 21876
rect 23440 21836 23446 21848
rect 23937 21845 23949 21848
rect 23983 21845 23995 21879
rect 23937 21839 23995 21845
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 26513 21879 26571 21885
rect 26513 21876 26525 21879
rect 26292 21848 26525 21876
rect 26292 21836 26298 21848
rect 26513 21845 26525 21848
rect 26559 21845 26571 21879
rect 26513 21839 26571 21845
rect 28074 21836 28080 21888
rect 28132 21836 28138 21888
rect 28350 21836 28356 21888
rect 28408 21836 28414 21888
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 2222 21632 2228 21684
rect 2280 21632 2286 21684
rect 2682 21632 2688 21684
rect 2740 21632 2746 21684
rect 4614 21632 4620 21684
rect 4672 21672 4678 21684
rect 4798 21672 4804 21684
rect 4672 21644 4804 21672
rect 4672 21632 4678 21644
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 6181 21675 6239 21681
rect 6181 21672 6193 21675
rect 5592 21644 6193 21672
rect 5592 21632 5598 21644
rect 6181 21641 6193 21644
rect 6227 21641 6239 21675
rect 6181 21635 6239 21641
rect 6365 21675 6423 21681
rect 6365 21641 6377 21675
rect 6411 21672 6423 21675
rect 7558 21672 7564 21684
rect 6411 21644 7564 21672
rect 6411 21641 6423 21644
rect 6365 21635 6423 21641
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 9582 21672 9588 21684
rect 8536 21644 9588 21672
rect 8536 21632 8542 21644
rect 9582 21632 9588 21644
rect 9640 21632 9646 21684
rect 9950 21632 9956 21684
rect 10008 21672 10014 21684
rect 11054 21672 11060 21684
rect 10008 21644 11060 21672
rect 10008 21632 10014 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21672 13875 21675
rect 14274 21672 14280 21684
rect 13863 21644 14280 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 15381 21675 15439 21681
rect 15381 21641 15393 21675
rect 15427 21672 15439 21675
rect 17313 21675 17371 21681
rect 15427 21644 15608 21672
rect 15427 21641 15439 21644
rect 15381 21635 15439 21641
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 2038 21496 2044 21548
rect 2096 21496 2102 21548
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 2700 21536 2728 21632
rect 4706 21564 4712 21616
rect 4764 21604 4770 21616
rect 4764 21576 5672 21604
rect 4764 21564 4770 21576
rect 2363 21508 2728 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 2958 21496 2964 21548
rect 3016 21536 3022 21548
rect 3513 21539 3571 21545
rect 3513 21536 3525 21539
rect 3016 21508 3525 21536
rect 3016 21496 3022 21508
rect 3513 21505 3525 21508
rect 3559 21505 3571 21539
rect 3513 21499 3571 21505
rect 4154 21496 4160 21548
rect 4212 21496 4218 21548
rect 4890 21496 4896 21548
rect 4948 21496 4954 21548
rect 4982 21496 4988 21548
rect 5040 21536 5046 21548
rect 5077 21539 5135 21545
rect 5077 21536 5089 21539
rect 5040 21508 5089 21536
rect 5040 21496 5046 21508
rect 5077 21505 5089 21508
rect 5123 21536 5135 21539
rect 5350 21536 5356 21548
rect 5123 21508 5356 21536
rect 5123 21505 5135 21508
rect 5077 21499 5135 21505
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 5445 21539 5503 21545
rect 5445 21505 5457 21539
rect 5491 21536 5503 21539
rect 5491 21508 5580 21536
rect 5491 21505 5503 21508
rect 5445 21499 5503 21505
rect 2056 21468 2084 21496
rect 2593 21471 2651 21477
rect 2593 21468 2605 21471
rect 2056 21440 2605 21468
rect 2593 21437 2605 21440
rect 2639 21437 2651 21471
rect 3329 21471 3387 21477
rect 3329 21468 3341 21471
rect 2593 21431 2651 21437
rect 2746 21440 3341 21468
rect 2409 21403 2467 21409
rect 2409 21369 2421 21403
rect 2455 21400 2467 21403
rect 2746 21400 2774 21440
rect 3329 21437 3341 21440
rect 3375 21437 3387 21471
rect 3329 21431 3387 21437
rect 3878 21428 3884 21480
rect 3936 21468 3942 21480
rect 4341 21471 4399 21477
rect 4341 21468 4353 21471
rect 3936 21440 4353 21468
rect 3936 21428 3942 21440
rect 4341 21437 4353 21440
rect 4387 21437 4399 21471
rect 4341 21431 4399 21437
rect 2455 21372 2774 21400
rect 4908 21400 4936 21496
rect 5552 21480 5580 21508
rect 5258 21428 5264 21480
rect 5316 21468 5322 21480
rect 5534 21468 5540 21480
rect 5316 21440 5540 21468
rect 5316 21428 5322 21440
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 5644 21468 5672 21576
rect 7006 21564 7012 21616
rect 7064 21604 7070 21616
rect 7101 21607 7159 21613
rect 7101 21604 7113 21607
rect 7064 21576 7113 21604
rect 7064 21564 7070 21576
rect 7101 21573 7113 21576
rect 7147 21573 7159 21607
rect 7101 21567 7159 21573
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 7708 21576 8800 21604
rect 7708 21564 7714 21576
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 6822 21536 6828 21548
rect 6779 21508 6828 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 7852 21545 7880 21576
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8772 21536 8800 21576
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 10781 21607 10839 21613
rect 10781 21604 10793 21607
rect 8996 21576 10793 21604
rect 8996 21564 9002 21576
rect 10781 21573 10793 21576
rect 10827 21573 10839 21607
rect 10781 21567 10839 21573
rect 12520 21607 12578 21613
rect 12520 21573 12532 21607
rect 12566 21604 12578 21607
rect 12894 21604 12900 21616
rect 12566 21576 12900 21604
rect 12566 21573 12578 21576
rect 12520 21567 12578 21573
rect 12894 21564 12900 21576
rect 12952 21564 12958 21616
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 8772 21508 9873 21536
rect 8665 21499 8723 21505
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 8128 21468 8156 21499
rect 5644 21440 8156 21468
rect 8202 21428 8208 21480
rect 8260 21428 8266 21480
rect 8680 21468 8708 21499
rect 10410 21496 10416 21548
rect 10468 21536 10474 21548
rect 10505 21539 10563 21545
rect 10505 21536 10517 21539
rect 10468 21508 10517 21536
rect 10468 21496 10474 21508
rect 10505 21505 10517 21508
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 11609 21539 11667 21545
rect 11609 21505 11621 21539
rect 11655 21536 11667 21539
rect 12986 21536 12992 21548
rect 11655 21508 12992 21536
rect 11655 21505 11667 21508
rect 11609 21499 11667 21505
rect 8938 21468 8944 21480
rect 8680 21440 8944 21468
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9030 21428 9036 21480
rect 9088 21428 9094 21480
rect 10686 21468 10692 21480
rect 9692 21440 10692 21468
rect 6454 21400 6460 21412
rect 4908 21372 6460 21400
rect 2455 21369 2467 21372
rect 2409 21363 2467 21369
rect 6454 21360 6460 21372
rect 6512 21360 6518 21412
rect 7653 21403 7711 21409
rect 7653 21369 7665 21403
rect 7699 21400 7711 21403
rect 7699 21372 8064 21400
rect 7699 21369 7711 21372
rect 7653 21363 7711 21369
rect 3237 21335 3295 21341
rect 3237 21301 3249 21335
rect 3283 21332 3295 21335
rect 3694 21332 3700 21344
rect 3283 21304 3700 21332
rect 3283 21301 3295 21304
rect 3237 21295 3295 21301
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 7558 21292 7564 21344
rect 7616 21332 7622 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7616 21304 7941 21332
rect 7616 21292 7622 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 8036 21332 8064 21372
rect 8110 21360 8116 21412
rect 8168 21400 8174 21412
rect 9585 21403 9643 21409
rect 9585 21400 9597 21403
rect 8168 21372 9597 21400
rect 8168 21360 8174 21372
rect 9585 21369 9597 21372
rect 9631 21369 9643 21403
rect 9585 21363 9643 21369
rect 8386 21332 8392 21344
rect 8036 21304 8392 21332
rect 7929 21295 7987 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 8481 21335 8539 21341
rect 8481 21301 8493 21335
rect 8527 21332 8539 21335
rect 8846 21332 8852 21344
rect 8527 21304 8852 21332
rect 8527 21301 8539 21304
rect 8481 21295 8539 21301
rect 8846 21292 8852 21304
rect 8904 21292 8910 21344
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 9692 21332 9720 21440
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 11624 21468 11652 21499
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 13722 21496 13728 21548
rect 13780 21496 13786 21548
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15010 21536 15016 21548
rect 14875 21508 15016 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 10796 21440 11652 21468
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 10796 21400 10824 21440
rect 12250 21428 12256 21480
rect 12308 21428 12314 21480
rect 15120 21468 15148 21499
rect 15194 21496 15200 21548
rect 15252 21496 15258 21548
rect 15580 21545 15608 21644
rect 17313 21641 17325 21675
rect 17359 21672 17371 21675
rect 18230 21672 18236 21684
rect 17359 21644 18236 21672
rect 17359 21641 17371 21644
rect 17313 21635 17371 21641
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 23293 21675 23351 21681
rect 20272 21644 22094 21672
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 19794 21604 19800 21616
rect 16632 21576 19800 21604
rect 16632 21564 16638 21576
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21536 15623 21539
rect 15930 21536 15936 21548
rect 15611 21508 15936 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 15930 21496 15936 21508
rect 15988 21536 15994 21548
rect 15988 21508 16528 21536
rect 15988 21496 15994 21508
rect 16500 21480 16528 21508
rect 17494 21496 17500 21548
rect 17552 21496 17558 21548
rect 17880 21545 17908 21576
rect 19794 21564 19800 21576
rect 19852 21564 19858 21616
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 18132 21539 18190 21545
rect 18132 21505 18144 21539
rect 18178 21536 18190 21539
rect 18690 21536 18696 21548
rect 18178 21508 18696 21536
rect 18178 21505 18190 21508
rect 18132 21499 18190 21505
rect 18690 21496 18696 21508
rect 18748 21496 18754 21548
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 19996 21536 20024 21632
rect 20272 21545 20300 21644
rect 22066 21604 22094 21644
rect 23293 21641 23305 21675
rect 23339 21672 23351 21675
rect 23750 21672 23756 21684
rect 23339 21644 23756 21672
rect 23339 21641 23351 21644
rect 23293 21635 23351 21641
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 24121 21675 24179 21681
rect 24121 21641 24133 21675
rect 24167 21672 24179 21675
rect 24946 21672 24952 21684
rect 24167 21644 24952 21672
rect 24167 21641 24179 21644
rect 24121 21635 24179 21641
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 25314 21632 25320 21684
rect 25372 21632 25378 21684
rect 26234 21632 26240 21684
rect 26292 21632 26298 21684
rect 26697 21675 26755 21681
rect 26697 21641 26709 21675
rect 26743 21672 26755 21675
rect 26786 21672 26792 21684
rect 26743 21644 26792 21672
rect 26743 21641 26755 21644
rect 26697 21635 26755 21641
rect 26786 21632 26792 21644
rect 26844 21632 26850 21684
rect 26970 21632 26976 21684
rect 27028 21672 27034 21684
rect 27028 21644 27292 21672
rect 27028 21632 27034 21644
rect 22066 21576 23796 21604
rect 19567 21508 20024 21536
rect 20257 21539 20315 21545
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 20257 21505 20269 21539
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 20441 21539 20499 21545
rect 20441 21505 20453 21539
rect 20487 21536 20499 21539
rect 20622 21536 20628 21548
rect 20487 21508 20628 21536
rect 20487 21505 20499 21508
rect 20441 21499 20499 21505
rect 14660 21440 15148 21468
rect 10652 21372 10824 21400
rect 10652 21360 10658 21372
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 14660 21409 14688 21440
rect 15746 21428 15752 21480
rect 15804 21428 15810 21480
rect 16482 21428 16488 21480
rect 16540 21428 16546 21480
rect 11241 21403 11299 21409
rect 11241 21400 11253 21403
rect 11112 21372 11253 21400
rect 11112 21360 11118 21372
rect 11241 21369 11253 21372
rect 11287 21369 11299 21403
rect 11241 21363 11299 21369
rect 14645 21403 14703 21409
rect 14645 21369 14657 21403
rect 14691 21369 14703 21403
rect 14645 21363 14703 21369
rect 19245 21403 19303 21409
rect 19245 21369 19257 21403
rect 19291 21400 19303 21403
rect 19536 21400 19564 21499
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20956 21508 21189 21536
rect 20956 21496 20962 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21634 21496 21640 21548
rect 21692 21536 21698 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21692 21508 22017 21536
rect 21692 21496 21698 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21536 22155 21539
rect 22186 21536 22192 21548
rect 22143 21508 22192 21536
rect 22143 21505 22155 21508
rect 22097 21499 22155 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 23382 21536 23388 21548
rect 22879 21508 23388 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 23768 21480 23796 21576
rect 24670 21564 24676 21616
rect 24728 21604 24734 21616
rect 27264 21604 27292 21644
rect 27402 21607 27460 21613
rect 27402 21604 27414 21607
rect 24728 21576 27200 21604
rect 27264 21576 27414 21604
rect 24728 21564 24734 21576
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25225 21539 25283 21545
rect 25225 21536 25237 21539
rect 24912 21508 25237 21536
rect 24912 21496 24918 21508
rect 25225 21505 25237 21508
rect 25271 21505 25283 21539
rect 25225 21499 25283 21505
rect 25501 21539 25559 21545
rect 25501 21505 25513 21539
rect 25547 21505 25559 21539
rect 25501 21499 25559 21505
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20588 21440 21005 21468
rect 20588 21428 20594 21440
rect 20993 21437 21005 21440
rect 21039 21468 21051 21471
rect 21039 21440 22094 21468
rect 21039 21437 21051 21440
rect 20993 21431 21051 21437
rect 19291 21372 19564 21400
rect 19291 21369 19303 21372
rect 19245 21363 19303 21369
rect 21082 21360 21088 21412
rect 21140 21400 21146 21412
rect 21821 21403 21879 21409
rect 21821 21400 21833 21403
rect 21140 21372 21833 21400
rect 21140 21360 21146 21372
rect 21821 21369 21833 21372
rect 21867 21369 21879 21403
rect 22066 21400 22094 21440
rect 22370 21428 22376 21480
rect 22428 21428 22434 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 22922 21468 22928 21480
rect 22704 21440 22928 21468
rect 22704 21428 22710 21440
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 23477 21471 23535 21477
rect 23477 21468 23489 21471
rect 23256 21440 23489 21468
rect 23256 21428 23262 21440
rect 23477 21437 23489 21440
rect 23523 21437 23535 21471
rect 23477 21431 23535 21437
rect 23658 21428 23664 21480
rect 23716 21428 23722 21480
rect 23750 21428 23756 21480
rect 23808 21468 23814 21480
rect 24305 21471 24363 21477
rect 24305 21468 24317 21471
rect 23808 21440 24317 21468
rect 23808 21428 23814 21440
rect 24305 21437 24317 21440
rect 24351 21437 24363 21471
rect 24305 21431 24363 21437
rect 24486 21428 24492 21480
rect 24544 21428 24550 21480
rect 25516 21468 25544 21499
rect 26326 21496 26332 21548
rect 26384 21536 26390 21548
rect 26513 21539 26571 21545
rect 26513 21536 26525 21539
rect 26384 21508 26525 21536
rect 26384 21496 26390 21508
rect 26513 21505 26525 21508
rect 26559 21505 26571 21539
rect 26513 21499 26571 21505
rect 26602 21496 26608 21548
rect 26660 21496 26666 21548
rect 27172 21545 27200 21576
rect 27402 21573 27414 21576
rect 27448 21573 27460 21607
rect 27402 21567 27460 21573
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 25056 21440 25544 21468
rect 25593 21471 25651 21477
rect 23216 21400 23244 21428
rect 25056 21409 25084 21440
rect 25593 21437 25605 21471
rect 25639 21437 25651 21471
rect 25593 21431 25651 21437
rect 25777 21471 25835 21477
rect 25777 21437 25789 21471
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 22066 21372 23244 21400
rect 25041 21403 25099 21409
rect 21821 21363 21879 21369
rect 25041 21369 25053 21403
rect 25087 21369 25099 21403
rect 25041 21363 25099 21369
rect 9180 21304 9720 21332
rect 9180 21292 9186 21304
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 9916 21304 12173 21332
rect 9916 21292 9922 21304
rect 12161 21301 12173 21304
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 13630 21292 13636 21344
rect 13688 21292 13694 21344
rect 14918 21292 14924 21344
rect 14976 21292 14982 21344
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20901 21335 20959 21341
rect 20901 21301 20913 21335
rect 20947 21332 20959 21335
rect 21358 21332 21364 21344
rect 20947 21304 21364 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 21450 21292 21456 21344
rect 21508 21332 21514 21344
rect 22281 21335 22339 21341
rect 22281 21332 22293 21335
rect 21508 21304 22293 21332
rect 21508 21292 21514 21304
rect 22281 21301 22293 21304
rect 22327 21301 22339 21335
rect 22281 21295 22339 21301
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 25608 21332 25636 21431
rect 25792 21400 25820 21431
rect 26329 21403 26387 21409
rect 26329 21400 26341 21403
rect 25792 21372 26341 21400
rect 26329 21369 26341 21372
rect 26375 21369 26387 21403
rect 26329 21363 26387 21369
rect 23992 21304 25636 21332
rect 28537 21335 28595 21341
rect 23992 21292 23998 21304
rect 28537 21301 28549 21335
rect 28583 21332 28595 21335
rect 28626 21332 28632 21344
rect 28583 21304 28632 21332
rect 28583 21301 28595 21304
rect 28537 21295 28595 21301
rect 28626 21292 28632 21304
rect 28684 21292 28690 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 1670 21088 1676 21140
rect 1728 21128 1734 21140
rect 2777 21131 2835 21137
rect 2777 21128 2789 21131
rect 1728 21100 2789 21128
rect 1728 21088 1734 21100
rect 2777 21097 2789 21100
rect 2823 21097 2835 21131
rect 2777 21091 2835 21097
rect 3513 21131 3571 21137
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 3878 21128 3884 21140
rect 3559 21100 3884 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 4338 21088 4344 21140
rect 4396 21128 4402 21140
rect 4525 21131 4583 21137
rect 4525 21128 4537 21131
rect 4396 21100 4537 21128
rect 4396 21088 4402 21100
rect 4525 21097 4537 21100
rect 4571 21097 4583 21131
rect 4525 21091 4583 21097
rect 4801 21131 4859 21137
rect 4801 21097 4813 21131
rect 4847 21128 4859 21131
rect 5074 21128 5080 21140
rect 4847 21100 5080 21128
rect 4847 21097 4859 21100
rect 4801 21091 4859 21097
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 6454 21088 6460 21140
rect 6512 21088 6518 21140
rect 6822 21088 6828 21140
rect 6880 21128 6886 21140
rect 8757 21131 8815 21137
rect 8757 21128 8769 21131
rect 6880 21100 8769 21128
rect 6880 21088 6886 21100
rect 8757 21097 8769 21100
rect 8803 21097 8815 21131
rect 8757 21091 8815 21097
rect 13262 21088 13268 21140
rect 13320 21088 13326 21140
rect 13722 21088 13728 21140
rect 13780 21088 13786 21140
rect 14918 21088 14924 21140
rect 14976 21088 14982 21140
rect 15289 21131 15347 21137
rect 15289 21097 15301 21131
rect 15335 21128 15347 21131
rect 15746 21128 15752 21140
rect 15335 21100 15752 21128
rect 15335 21097 15347 21100
rect 15289 21091 15347 21097
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16114 21088 16120 21140
rect 16172 21088 16178 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 20898 21128 20904 21140
rect 16356 21100 20904 21128
rect 16356 21088 16362 21100
rect 20898 21088 20904 21100
rect 20956 21088 20962 21140
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 22278 21128 22284 21140
rect 21775 21100 22284 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 22278 21088 22284 21100
rect 22336 21088 22342 21140
rect 23474 21128 23480 21140
rect 22664 21100 23480 21128
rect 1394 20952 1400 21004
rect 1452 20952 1458 21004
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20992 3295 20995
rect 3973 20995 4031 21001
rect 3973 20992 3985 20995
rect 3283 20964 3985 20992
rect 3283 20961 3295 20964
rect 3237 20955 3295 20961
rect 3973 20961 3985 20964
rect 4019 20961 4031 20995
rect 6472 20992 6500 21088
rect 6641 20995 6699 21001
rect 6641 20992 6653 20995
rect 6472 20964 6653 20992
rect 3973 20955 4031 20961
rect 6641 20961 6653 20964
rect 6687 20961 6699 20995
rect 6641 20955 6699 20961
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20893 3111 20927
rect 3053 20887 3111 20893
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20924 3203 20927
rect 3418 20924 3424 20936
rect 3191 20896 3424 20924
rect 3191 20893 3203 20896
rect 3145 20887 3203 20893
rect 1664 20859 1722 20865
rect 1664 20825 1676 20859
rect 1710 20856 1722 20859
rect 2590 20856 2596 20868
rect 1710 20828 2596 20856
rect 1710 20825 1722 20828
rect 1664 20819 1722 20825
rect 2590 20816 2596 20828
rect 2648 20816 2654 20868
rect 3068 20856 3096 20887
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 3694 20884 3700 20936
rect 3752 20924 3758 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3752 20896 3801 20924
rect 3752 20884 3758 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4062 20884 4068 20936
rect 4120 20924 4126 20936
rect 4709 20927 4767 20933
rect 4709 20924 4721 20927
rect 4120 20896 4721 20924
rect 4120 20884 4126 20896
rect 4709 20893 4721 20896
rect 4755 20893 4767 20927
rect 4709 20887 4767 20893
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 3326 20856 3332 20868
rect 3068 20828 3332 20856
rect 3326 20816 3332 20828
rect 3384 20816 3390 20868
rect 3436 20856 3464 20884
rect 5000 20856 5028 20887
rect 5074 20884 5080 20936
rect 5132 20884 5138 20936
rect 5344 20927 5402 20933
rect 5344 20893 5356 20927
rect 5390 20924 5402 20927
rect 5902 20924 5908 20936
rect 5390 20896 5908 20924
rect 5390 20893 5402 20896
rect 5344 20887 5402 20893
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 6840 20856 6868 21088
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 10318 21060 10324 21072
rect 9732 21032 10324 21060
rect 9732 21020 9738 21032
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 10410 21020 10416 21072
rect 10468 21060 10474 21072
rect 12529 21063 12587 21069
rect 10468 21032 11100 21060
rect 10468 21020 10474 21032
rect 10873 20995 10931 21001
rect 10873 20992 10885 20995
rect 8864 20964 10885 20992
rect 7377 20927 7435 20933
rect 7377 20893 7389 20927
rect 7423 20924 7435 20927
rect 8864 20924 8892 20964
rect 10873 20961 10885 20964
rect 10919 20992 10931 20995
rect 10962 20992 10968 21004
rect 10919 20964 10968 20992
rect 10919 20961 10931 20964
rect 10873 20955 10931 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 7423 20896 8892 20924
rect 7423 20893 7435 20896
rect 7377 20887 7435 20893
rect 3436 20828 3924 20856
rect 5000 20828 6868 20856
rect 7644 20859 7702 20865
rect 3896 20800 3924 20828
rect 7644 20825 7656 20859
rect 7690 20856 7702 20859
rect 8110 20856 8116 20868
rect 7690 20828 8116 20856
rect 7690 20825 7702 20828
rect 7644 20819 7702 20825
rect 8110 20816 8116 20828
rect 8168 20816 8174 20868
rect 8202 20816 8208 20868
rect 8260 20856 8266 20868
rect 9033 20859 9091 20865
rect 9033 20856 9045 20859
rect 8260 20828 9045 20856
rect 8260 20816 8266 20828
rect 9033 20825 9045 20828
rect 9079 20825 9091 20859
rect 9033 20819 9091 20825
rect 9122 20816 9128 20868
rect 9180 20816 9186 20868
rect 10042 20816 10048 20868
rect 10100 20816 10106 20868
rect 10137 20859 10195 20865
rect 10137 20825 10149 20859
rect 10183 20856 10195 20859
rect 10410 20856 10416 20868
rect 10183 20828 10416 20856
rect 10183 20825 10195 20828
rect 10137 20819 10195 20825
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 10686 20816 10692 20868
rect 10744 20856 10750 20868
rect 11072 20856 11100 21032
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 12575 21032 12756 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 12728 21001 12756 21032
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 13740 20992 13768 21088
rect 12759 20964 13768 20992
rect 14936 20992 14964 21088
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 14936 20964 15669 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 16132 20992 16160 21088
rect 18322 21020 18328 21072
rect 18380 21020 18386 21072
rect 18693 21063 18751 21069
rect 18693 21029 18705 21063
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 20717 21063 20775 21069
rect 20717 21029 20729 21063
rect 20763 21060 20775 21063
rect 22664 21060 22692 21100
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 24121 21131 24179 21137
rect 24121 21128 24133 21131
rect 23716 21100 24133 21128
rect 23716 21088 23722 21100
rect 24121 21097 24133 21100
rect 24167 21097 24179 21131
rect 24121 21091 24179 21097
rect 24486 21088 24492 21140
rect 24544 21128 24550 21140
rect 24949 21131 25007 21137
rect 24949 21128 24961 21131
rect 24544 21100 24961 21128
rect 24544 21088 24550 21100
rect 24949 21097 24961 21100
rect 24995 21097 25007 21131
rect 24949 21091 25007 21097
rect 24302 21060 24308 21072
rect 20763 21032 22692 21060
rect 22756 21032 24308 21060
rect 20763 21029 20775 21032
rect 20717 21023 20775 21029
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 16132 20964 16313 20992
rect 15657 20955 15715 20961
rect 16301 20961 16313 20964
rect 16347 20961 16359 20995
rect 18708 20992 18736 21023
rect 16301 20955 16359 20961
rect 18156 20964 18736 20992
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20924 11207 20927
rect 11238 20924 11244 20936
rect 11195 20896 11244 20924
rect 11195 20893 11207 20896
rect 11149 20887 11207 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 12986 20884 12992 20936
rect 13044 20924 13050 20936
rect 13817 20927 13875 20933
rect 13817 20924 13829 20927
rect 13044 20896 13829 20924
rect 13044 20884 13050 20896
rect 13817 20893 13829 20896
rect 13863 20893 13875 20927
rect 13817 20887 13875 20893
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 15286 20884 15292 20936
rect 15344 20924 15350 20936
rect 15473 20927 15531 20933
rect 15473 20924 15485 20927
rect 15344 20896 15485 20924
rect 15344 20884 15350 20896
rect 15473 20893 15485 20896
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 16482 20884 16488 20936
rect 16540 20884 16546 20936
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20924 17003 20927
rect 17218 20924 17224 20936
rect 16991 20896 17224 20924
rect 16991 20893 17003 20896
rect 16945 20887 17003 20893
rect 17218 20884 17224 20896
rect 17276 20924 17282 20936
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 17276 20896 17325 20924
rect 17276 20884 17282 20896
rect 17313 20893 17325 20896
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 18156 20933 18184 20964
rect 20806 20952 20812 21004
rect 20864 20952 20870 21004
rect 22756 21001 22784 21032
rect 24302 21020 24308 21032
rect 24360 21020 24366 21072
rect 26970 21020 26976 21072
rect 27028 21020 27034 21072
rect 21085 20995 21143 21001
rect 21085 20961 21097 20995
rect 21131 20992 21143 20995
rect 22005 20995 22063 21001
rect 21131 20964 21956 20992
rect 21131 20961 21143 20964
rect 21085 20955 21143 20961
rect 18141 20927 18199 20933
rect 18141 20893 18153 20927
rect 18187 20893 18199 20927
rect 18141 20887 18199 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20924 18475 20927
rect 18874 20924 18880 20936
rect 18463 20896 18880 20924
rect 18463 20893 18475 20896
rect 18417 20887 18475 20893
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19794 20924 19800 20936
rect 19291 20896 19800 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20824 20924 20852 20952
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20824 20896 20913 20924
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 11394 20859 11452 20865
rect 11394 20856 11406 20859
rect 10744 20828 11008 20856
rect 11072 20828 11406 20856
rect 10744 20816 10750 20828
rect 2869 20791 2927 20797
rect 2869 20757 2881 20791
rect 2915 20788 2927 20791
rect 3050 20788 3056 20800
rect 2915 20760 3056 20788
rect 2915 20757 2927 20760
rect 2869 20751 2927 20757
rect 3050 20748 3056 20760
rect 3108 20748 3114 20800
rect 3878 20748 3884 20800
rect 3936 20748 3942 20800
rect 4246 20748 4252 20800
rect 4304 20788 4310 20800
rect 4433 20791 4491 20797
rect 4433 20788 4445 20791
rect 4304 20760 4445 20788
rect 4304 20748 4310 20760
rect 4433 20757 4445 20760
rect 4479 20757 4491 20791
rect 4433 20751 4491 20757
rect 7282 20748 7288 20800
rect 7340 20748 7346 20800
rect 9582 20748 9588 20800
rect 9640 20788 9646 20800
rect 10870 20788 10876 20800
rect 9640 20760 10876 20788
rect 9640 20748 9646 20760
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 10980 20788 11008 20828
rect 11394 20825 11406 20828
rect 11440 20825 11452 20859
rect 15654 20856 15660 20868
rect 11394 20819 11452 20825
rect 11532 20828 15660 20856
rect 11532 20788 11560 20828
rect 15654 20816 15660 20828
rect 15712 20856 15718 20868
rect 15712 20828 18092 20856
rect 15712 20816 15718 20828
rect 10980 20760 11560 20788
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 13357 20791 13415 20797
rect 13357 20788 13369 20791
rect 12952 20760 13369 20788
rect 12952 20748 12958 20760
rect 13357 20757 13369 20760
rect 13403 20757 13415 20791
rect 13357 20751 13415 20757
rect 13633 20791 13691 20797
rect 13633 20757 13645 20791
rect 13679 20788 13691 20791
rect 13814 20788 13820 20800
rect 13679 20760 13820 20788
rect 13679 20757 13691 20760
rect 13633 20751 13691 20757
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 17034 20748 17040 20800
rect 17092 20748 17098 20800
rect 17954 20748 17960 20800
rect 18012 20748 18018 20800
rect 18064 20788 18092 20828
rect 18230 20816 18236 20868
rect 18288 20856 18294 20868
rect 18509 20859 18567 20865
rect 18509 20856 18521 20859
rect 18288 20828 18521 20856
rect 18288 20816 18294 20828
rect 18509 20825 18521 20828
rect 18555 20825 18567 20859
rect 18509 20819 18567 20825
rect 19512 20859 19570 20865
rect 19512 20825 19524 20859
rect 19558 20856 19570 20859
rect 20088 20856 20116 20884
rect 21100 20856 21128 20955
rect 21269 20927 21327 20933
rect 21269 20893 21281 20927
rect 21315 20893 21327 20927
rect 21269 20887 21327 20893
rect 19558 20828 20116 20856
rect 20180 20828 21128 20856
rect 19558 20825 19570 20828
rect 19512 20819 19570 20825
rect 20180 20788 20208 20828
rect 18064 20760 20208 20788
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20788 20683 20791
rect 20990 20788 20996 20800
rect 20671 20760 20996 20788
rect 20671 20757 20683 20760
rect 20625 20751 20683 20757
rect 20990 20748 20996 20760
rect 21048 20748 21054 20800
rect 21284 20788 21312 20887
rect 21358 20884 21364 20936
rect 21416 20924 21422 20936
rect 21821 20927 21879 20933
rect 21821 20924 21833 20927
rect 21416 20896 21833 20924
rect 21416 20884 21422 20896
rect 21821 20893 21833 20896
rect 21867 20893 21879 20927
rect 21928 20924 21956 20964
rect 22005 20961 22017 20995
rect 22051 20992 22063 20995
rect 22741 20995 22799 21001
rect 22051 20964 22692 20992
rect 22051 20961 22063 20964
rect 22005 20955 22063 20961
rect 22557 20927 22615 20933
rect 22557 20924 22569 20927
rect 21928 20896 22569 20924
rect 21821 20887 21879 20893
rect 22557 20893 22569 20896
rect 22603 20893 22615 20927
rect 22664 20924 22692 20964
rect 22741 20961 22753 20995
rect 22787 20961 22799 20995
rect 22741 20955 22799 20961
rect 23014 20952 23020 21004
rect 23072 20952 23078 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 23477 20995 23535 21001
rect 23247 20964 23428 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 23032 20924 23060 20952
rect 22664 20896 23060 20924
rect 23293 20927 23351 20933
rect 22557 20887 22615 20893
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23400 20924 23428 20964
rect 23477 20961 23489 20995
rect 23523 20992 23535 20995
rect 24118 20992 24124 21004
rect 23523 20964 24124 20992
rect 23523 20961 23535 20964
rect 23477 20955 23535 20961
rect 24118 20952 24124 20964
rect 24176 20952 24182 21004
rect 25038 20992 25044 21004
rect 24596 20964 25044 20992
rect 23934 20924 23940 20936
rect 23400 20896 23940 20924
rect 23293 20887 23351 20893
rect 21836 20856 21864 20887
rect 23308 20856 23336 20887
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 24026 20884 24032 20936
rect 24084 20884 24090 20936
rect 24596 20933 24624 20964
rect 25038 20952 25044 20964
rect 25096 20952 25102 21004
rect 26789 20995 26847 21001
rect 26789 20961 26801 20995
rect 26835 20992 26847 20995
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 26835 20964 27997 20992
rect 26835 20961 26847 20964
rect 26789 20955 26847 20961
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24857 20927 24915 20933
rect 24857 20893 24869 20927
rect 24903 20893 24915 20927
rect 24857 20887 24915 20893
rect 25133 20927 25191 20933
rect 25133 20893 25145 20927
rect 25179 20924 25191 20927
rect 25774 20924 25780 20936
rect 25179 20896 25780 20924
rect 25179 20893 25191 20896
rect 25133 20887 25191 20893
rect 24872 20856 24900 20887
rect 25774 20884 25780 20896
rect 25832 20884 25838 20936
rect 26605 20927 26663 20933
rect 26605 20893 26617 20927
rect 26651 20893 26663 20927
rect 26605 20887 26663 20893
rect 21836 20828 23336 20856
rect 24412 20828 24900 20856
rect 26620 20856 26648 20887
rect 26878 20884 26884 20936
rect 26936 20924 26942 20936
rect 27341 20927 27399 20933
rect 27341 20924 27353 20927
rect 26936 20896 27353 20924
rect 26936 20884 26942 20896
rect 27341 20893 27353 20896
rect 27387 20893 27399 20927
rect 27341 20887 27399 20893
rect 27522 20884 27528 20936
rect 27580 20924 27586 20936
rect 27801 20927 27859 20933
rect 27801 20924 27813 20927
rect 27580 20896 27813 20924
rect 27580 20884 27586 20896
rect 27801 20893 27813 20896
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 28537 20927 28595 20933
rect 28537 20924 28549 20927
rect 27948 20896 28549 20924
rect 27948 20884 27954 20896
rect 28537 20893 28549 20896
rect 28583 20893 28595 20927
rect 28537 20887 28595 20893
rect 27706 20856 27712 20868
rect 26620 20828 27712 20856
rect 24026 20788 24032 20800
rect 21284 20760 24032 20788
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 24412 20797 24440 20828
rect 27706 20816 27712 20828
rect 27764 20816 27770 20868
rect 24397 20791 24455 20797
rect 24397 20757 24409 20791
rect 24443 20757 24455 20791
rect 24397 20751 24455 20757
rect 24673 20791 24731 20797
rect 24673 20757 24685 20791
rect 24719 20788 24731 20791
rect 24854 20788 24860 20800
rect 24719 20760 24860 20788
rect 24719 20757 24731 20760
rect 24673 20751 24731 20757
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 27430 20748 27436 20800
rect 27488 20748 27494 20800
rect 27614 20748 27620 20800
rect 27672 20748 27678 20800
rect 28353 20791 28411 20797
rect 28353 20757 28365 20791
rect 28399 20788 28411 20791
rect 28442 20788 28448 20800
rect 28399 20760 28448 20788
rect 28399 20757 28411 20760
rect 28353 20751 28411 20757
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 2590 20544 2596 20596
rect 2648 20544 2654 20596
rect 3326 20544 3332 20596
rect 3384 20584 3390 20596
rect 3513 20587 3571 20593
rect 3513 20584 3525 20587
rect 3384 20556 3525 20584
rect 3384 20544 3390 20556
rect 3513 20553 3525 20556
rect 3559 20553 3571 20587
rect 3513 20547 3571 20553
rect 6914 20544 6920 20596
rect 6972 20544 6978 20596
rect 7650 20544 7656 20596
rect 7708 20584 7714 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7708 20556 8217 20584
rect 7708 20544 7714 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8205 20547 8263 20553
rect 8386 20544 8392 20596
rect 8444 20544 8450 20596
rect 8757 20587 8815 20593
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 13173 20587 13231 20593
rect 8803 20556 13124 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 3602 20476 3608 20528
rect 3660 20516 3666 20528
rect 3660 20488 4108 20516
rect 3660 20476 3666 20488
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 1719 20420 2774 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 1412 20380 1440 20411
rect 2746 20392 2774 20420
rect 3234 20408 3240 20460
rect 3292 20448 3298 20460
rect 3694 20448 3700 20460
rect 3292 20420 3700 20448
rect 3292 20408 3298 20420
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 4080 20457 4108 20488
rect 5074 20476 5080 20528
rect 5132 20516 5138 20528
rect 5132 20488 6868 20516
rect 5132 20476 5138 20488
rect 3973 20451 4031 20457
rect 3973 20448 3985 20451
rect 3936 20420 3985 20448
rect 3936 20408 3942 20420
rect 3973 20417 3985 20420
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 4065 20451 4123 20457
rect 4065 20417 4077 20451
rect 4111 20417 4123 20451
rect 4065 20411 4123 20417
rect 4338 20408 4344 20460
rect 4396 20448 4402 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4396 20420 4537 20448
rect 4396 20408 4402 20420
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 4617 20451 4675 20457
rect 4617 20417 4629 20451
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 2038 20380 2044 20392
rect 1412 20352 2044 20380
rect 2038 20340 2044 20352
rect 2096 20340 2102 20392
rect 2746 20352 2780 20392
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 4632 20380 4660 20411
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4856 20420 4905 20448
rect 4856 20408 4862 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 5997 20451 6055 20457
rect 5997 20448 6009 20451
rect 5859 20420 6009 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 5997 20417 6009 20420
rect 6043 20417 6055 20451
rect 5997 20411 6055 20417
rect 4982 20380 4988 20392
rect 4632 20352 4988 20380
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20349 5135 20383
rect 6012 20380 6040 20411
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 6840 20457 6868 20488
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6512 20420 6561 20448
rect 6512 20408 6518 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 6932 20380 6960 20544
rect 7092 20519 7150 20525
rect 7092 20485 7104 20519
rect 7138 20516 7150 20519
rect 7282 20516 7288 20528
rect 7138 20488 7288 20516
rect 7138 20485 7150 20488
rect 7092 20479 7150 20485
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 8404 20516 8432 20544
rect 11238 20516 11244 20528
rect 8404 20488 9076 20516
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 8754 20448 8760 20460
rect 8711 20420 8760 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 8938 20408 8944 20460
rect 8996 20408 9002 20460
rect 9048 20457 9076 20488
rect 9232 20488 11244 20516
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 6012 20352 6960 20380
rect 9232 20380 9260 20488
rect 11238 20476 11244 20488
rect 11296 20516 11302 20528
rect 11296 20488 11560 20516
rect 11296 20476 11302 20488
rect 9582 20457 9588 20460
rect 9576 20448 9588 20457
rect 9543 20420 9588 20448
rect 9576 20411 9588 20420
rect 9582 20408 9588 20411
rect 9640 20408 9646 20460
rect 10778 20408 10784 20460
rect 10836 20408 10842 20460
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 11532 20457 11560 20488
rect 11790 20457 11796 20460
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 10928 20420 11161 20448
rect 10928 20408 10934 20420
rect 11149 20417 11161 20420
rect 11195 20417 11207 20451
rect 11149 20411 11207 20417
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11784 20411 11796 20457
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 9232 20352 9321 20380
rect 5077 20343 5135 20349
rect 9309 20349 9321 20352
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 1765 20315 1823 20321
rect 1765 20281 1777 20315
rect 1811 20312 1823 20315
rect 4709 20315 4767 20321
rect 1811 20284 2774 20312
rect 1811 20281 1823 20284
rect 1765 20275 1823 20281
rect 1486 20204 1492 20256
rect 1544 20204 1550 20256
rect 2746 20244 2774 20284
rect 4709 20281 4721 20315
rect 4755 20312 4767 20315
rect 5092 20312 5120 20343
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 11241 20383 11299 20389
rect 11241 20380 11253 20383
rect 10376 20352 11253 20380
rect 10376 20340 10382 20352
rect 11241 20349 11253 20352
rect 11287 20349 11299 20383
rect 11241 20343 11299 20349
rect 4755 20284 5120 20312
rect 8481 20315 8539 20321
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 8481 20281 8493 20315
rect 8527 20312 8539 20315
rect 8527 20284 9352 20312
rect 8527 20281 8539 20284
rect 8481 20275 8539 20281
rect 2958 20244 2964 20256
rect 2746 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 3326 20204 3332 20256
rect 3384 20204 3390 20256
rect 3786 20204 3792 20256
rect 3844 20204 3850 20256
rect 4154 20204 4160 20256
rect 4212 20204 4218 20256
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 4798 20244 4804 20256
rect 4387 20216 4804 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 4890 20204 4896 20256
rect 4948 20244 4954 20256
rect 5261 20247 5319 20253
rect 5261 20244 5273 20247
rect 4948 20216 5273 20244
rect 4948 20204 4954 20216
rect 5261 20213 5273 20216
rect 5307 20213 5319 20247
rect 5261 20207 5319 20213
rect 5626 20204 5632 20256
rect 5684 20204 5690 20256
rect 6086 20204 6092 20256
rect 6144 20204 6150 20256
rect 6546 20204 6552 20256
rect 6604 20244 6610 20256
rect 6641 20247 6699 20253
rect 6641 20244 6653 20247
rect 6604 20216 6653 20244
rect 6604 20204 6610 20216
rect 6641 20213 6653 20216
rect 6687 20213 6699 20247
rect 6641 20207 6699 20213
rect 9122 20204 9128 20256
rect 9180 20244 9186 20256
rect 9217 20247 9275 20253
rect 9217 20244 9229 20247
rect 9180 20216 9229 20244
rect 9180 20204 9186 20216
rect 9217 20213 9229 20216
rect 9263 20213 9275 20247
rect 9324 20244 9352 20284
rect 10042 20244 10048 20256
rect 9324 20216 10048 20244
rect 9217 20207 9275 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 10686 20204 10692 20256
rect 10744 20204 10750 20256
rect 10962 20204 10968 20256
rect 11020 20204 11026 20256
rect 11532 20244 11560 20411
rect 11790 20408 11796 20411
rect 11848 20408 11854 20460
rect 13096 20380 13124 20556
rect 13173 20553 13185 20587
rect 13219 20553 13231 20587
rect 13173 20547 13231 20553
rect 13188 20516 13216 20547
rect 13538 20544 13544 20596
rect 13596 20584 13602 20596
rect 15194 20584 15200 20596
rect 13596 20556 15200 20584
rect 13596 20544 13602 20556
rect 13188 20488 13676 20516
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 13538 20448 13544 20460
rect 13403 20420 13544 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13648 20457 13676 20488
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 13924 20380 13952 20411
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 14056 20420 14197 20448
rect 14056 20408 14062 20420
rect 14185 20417 14197 20420
rect 14231 20448 14243 20451
rect 14642 20448 14648 20460
rect 14231 20420 14648 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 14936 20457 14964 20556
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 16025 20587 16083 20593
rect 16025 20553 16037 20587
rect 16071 20584 16083 20587
rect 16482 20584 16488 20596
rect 16071 20556 16488 20584
rect 16071 20553 16083 20556
rect 16025 20547 16083 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 17276 20556 17325 20584
rect 17276 20544 17282 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 17405 20587 17463 20593
rect 17405 20553 17417 20587
rect 17451 20584 17463 20587
rect 17494 20584 17500 20596
rect 17451 20556 17500 20584
rect 17451 20553 17463 20556
rect 17405 20547 17463 20553
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 18322 20584 18328 20596
rect 18248 20556 18328 20584
rect 18248 20525 18276 20556
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 20312 20556 21128 20584
rect 20312 20544 20318 20556
rect 18233 20519 18291 20525
rect 18233 20485 18245 20519
rect 18279 20485 18291 20519
rect 18233 20479 18291 20485
rect 19794 20476 19800 20528
rect 19852 20516 19858 20528
rect 20717 20519 20775 20525
rect 20717 20516 20729 20519
rect 19852 20488 20729 20516
rect 19852 20476 19858 20488
rect 20717 20485 20729 20488
rect 20763 20485 20775 20519
rect 21100 20516 21128 20556
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21542 20584 21548 20596
rect 21232 20556 21548 20584
rect 21232 20544 21238 20556
rect 21542 20544 21548 20556
rect 21600 20584 21606 20596
rect 22278 20584 22284 20596
rect 21600 20556 22284 20584
rect 21600 20544 21606 20556
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 24026 20544 24032 20596
rect 24084 20544 24090 20596
rect 24302 20544 24308 20596
rect 24360 20544 24366 20596
rect 24854 20544 24860 20596
rect 24912 20544 24918 20596
rect 25038 20544 25044 20596
rect 25096 20544 25102 20596
rect 26605 20587 26663 20593
rect 26605 20553 26617 20587
rect 26651 20584 26663 20587
rect 27522 20584 27528 20596
rect 26651 20556 27528 20584
rect 26651 20553 26663 20556
rect 26605 20547 26663 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 27706 20584 27712 20596
rect 27663 20556 27712 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 27706 20544 27712 20556
rect 27764 20584 27770 20596
rect 28353 20587 28411 20593
rect 28353 20584 28365 20587
rect 27764 20556 28365 20584
rect 27764 20544 27770 20556
rect 28353 20553 28365 20556
rect 28399 20553 28411 20587
rect 28353 20547 28411 20553
rect 21266 20516 21272 20528
rect 21100 20488 21272 20516
rect 20717 20479 20775 20485
rect 21266 20476 21272 20488
rect 21324 20516 21330 20528
rect 21913 20519 21971 20525
rect 21913 20516 21925 20519
rect 21324 20488 21925 20516
rect 21324 20476 21330 20488
rect 21913 20485 21925 20488
rect 21959 20485 21971 20519
rect 21913 20479 21971 20485
rect 22005 20519 22063 20525
rect 22005 20485 22017 20519
rect 22051 20516 22063 20519
rect 22830 20516 22836 20528
rect 22051 20488 22836 20516
rect 22051 20485 22063 20488
rect 22005 20479 22063 20485
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 23842 20476 23848 20528
rect 23900 20516 23906 20528
rect 24670 20516 24676 20528
rect 23900 20488 24676 20516
rect 23900 20476 23906 20488
rect 24670 20476 24676 20488
rect 24728 20476 24734 20528
rect 14921 20451 14979 20457
rect 14921 20417 14933 20451
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16298 20448 16304 20460
rect 15979 20420 16304 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16298 20408 16304 20420
rect 16356 20448 16362 20460
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 16356 20420 16405 20448
rect 16356 20408 16362 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17034 20448 17040 20460
rect 16715 20420 17040 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17586 20408 17592 20460
rect 17644 20408 17650 20460
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 18012 20420 18061 20448
rect 18012 20408 18018 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20417 20039 20451
rect 19981 20411 20039 20417
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23106 20448 23112 20460
rect 23063 20420 23112 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 13096 20352 13952 20380
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14415 20352 15025 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 15197 20383 15255 20389
rect 15197 20349 15209 20383
rect 15243 20349 15255 20383
rect 15197 20343 15255 20349
rect 12897 20315 12955 20321
rect 12897 20281 12909 20315
rect 12943 20312 12955 20315
rect 12986 20312 12992 20324
rect 12943 20284 12992 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 12986 20272 12992 20284
rect 13044 20312 13050 20324
rect 13354 20312 13360 20324
rect 13044 20284 13360 20312
rect 13044 20272 13050 20284
rect 13354 20272 13360 20284
rect 13412 20272 13418 20324
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15212 20312 15240 20343
rect 15378 20340 15384 20392
rect 15436 20340 15442 20392
rect 16850 20340 16856 20392
rect 16908 20340 16914 20392
rect 18966 20340 18972 20392
rect 19024 20340 19030 20392
rect 16574 20312 16580 20324
rect 14884 20284 15240 20312
rect 15764 20284 16580 20312
rect 14884 20272 14890 20284
rect 12250 20244 12256 20256
rect 11532 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20244 12314 20256
rect 12710 20244 12716 20256
rect 12308 20216 12716 20244
rect 12308 20204 12314 20216
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13446 20204 13452 20256
rect 13504 20204 13510 20256
rect 13722 20204 13728 20256
rect 13780 20204 13786 20256
rect 13906 20204 13912 20256
rect 13964 20244 13970 20256
rect 15764 20244 15792 20284
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 19996 20312 20024 20411
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20380 22247 20383
rect 22278 20380 22284 20392
rect 22235 20352 22284 20380
rect 22235 20349 22247 20352
rect 22189 20343 22247 20349
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 20070 20312 20076 20324
rect 19996 20284 20076 20312
rect 20070 20272 20076 20284
rect 20128 20312 20134 20324
rect 23032 20312 23060 20411
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23532 20420 24225 20448
rect 23532 20408 23538 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20448 24547 20451
rect 24535 20420 24624 20448
rect 24535 20417 24547 20420
rect 24489 20411 24547 20417
rect 24596 20321 24624 20420
rect 24762 20408 24768 20460
rect 24820 20408 24826 20460
rect 24872 20448 24900 20544
rect 25056 20516 25084 20544
rect 26878 20516 26884 20528
rect 25056 20488 26884 20516
rect 25041 20451 25099 20457
rect 25041 20448 25053 20451
rect 24872 20420 25053 20448
rect 25041 20417 25053 20420
rect 25087 20417 25099 20451
rect 25041 20411 25099 20417
rect 25148 20420 25728 20448
rect 24857 20383 24915 20389
rect 24857 20349 24869 20383
rect 24903 20380 24915 20383
rect 25148 20380 25176 20420
rect 25700 20392 25728 20420
rect 26510 20408 26516 20460
rect 26568 20408 26574 20460
rect 26804 20457 26832 20488
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 26789 20451 26847 20457
rect 26789 20417 26801 20451
rect 26835 20417 26847 20451
rect 26789 20411 26847 20417
rect 27062 20408 27068 20460
rect 27120 20408 27126 20460
rect 27157 20451 27215 20457
rect 27157 20417 27169 20451
rect 27203 20448 27215 20451
rect 27430 20448 27436 20460
rect 27203 20420 27436 20448
rect 27203 20417 27215 20420
rect 27157 20411 27215 20417
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 27614 20408 27620 20460
rect 27672 20448 27678 20460
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 27672 20420 27905 20448
rect 27672 20408 27678 20420
rect 27893 20417 27905 20420
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 24903 20352 25176 20380
rect 24903 20349 24915 20352
rect 24857 20343 24915 20349
rect 25590 20340 25596 20392
rect 25648 20340 25654 20392
rect 25682 20340 25688 20392
rect 25740 20340 25746 20392
rect 25774 20340 25780 20392
rect 25832 20340 25838 20392
rect 26602 20340 26608 20392
rect 26660 20380 26666 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26660 20352 26985 20380
rect 26660 20340 26666 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 27080 20380 27108 20408
rect 27706 20380 27712 20392
rect 27080 20352 27712 20380
rect 26973 20343 27031 20349
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 20128 20284 23060 20312
rect 24581 20315 24639 20321
rect 20128 20272 20134 20284
rect 24581 20281 24593 20315
rect 24627 20281 24639 20315
rect 24581 20275 24639 20281
rect 24780 20284 27568 20312
rect 13964 20216 15792 20244
rect 13964 20204 13970 20216
rect 15838 20204 15844 20256
rect 15896 20204 15902 20256
rect 16206 20204 16212 20256
rect 16264 20204 16270 20256
rect 20530 20204 20536 20256
rect 20588 20244 20594 20256
rect 21637 20247 21695 20253
rect 21637 20244 21649 20247
rect 20588 20216 21649 20244
rect 20588 20204 20594 20216
rect 21637 20213 21649 20216
rect 21683 20213 21695 20247
rect 21637 20207 21695 20213
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 24780 20244 24808 20284
rect 27540 20256 27568 20284
rect 21784 20216 24808 20244
rect 25501 20247 25559 20253
rect 21784 20204 21790 20216
rect 25501 20213 25513 20247
rect 25547 20244 25559 20247
rect 25958 20244 25964 20256
rect 25547 20216 25964 20244
rect 25547 20213 25559 20216
rect 25501 20207 25559 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26326 20204 26332 20256
rect 26384 20204 26390 20256
rect 27522 20204 27528 20256
rect 27580 20204 27586 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 2038 20000 2044 20052
rect 2096 20040 2102 20052
rect 2777 20043 2835 20049
rect 2777 20040 2789 20043
rect 2096 20012 2789 20040
rect 2096 20000 2102 20012
rect 2777 20009 2789 20012
rect 2823 20009 2835 20043
rect 2777 20003 2835 20009
rect 4246 20000 4252 20052
rect 4304 20000 4310 20052
rect 4338 20000 4344 20052
rect 4396 20040 4402 20052
rect 4525 20043 4583 20049
rect 4525 20040 4537 20043
rect 4396 20012 4537 20040
rect 4396 20000 4402 20012
rect 4525 20009 4537 20012
rect 4571 20009 4583 20043
rect 4525 20003 4583 20009
rect 7837 20043 7895 20049
rect 7837 20009 7849 20043
rect 7883 20040 7895 20043
rect 10778 20040 10784 20052
rect 7883 20012 10784 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 13504 20012 14412 20040
rect 13504 20000 13510 20012
rect 4706 19932 4712 19984
rect 4764 19972 4770 19984
rect 4982 19972 4988 19984
rect 4764 19944 4988 19972
rect 4764 19932 4770 19944
rect 4982 19932 4988 19944
rect 5040 19972 5046 19984
rect 5442 19972 5448 19984
rect 5040 19944 5448 19972
rect 5040 19932 5046 19944
rect 5442 19932 5448 19944
rect 5500 19972 5506 19984
rect 8386 19972 8392 19984
rect 5500 19944 8392 19972
rect 5500 19932 5506 19944
rect 8386 19932 8392 19944
rect 8444 19932 8450 19984
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 9582 19972 9588 19984
rect 8812 19944 9588 19972
rect 8812 19932 8818 19944
rect 9582 19932 9588 19944
rect 9640 19932 9646 19984
rect 9769 19975 9827 19981
rect 9769 19941 9781 19975
rect 9815 19972 9827 19975
rect 9950 19972 9956 19984
rect 9815 19944 9956 19972
rect 9815 19941 9827 19944
rect 9769 19935 9827 19941
rect 9950 19932 9956 19944
rect 10008 19972 10014 19984
rect 10229 19975 10287 19981
rect 10229 19972 10241 19975
rect 10008 19944 10241 19972
rect 10008 19932 10014 19944
rect 10229 19941 10241 19944
rect 10275 19941 10287 19975
rect 10229 19935 10287 19941
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19941 13783 19975
rect 13725 19935 13783 19941
rect 5074 19904 5080 19916
rect 2746 19876 5080 19904
rect 1394 19796 1400 19848
rect 1452 19836 1458 19848
rect 2746 19836 2774 19876
rect 5074 19864 5080 19876
rect 5132 19904 5138 19916
rect 6365 19907 6423 19913
rect 6365 19904 6377 19907
rect 5132 19876 6377 19904
rect 5132 19864 5138 19876
rect 6365 19873 6377 19876
rect 6411 19873 6423 19907
rect 6365 19867 6423 19873
rect 6730 19864 6736 19916
rect 6788 19904 6794 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 6788 19876 7389 19904
rect 6788 19864 6794 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 8036 19876 9076 19904
rect 1452 19808 2774 19836
rect 1452 19796 1458 19808
rect 2958 19796 2964 19848
rect 3016 19796 3022 19848
rect 3050 19796 3056 19848
rect 3108 19836 3114 19848
rect 3145 19839 3203 19845
rect 3145 19836 3157 19839
rect 3108 19808 3157 19836
rect 3108 19796 3114 19808
rect 3145 19805 3157 19808
rect 3191 19805 3203 19839
rect 3145 19799 3203 19805
rect 3326 19796 3332 19848
rect 3384 19796 3390 19848
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3620 19808 3801 19836
rect 1664 19771 1722 19777
rect 1664 19737 1676 19771
rect 1710 19768 1722 19771
rect 3344 19768 3372 19796
rect 1710 19740 3372 19768
rect 1710 19737 1722 19740
rect 1664 19731 1722 19737
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 3620 19709 3648 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4706 19796 4712 19848
rect 4764 19796 4770 19848
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19836 5687 19839
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 5675 19808 6653 19836
rect 5675 19805 5687 19808
rect 5629 19799 5687 19805
rect 6641 19805 6653 19808
rect 6687 19836 6699 19839
rect 7282 19836 7288 19848
rect 6687 19808 7288 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 8036 19845 8064 19876
rect 9048 19848 9076 19876
rect 10410 19864 10416 19916
rect 10468 19904 10474 19916
rect 10468 19876 12020 19904
rect 10468 19864 10474 19876
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19836 8171 19839
rect 8202 19836 8208 19848
rect 8159 19808 8208 19836
rect 8159 19805 8171 19808
rect 8113 19799 8171 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 4890 19728 4896 19780
rect 4948 19728 4954 19780
rect 4985 19771 5043 19777
rect 4985 19737 4997 19771
rect 5031 19737 5043 19771
rect 4985 19731 5043 19737
rect 5537 19771 5595 19777
rect 5537 19737 5549 19771
rect 5583 19768 5595 19771
rect 5994 19768 6000 19780
rect 5583 19740 6000 19768
rect 5583 19737 5595 19740
rect 5537 19731 5595 19737
rect 3605 19703 3663 19709
rect 3605 19700 3617 19703
rect 3568 19672 3617 19700
rect 3568 19660 3574 19672
rect 3605 19669 3617 19672
rect 3651 19669 3663 19703
rect 5000 19700 5028 19731
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 6086 19728 6092 19780
rect 6144 19728 6150 19780
rect 7190 19728 7196 19780
rect 7248 19768 7254 19780
rect 8312 19768 8340 19799
rect 9030 19796 9036 19848
rect 9088 19796 9094 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 10045 19839 10103 19845
rect 10045 19805 10057 19839
rect 10091 19836 10103 19839
rect 10502 19836 10508 19848
rect 10091 19808 10508 19836
rect 10091 19805 10103 19808
rect 10045 19799 10103 19805
rect 7248 19740 8340 19768
rect 7248 19728 7254 19740
rect 6104 19700 6132 19728
rect 5000 19672 6132 19700
rect 3605 19663 3663 19669
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 9876 19700 9904 19799
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 10873 19771 10931 19777
rect 10873 19737 10885 19771
rect 10919 19737 10931 19771
rect 10873 19731 10931 19737
rect 8812 19672 9904 19700
rect 10888 19700 10916 19731
rect 10962 19728 10968 19780
rect 11020 19728 11026 19780
rect 11330 19728 11336 19780
rect 11388 19768 11394 19780
rect 11992 19777 12020 19876
rect 12710 19864 12716 19916
rect 12768 19864 12774 19916
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13740 19904 13768 19935
rect 13906 19932 13912 19984
rect 13964 19932 13970 19984
rect 13219 19876 13768 19904
rect 13924 19904 13952 19932
rect 14384 19913 14412 20012
rect 14826 20000 14832 20052
rect 14884 20000 14890 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15436 20012 16037 20040
rect 15436 20000 15442 20012
rect 16025 20009 16037 20012
rect 16071 20009 16083 20043
rect 16025 20003 16083 20009
rect 16206 20000 16212 20052
rect 16264 20000 16270 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 16850 20040 16856 20052
rect 16531 20012 16856 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17586 20000 17592 20052
rect 17644 20000 17650 20052
rect 17954 20000 17960 20052
rect 18012 20000 18018 20052
rect 20625 20043 20683 20049
rect 20625 20009 20637 20043
rect 20671 20040 20683 20043
rect 20806 20040 20812 20052
rect 20671 20012 20812 20040
rect 20671 20009 20683 20012
rect 20625 20003 20683 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 21634 20000 21640 20052
rect 21692 20040 21698 20052
rect 25593 20043 25651 20049
rect 21692 20012 23980 20040
rect 21692 20000 21698 20012
rect 15838 19932 15844 19984
rect 15896 19932 15902 19984
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 13924 19876 14197 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 14369 19907 14427 19913
rect 14369 19873 14381 19907
rect 14415 19873 14427 19907
rect 16224 19904 16252 20000
rect 17604 19972 17632 20000
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 17604 19944 18797 19972
rect 18785 19941 18797 19944
rect 18831 19941 18843 19975
rect 18785 19935 18843 19941
rect 20898 19932 20904 19984
rect 20956 19972 20962 19984
rect 21726 19972 21732 19984
rect 20956 19944 21732 19972
rect 20956 19932 20962 19944
rect 21726 19932 21732 19944
rect 21784 19932 21790 19984
rect 17129 19907 17187 19913
rect 16224 19876 16712 19904
rect 14369 19867 14427 19873
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13872 19808 13921 19836
rect 13872 19796 13878 19808
rect 13909 19805 13921 19808
rect 13955 19805 13967 19839
rect 13909 19799 13967 19805
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15378 19796 15384 19848
rect 15436 19796 15442 19848
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19836 15991 19839
rect 16206 19836 16212 19848
rect 15979 19808 16212 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16684 19845 16712 19876
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 17175 19876 17509 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 22370 19904 22376 19916
rect 20855 19876 22376 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 23842 19864 23848 19916
rect 23900 19864 23906 19916
rect 23952 19904 23980 20012
rect 25593 20009 25605 20043
rect 25639 20040 25651 20043
rect 25774 20040 25780 20052
rect 25639 20012 25780 20040
rect 25639 20009 25651 20012
rect 25593 20003 25651 20009
rect 25774 20000 25780 20012
rect 25832 20000 25838 20052
rect 25958 20000 25964 20052
rect 26016 20000 26022 20052
rect 26326 20000 26332 20052
rect 26384 20000 26390 20052
rect 26510 20000 26516 20052
rect 26568 20040 26574 20052
rect 26697 20043 26755 20049
rect 26697 20040 26709 20043
rect 26568 20012 26709 20040
rect 26568 20000 26574 20012
rect 26697 20009 26709 20012
rect 26743 20009 26755 20043
rect 26697 20003 26755 20009
rect 26970 20000 26976 20052
rect 27028 20000 27034 20052
rect 27249 20043 27307 20049
rect 27249 20009 27261 20043
rect 27295 20040 27307 20043
rect 27338 20040 27344 20052
rect 27295 20012 27344 20040
rect 27295 20009 27307 20012
rect 27249 20003 27307 20009
rect 27338 20000 27344 20012
rect 27396 20000 27402 20052
rect 24121 19975 24179 19981
rect 24121 19941 24133 19975
rect 24167 19972 24179 19975
rect 24167 19944 24900 19972
rect 24167 19941 24179 19944
rect 24121 19935 24179 19941
rect 23952 19876 24716 19904
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 11388 19740 11897 19768
rect 11388 19728 11394 19740
rect 11885 19737 11897 19740
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 11977 19771 12035 19777
rect 11977 19737 11989 19771
rect 12023 19768 12035 19771
rect 16298 19768 16304 19780
rect 12023 19740 16304 19768
rect 12023 19737 12035 19740
rect 11977 19731 12035 19737
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 17052 19768 17080 19799
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 17313 19839 17371 19845
rect 17313 19836 17325 19839
rect 17276 19808 17325 19836
rect 17276 19796 17282 19808
rect 17313 19805 17325 19808
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 18046 19796 18052 19848
rect 18104 19836 18110 19848
rect 18141 19839 18199 19845
rect 18141 19836 18153 19839
rect 18104 19808 18153 19836
rect 18104 19796 18110 19808
rect 18141 19805 18153 19808
rect 18187 19836 18199 19839
rect 18969 19839 19027 19845
rect 18969 19836 18981 19839
rect 18187 19808 18981 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 18969 19805 18981 19808
rect 19015 19805 19027 19839
rect 18969 19799 19027 19805
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 18064 19768 18092 19796
rect 17052 19740 18092 19768
rect 13078 19700 13084 19712
rect 10888 19672 13084 19700
rect 8812 19660 8818 19672
rect 13078 19660 13084 19672
rect 13136 19700 13142 19712
rect 13633 19703 13691 19709
rect 13633 19700 13645 19703
rect 13136 19672 13645 19700
rect 13136 19660 13142 19672
rect 13633 19669 13645 19672
rect 13679 19669 13691 19703
rect 13633 19663 13691 19669
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 17218 19700 17224 19712
rect 15896 19672 17224 19700
rect 15896 19660 15902 19672
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 19260 19700 19288 19799
rect 21726 19796 21732 19848
rect 21784 19796 21790 19848
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19836 22063 19839
rect 22741 19839 22799 19845
rect 22051 19808 22692 19836
rect 22051 19805 22063 19808
rect 22005 19799 22063 19805
rect 19512 19771 19570 19777
rect 19512 19737 19524 19771
rect 19558 19768 19570 19771
rect 20901 19771 20959 19777
rect 19558 19740 20852 19768
rect 19558 19737 19570 19740
rect 19512 19731 19570 19737
rect 19610 19700 19616 19712
rect 19260 19672 19616 19700
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 20824 19700 20852 19740
rect 20901 19737 20913 19771
rect 20947 19768 20959 19771
rect 21450 19768 21456 19780
rect 20947 19740 21456 19768
rect 20947 19737 20959 19740
rect 20901 19731 20959 19737
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 21744 19768 21772 19796
rect 21821 19771 21879 19777
rect 21821 19768 21833 19771
rect 21744 19740 21833 19768
rect 21821 19737 21833 19740
rect 21867 19737 21879 19771
rect 21821 19731 21879 19737
rect 22554 19728 22560 19780
rect 22612 19728 22618 19780
rect 22664 19768 22692 19808
rect 22741 19805 22753 19839
rect 22787 19836 22799 19839
rect 23860 19836 23888 19864
rect 24688 19845 24716 19876
rect 24872 19848 24900 19944
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 25314 19904 25320 19916
rect 25096 19876 25320 19904
rect 25096 19864 25102 19876
rect 25314 19864 25320 19876
rect 25372 19904 25378 19916
rect 25976 19913 26004 20000
rect 25961 19907 26019 19913
rect 25372 19876 25544 19904
rect 25372 19864 25378 19876
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 22787 19808 23888 19836
rect 23952 19808 24593 19836
rect 22787 19805 22799 19808
rect 22741 19799 22799 19805
rect 23008 19771 23066 19777
rect 22664 19740 22784 19768
rect 22756 19712 22784 19740
rect 23008 19737 23020 19771
rect 23054 19768 23066 19771
rect 23474 19768 23480 19780
rect 23054 19740 23480 19768
rect 23054 19737 23066 19740
rect 23008 19731 23066 19737
rect 23474 19728 23480 19740
rect 23532 19728 23538 19780
rect 22462 19700 22468 19712
rect 20824 19672 22468 19700
rect 22462 19660 22468 19672
rect 22520 19660 22526 19712
rect 22738 19660 22744 19712
rect 22796 19700 22802 19712
rect 23952 19700 23980 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 24596 19768 24624 19799
rect 24854 19796 24860 19848
rect 24912 19796 24918 19848
rect 25516 19845 25544 19876
rect 25961 19873 25973 19907
rect 26007 19873 26019 19907
rect 25961 19867 26019 19873
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19904 26203 19907
rect 26344 19904 26372 20000
rect 26605 19975 26663 19981
rect 26605 19941 26617 19975
rect 26651 19972 26663 19975
rect 26988 19972 27016 20000
rect 27890 19972 27896 19984
rect 26651 19944 27016 19972
rect 27080 19944 27896 19972
rect 26651 19941 26663 19944
rect 26605 19935 26663 19941
rect 27080 19904 27108 19944
rect 27890 19932 27896 19944
rect 27948 19932 27954 19984
rect 26191 19876 26372 19904
rect 26896 19876 27108 19904
rect 26191 19873 26203 19876
rect 26145 19867 26203 19873
rect 26896 19845 26924 19876
rect 27154 19864 27160 19916
rect 27212 19904 27218 19916
rect 27212 19876 28212 19904
rect 27212 19864 27218 19876
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19805 25191 19839
rect 25133 19799 25191 19805
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 26881 19839 26939 19845
rect 25547 19808 26832 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25148 19768 25176 19799
rect 24596 19740 25176 19768
rect 25424 19768 25452 19799
rect 26418 19768 26424 19780
rect 25424 19740 26424 19768
rect 26418 19728 26424 19740
rect 26476 19728 26482 19780
rect 26804 19768 26832 19808
rect 26881 19805 26893 19839
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27019 19808 27445 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27433 19805 27445 19808
rect 27479 19805 27491 19839
rect 27433 19799 27491 19805
rect 26988 19768 27016 19799
rect 27522 19796 27528 19848
rect 27580 19796 27586 19848
rect 27890 19796 27896 19848
rect 27948 19796 27954 19848
rect 28184 19845 28212 19876
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 26804 19740 27016 19768
rect 27246 19728 27252 19780
rect 27304 19728 27310 19780
rect 27614 19728 27620 19780
rect 27672 19768 27678 19780
rect 28261 19771 28319 19777
rect 28261 19768 28273 19771
rect 27672 19740 28273 19768
rect 27672 19728 27678 19740
rect 28261 19737 28273 19740
rect 28307 19737 28319 19771
rect 28261 19731 28319 19737
rect 22796 19672 23980 19700
rect 22796 19660 22802 19672
rect 24302 19660 24308 19712
rect 24360 19700 24366 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 24360 19672 24409 19700
rect 24360 19660 24366 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 24762 19660 24768 19712
rect 24820 19660 24826 19712
rect 24946 19660 24952 19712
rect 25004 19660 25010 19712
rect 25222 19660 25228 19712
rect 25280 19660 25286 19712
rect 27062 19660 27068 19712
rect 27120 19660 27126 19712
rect 27264 19700 27292 19728
rect 27706 19700 27712 19712
rect 27264 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 27982 19660 27988 19712
rect 28040 19660 28046 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 1486 19456 1492 19508
rect 1544 19456 1550 19508
rect 2774 19456 2780 19508
rect 2832 19456 2838 19508
rect 3510 19456 3516 19508
rect 3568 19456 3574 19508
rect 3786 19456 3792 19508
rect 3844 19456 3850 19508
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 3970 19496 3976 19508
rect 3927 19468 3976 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 4948 19468 5365 19496
rect 4948 19456 4954 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5353 19459 5411 19465
rect 5442 19456 5448 19508
rect 5500 19456 5506 19508
rect 5626 19456 5632 19508
rect 5684 19456 5690 19508
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 5767 19468 6592 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 1504 19428 1532 19456
rect 3804 19428 3832 19456
rect 1504 19400 2774 19428
rect 3804 19400 4108 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 1664 19363 1722 19369
rect 1664 19329 1676 19363
rect 1710 19360 1722 19363
rect 2222 19360 2228 19372
rect 1710 19332 2228 19360
rect 1710 19329 1722 19332
rect 1664 19323 1722 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 2746 19360 2774 19400
rect 2869 19363 2927 19369
rect 2869 19360 2881 19363
rect 2746 19332 2881 19360
rect 2869 19329 2881 19332
rect 2915 19329 2927 19363
rect 2869 19323 2927 19329
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 3694 19360 3700 19372
rect 3568 19332 3700 19360
rect 3568 19320 3574 19332
rect 3694 19320 3700 19332
rect 3752 19360 3758 19372
rect 4080 19369 4108 19400
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3752 19332 3801 19360
rect 3752 19320 3758 19332
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4154 19320 4160 19372
rect 4212 19320 4218 19372
rect 4246 19320 4252 19372
rect 4304 19360 4310 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4304 19332 4721 19360
rect 4304 19320 4310 19332
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 4798 19320 4804 19372
rect 4856 19360 4862 19372
rect 4893 19363 4951 19369
rect 4893 19360 4905 19363
rect 4856 19332 4905 19360
rect 4856 19320 4862 19332
rect 4893 19329 4905 19332
rect 4939 19329 4951 19363
rect 5460 19360 5488 19456
rect 5644 19428 5672 19456
rect 6564 19437 6592 19468
rect 7742 19456 7748 19508
rect 7800 19456 7806 19508
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 10686 19496 10692 19508
rect 9088 19468 10692 19496
rect 9088 19456 9094 19468
rect 6549 19431 6607 19437
rect 5644 19400 5948 19428
rect 5920 19369 5948 19400
rect 6549 19397 6561 19431
rect 6595 19397 6607 19431
rect 7760 19428 7788 19456
rect 7837 19431 7895 19437
rect 7837 19428 7849 19431
rect 7760 19400 7849 19428
rect 6549 19391 6607 19397
rect 7837 19397 7849 19400
rect 7883 19397 7895 19431
rect 7837 19391 7895 19397
rect 8294 19388 8300 19440
rect 8352 19428 8358 19440
rect 9398 19428 9404 19440
rect 8352 19400 9404 19428
rect 8352 19388 8358 19400
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5460 19332 5641 19360
rect 4893 19323 4951 19329
rect 5629 19329 5641 19332
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 6052 19332 6316 19360
rect 6052 19320 6058 19332
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 4172 19292 4200 19320
rect 3099 19264 4200 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 6288 19224 6316 19332
rect 7282 19320 7288 19372
rect 7340 19360 7346 19372
rect 7561 19363 7619 19369
rect 7561 19360 7573 19363
rect 7340 19332 7573 19360
rect 7340 19320 7346 19332
rect 7561 19329 7573 19332
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 9600 19369 9628 19468
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 12894 19496 12900 19508
rect 11624 19468 12900 19496
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19428 9735 19431
rect 10413 19431 10471 19437
rect 10413 19428 10425 19431
rect 9723 19400 10425 19428
rect 9723 19397 9735 19400
rect 9677 19391 9735 19397
rect 10413 19397 10425 19400
rect 10459 19397 10471 19431
rect 10413 19391 10471 19397
rect 11330 19388 11336 19440
rect 11388 19388 11394 19440
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19329 9643 19363
rect 9858 19360 9864 19372
rect 9585 19323 9643 19329
rect 9692 19332 9864 19360
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 9508 19292 9536 19323
rect 9692 19292 9720 19332
rect 9858 19320 9864 19332
rect 9916 19360 9922 19372
rect 9916 19332 9996 19360
rect 9916 19320 9922 19332
rect 9508 19264 9720 19292
rect 7006 19224 7012 19236
rect 6288 19196 7012 19224
rect 7006 19184 7012 19196
rect 7064 19184 7070 19236
rect 9968 19224 9996 19332
rect 10042 19320 10048 19372
rect 10100 19320 10106 19372
rect 11624 19369 11652 19468
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 12986 19456 12992 19508
rect 13044 19456 13050 19508
rect 14921 19499 14979 19505
rect 14921 19465 14933 19499
rect 14967 19496 14979 19499
rect 15194 19496 15200 19508
rect 14967 19468 15200 19496
rect 14967 19465 14979 19468
rect 14921 19459 14979 19465
rect 15194 19456 15200 19468
rect 15252 19496 15258 19508
rect 15252 19468 15332 19496
rect 15252 19456 15258 19468
rect 12253 19431 12311 19437
rect 12253 19397 12265 19431
rect 12299 19428 12311 19431
rect 13004 19428 13032 19456
rect 12299 19400 13032 19428
rect 13357 19431 13415 19437
rect 12299 19397 12311 19400
rect 12253 19391 12311 19397
rect 13357 19397 13369 19431
rect 13403 19428 13415 19431
rect 13403 19400 14320 19428
rect 13403 19397 13415 19400
rect 13357 19391 13415 19397
rect 11609 19363 11667 19369
rect 11609 19329 11621 19363
rect 11655 19329 11667 19363
rect 11609 19323 11667 19329
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19360 12403 19363
rect 12434 19360 12440 19372
rect 12391 19332 12440 19360
rect 12391 19329 12403 19332
rect 12345 19323 12403 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 13265 19363 13323 19369
rect 13265 19329 13277 19363
rect 13311 19360 13323 19363
rect 13538 19360 13544 19372
rect 13311 19332 13544 19360
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 13538 19320 13544 19332
rect 13596 19360 13602 19372
rect 13596 19332 13860 19360
rect 13596 19320 13602 19332
rect 13832 19304 13860 19332
rect 14182 19320 14188 19372
rect 14240 19320 14246 19372
rect 14292 19360 14320 19400
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 14608 19400 15056 19428
rect 14608 19388 14614 19400
rect 14292 19332 14872 19360
rect 10318 19252 10324 19304
rect 10376 19252 10382 19304
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12529 19295 12587 19301
rect 11839 19264 12434 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 11054 19224 11060 19236
rect 9968 19196 11060 19224
rect 11054 19184 11060 19196
rect 11112 19184 11118 19236
rect 12406 19224 12434 19264
rect 12529 19261 12541 19295
rect 12575 19292 12587 19295
rect 13170 19292 13176 19304
rect 12575 19264 13176 19292
rect 12575 19261 12587 19264
rect 12529 19255 12587 19261
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 13630 19252 13636 19304
rect 13688 19252 13694 19304
rect 13814 19252 13820 19304
rect 13872 19252 13878 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 13722 19224 13728 19236
rect 12406 19196 13728 19224
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 3602 19116 3608 19168
rect 3660 19116 3666 19168
rect 5442 19116 5448 19168
rect 5500 19116 5506 19168
rect 6086 19116 6092 19168
rect 6144 19116 6150 19168
rect 7377 19159 7435 19165
rect 7377 19125 7389 19159
rect 7423 19156 7435 19159
rect 8294 19156 8300 19168
rect 7423 19128 8300 19156
rect 7423 19125 7435 19128
rect 7377 19119 7435 19125
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 9030 19156 9036 19168
rect 8628 19128 9036 19156
rect 8628 19116 8634 19128
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9858 19116 9864 19168
rect 9916 19116 9922 19168
rect 14292 19156 14320 19255
rect 14458 19252 14464 19304
rect 14516 19252 14522 19304
rect 14844 19224 14872 19332
rect 15028 19301 15056 19400
rect 15304 19360 15332 19468
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15436 19468 15761 19496
rect 15436 19456 15442 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 15749 19459 15807 19465
rect 16025 19499 16083 19505
rect 16025 19465 16037 19499
rect 16071 19465 16083 19499
rect 16025 19459 16083 19465
rect 15657 19363 15715 19369
rect 15657 19360 15669 19363
rect 15304 19332 15669 19360
rect 15657 19329 15669 19332
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 16040 19360 16068 19459
rect 18046 19456 18052 19508
rect 18104 19456 18110 19508
rect 19886 19456 19892 19508
rect 19944 19496 19950 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 19944 19468 21465 19496
rect 19944 19456 19950 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22462 19456 22468 19508
rect 22520 19456 22526 19508
rect 22557 19499 22615 19505
rect 22557 19465 22569 19499
rect 22603 19496 22615 19499
rect 22603 19468 23336 19496
rect 22603 19465 22615 19468
rect 22557 19459 22615 19465
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 16356 19400 19564 19428
rect 16356 19388 16362 19400
rect 15979 19332 16068 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 16206 19320 16212 19372
rect 16264 19320 16270 19372
rect 16936 19363 16994 19369
rect 16936 19329 16948 19363
rect 16982 19360 16994 19363
rect 17310 19360 17316 19372
rect 16982 19332 17316 19360
rect 16982 19329 16994 19332
rect 16936 19323 16994 19329
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 19536 19360 19564 19400
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 20809 19431 20867 19437
rect 20809 19428 20821 19431
rect 19668 19400 20821 19428
rect 19668 19388 19674 19400
rect 20809 19397 20821 19400
rect 20855 19397 20867 19431
rect 20809 19391 20867 19397
rect 23106 19388 23112 19440
rect 23164 19428 23170 19440
rect 23201 19431 23259 19437
rect 23201 19428 23213 19431
rect 23164 19400 23213 19428
rect 23164 19388 23170 19400
rect 23201 19397 23213 19400
rect 23247 19397 23259 19431
rect 23201 19391 23259 19397
rect 20070 19360 20076 19372
rect 19536 19332 20076 19360
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20990 19320 20996 19372
rect 21048 19360 21054 19372
rect 21353 19369 21411 19375
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 21048 19332 21097 19360
rect 21048 19320 21054 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21353 19346 21365 19369
rect 21399 19346 21411 19369
rect 21353 19329 21364 19346
rect 21085 19323 21143 19329
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19261 15255 19295
rect 15197 19255 15255 19261
rect 16669 19295 16727 19301
rect 16669 19261 16681 19295
rect 16715 19261 16727 19295
rect 16669 19255 16727 19261
rect 15212 19224 15240 19255
rect 14844 19196 15240 19224
rect 15378 19156 15384 19168
rect 14292 19128 15384 19156
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 16684 19156 16712 19255
rect 18322 19252 18328 19304
rect 18380 19252 18386 19304
rect 18966 19252 18972 19304
rect 19024 19252 19030 19304
rect 21358 19294 21364 19329
rect 21416 19294 21422 19346
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 22741 19363 22799 19369
rect 22741 19360 22753 19363
rect 21508 19332 22753 19360
rect 21508 19320 21514 19332
rect 22741 19329 22753 19332
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 23017 19363 23075 19369
rect 23017 19329 23029 19363
rect 23063 19360 23075 19363
rect 23308 19360 23336 19468
rect 25590 19388 25596 19440
rect 25648 19428 25654 19440
rect 25774 19428 25780 19440
rect 25648 19400 25780 19428
rect 25648 19388 25654 19400
rect 25774 19388 25780 19400
rect 25832 19388 25838 19440
rect 27890 19428 27896 19440
rect 26436 19400 27896 19428
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23063 19332 23336 19360
rect 23952 19332 24041 19360
rect 23063 19329 23075 19332
rect 23017 19323 23075 19329
rect 21821 19295 21879 19301
rect 21821 19261 21833 19295
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 18932 19196 21312 19224
rect 18932 19184 18938 19196
rect 17586 19156 17592 19168
rect 16684 19128 17592 19156
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21177 19159 21235 19165
rect 21177 19156 21189 19159
rect 20864 19128 21189 19156
rect 20864 19116 20870 19128
rect 21177 19125 21189 19128
rect 21223 19125 21235 19159
rect 21284 19156 21312 19196
rect 21836 19156 21864 19255
rect 22830 19184 22836 19236
rect 22888 19184 22894 19236
rect 23952 19168 23980 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19360 24271 19363
rect 25130 19360 25136 19372
rect 24259 19332 25136 19360
rect 24259 19329 24271 19332
rect 24213 19323 24271 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25222 19320 25228 19372
rect 25280 19360 25286 19372
rect 26436 19369 26464 19400
rect 27890 19388 27896 19400
rect 27948 19388 27954 19440
rect 25869 19363 25927 19369
rect 25869 19360 25881 19363
rect 25280 19332 25881 19360
rect 25280 19320 25286 19332
rect 25869 19329 25881 19332
rect 25915 19329 25927 19363
rect 26421 19363 26479 19369
rect 26421 19360 26433 19363
rect 25869 19323 25927 19329
rect 26160 19332 26433 19360
rect 24394 19252 24400 19304
rect 24452 19252 24458 19304
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 24949 19295 25007 19301
rect 24949 19292 24961 19295
rect 24912 19264 24961 19292
rect 24912 19252 24918 19264
rect 24949 19261 24961 19264
rect 24995 19261 25007 19295
rect 24949 19255 25007 19261
rect 24964 19224 24992 19255
rect 25038 19252 25044 19304
rect 25096 19292 25102 19304
rect 25685 19295 25743 19301
rect 25685 19292 25697 19295
rect 25096 19264 25697 19292
rect 25096 19252 25102 19264
rect 25685 19261 25697 19264
rect 25731 19261 25743 19295
rect 25685 19255 25743 19261
rect 26050 19224 26056 19236
rect 24964 19196 26056 19224
rect 26050 19184 26056 19196
rect 26108 19224 26114 19236
rect 26160 19224 26188 19332
rect 26421 19329 26433 19332
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 26694 19320 26700 19372
rect 26752 19360 26758 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26752 19332 26985 19360
rect 26752 19320 26758 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 27062 19320 27068 19372
rect 27120 19360 27126 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 27120 19332 27169 19360
rect 27120 19320 27126 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27522 19320 27528 19372
rect 27580 19360 27586 19372
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 27580 19332 27629 19360
rect 27580 19320 27586 19332
rect 27617 19329 27629 19332
rect 27663 19360 27675 19363
rect 28353 19363 28411 19369
rect 28353 19360 28365 19363
rect 27663 19332 28365 19360
rect 27663 19329 27675 19332
rect 27617 19323 27675 19329
rect 28353 19329 28365 19332
rect 28399 19329 28411 19363
rect 28353 19323 28411 19329
rect 27706 19252 27712 19304
rect 27764 19252 27770 19304
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 28074 19292 28080 19304
rect 27939 19264 28080 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 28166 19252 28172 19304
rect 28224 19252 28230 19304
rect 26108 19196 26188 19224
rect 27724 19224 27752 19252
rect 28184 19224 28212 19252
rect 27724 19196 28212 19224
rect 26108 19184 26114 19196
rect 21284 19128 21864 19156
rect 21177 19119 21235 19125
rect 23934 19116 23940 19168
rect 23992 19116 23998 19168
rect 24854 19116 24860 19168
rect 24912 19116 24918 19168
rect 25590 19116 25596 19168
rect 25648 19116 25654 19168
rect 26326 19116 26332 19168
rect 26384 19116 26390 19168
rect 26510 19116 26516 19168
rect 26568 19116 26574 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 2222 18912 2228 18964
rect 2280 18912 2286 18964
rect 5445 18955 5503 18961
rect 5445 18921 5457 18955
rect 5491 18952 5503 18955
rect 6181 18955 6239 18961
rect 6181 18952 6193 18955
rect 5491 18924 6193 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 6181 18921 6193 18924
rect 6227 18952 6239 18955
rect 6454 18952 6460 18964
rect 6227 18924 6460 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 9033 18955 9091 18961
rect 9033 18921 9045 18955
rect 9079 18921 9091 18955
rect 9033 18915 9091 18921
rect 10229 18955 10287 18961
rect 10229 18921 10241 18955
rect 10275 18952 10287 18955
rect 10318 18952 10324 18964
rect 10275 18924 10324 18952
rect 10275 18921 10287 18924
rect 10229 18915 10287 18921
rect 4525 18887 4583 18893
rect 4525 18853 4537 18887
rect 4571 18884 4583 18887
rect 9048 18884 9076 18915
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 10502 18912 10508 18964
rect 10560 18912 10566 18964
rect 10965 18955 11023 18961
rect 10965 18921 10977 18955
rect 11011 18952 11023 18955
rect 11790 18952 11796 18964
rect 11011 18924 11796 18952
rect 11011 18921 11023 18924
rect 10965 18915 11023 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 12434 18912 12440 18964
rect 12492 18912 12498 18964
rect 13078 18912 13084 18964
rect 13136 18912 13142 18964
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 14458 18952 14464 18964
rect 14139 18924 14464 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 17862 18952 17868 18964
rect 17420 18924 17868 18952
rect 10520 18884 10548 18912
rect 4571 18856 5028 18884
rect 9048 18856 10548 18884
rect 4571 18853 4583 18856
rect 4525 18847 4583 18853
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18816 1731 18819
rect 2866 18816 2872 18828
rect 1719 18788 2872 18816
rect 1719 18785 1731 18788
rect 1673 18779 1731 18785
rect 2866 18776 2872 18788
rect 2924 18816 2930 18828
rect 5000 18825 5028 18856
rect 4985 18819 5043 18825
rect 2924 18788 3464 18816
rect 2924 18776 2930 18788
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2455 18720 2697 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 2685 18717 2697 18720
rect 2731 18748 2743 18751
rect 2774 18748 2780 18760
rect 2731 18720 2780 18748
rect 2731 18717 2743 18720
rect 2685 18711 2743 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 3436 18757 3464 18788
rect 4985 18785 4997 18819
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 5166 18776 5172 18828
rect 5224 18816 5230 18828
rect 5537 18819 5595 18825
rect 5537 18816 5549 18819
rect 5224 18788 5549 18816
rect 5224 18776 5230 18788
rect 5537 18785 5549 18788
rect 5583 18785 5595 18819
rect 5537 18779 5595 18785
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 6604 18788 6653 18816
rect 6604 18776 6610 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 7006 18776 7012 18828
rect 7064 18776 7070 18828
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7147 18788 7573 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7561 18785 7573 18788
rect 7607 18816 7619 18819
rect 7650 18816 7656 18828
rect 7607 18788 7656 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 8938 18776 8944 18828
rect 8996 18816 9002 18828
rect 9769 18819 9827 18825
rect 8996 18788 9720 18816
rect 8996 18776 9002 18788
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 3513 18751 3571 18757
rect 3513 18717 3525 18751
rect 3559 18748 3571 18751
rect 3789 18751 3847 18757
rect 3789 18748 3801 18751
rect 3559 18720 3801 18748
rect 3559 18717 3571 18720
rect 3513 18711 3571 18717
rect 3789 18717 3801 18720
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 3970 18708 3976 18760
rect 4028 18708 4034 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 4890 18748 4896 18760
rect 4847 18720 4896 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 3329 18683 3387 18689
rect 3329 18680 3341 18683
rect 2372 18652 3341 18680
rect 2372 18640 2378 18652
rect 3329 18649 3341 18652
rect 3375 18649 3387 18683
rect 4724 18680 4752 18711
rect 4890 18708 4896 18720
rect 4948 18708 4954 18760
rect 5442 18708 5448 18760
rect 5500 18708 5506 18760
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 5460 18680 5488 18708
rect 4724 18652 5488 18680
rect 3329 18643 3387 18649
rect 2498 18572 2504 18624
rect 2556 18572 2562 18624
rect 4430 18572 4436 18624
rect 4488 18572 4494 18624
rect 6472 18612 6500 18711
rect 7024 18680 7052 18776
rect 8570 18708 8576 18760
rect 8628 18708 8634 18760
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8904 18720 9229 18748
rect 8904 18708 8910 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9692 18748 9720 18788
rect 9769 18785 9781 18819
rect 9815 18816 9827 18819
rect 9858 18816 9864 18828
rect 9815 18788 9864 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 12805 18819 12863 18825
rect 12805 18785 12817 18819
rect 12851 18816 12863 18819
rect 13449 18819 13507 18825
rect 13449 18816 13461 18819
rect 12851 18788 13461 18816
rect 12851 18785 12863 18788
rect 12805 18779 12863 18785
rect 13449 18785 13461 18788
rect 13495 18785 13507 18819
rect 13449 18779 13507 18785
rect 10134 18748 10140 18760
rect 9692 18720 10140 18748
rect 9585 18711 9643 18717
rect 7285 18683 7343 18689
rect 7285 18680 7297 18683
rect 7024 18652 7297 18680
rect 7285 18649 7297 18652
rect 7331 18649 7343 18683
rect 7285 18643 7343 18649
rect 7377 18683 7435 18689
rect 7377 18649 7389 18683
rect 7423 18680 7435 18683
rect 7558 18680 7564 18692
rect 7423 18652 7564 18680
rect 7423 18649 7435 18652
rect 7377 18643 7435 18649
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 9324 18680 9352 18711
rect 8496 18652 9352 18680
rect 9600 18680 9628 18711
rect 10134 18708 10140 18720
rect 10192 18748 10198 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 10192 18720 10333 18748
rect 10192 18708 10198 18720
rect 10321 18717 10333 18720
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 11112 18720 11161 18748
rect 11112 18708 11118 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 11885 18751 11943 18757
rect 11885 18717 11897 18751
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 9858 18680 9864 18692
rect 9600 18652 9864 18680
rect 8496 18624 8524 18652
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 11701 18683 11759 18689
rect 11701 18649 11713 18683
rect 11747 18680 11759 18683
rect 11790 18680 11796 18692
rect 11747 18652 11796 18680
rect 11747 18649 11759 18652
rect 11701 18643 11759 18649
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 7466 18612 7472 18624
rect 6472 18584 7472 18612
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 8386 18572 8392 18624
rect 8444 18572 8450 18624
rect 8478 18572 8484 18624
rect 8536 18572 8542 18624
rect 9401 18615 9459 18621
rect 9401 18581 9413 18615
rect 9447 18612 9459 18615
rect 10778 18612 10784 18624
rect 9447 18584 10784 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11900 18612 11928 18711
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12618 18708 12624 18760
rect 12676 18708 12682 18760
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 13817 18751 13875 18757
rect 13817 18748 13829 18751
rect 13780 18720 13829 18748
rect 13780 18708 13786 18720
rect 13817 18717 13829 18720
rect 13863 18717 13875 18751
rect 13817 18711 13875 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14292 18680 14320 18711
rect 14642 18708 14648 18760
rect 14700 18748 14706 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 14700 18720 15393 18748
rect 14700 18708 14706 18720
rect 15381 18717 15393 18720
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 13648 18652 14320 18680
rect 15396 18680 15424 18711
rect 15562 18708 15568 18760
rect 15620 18708 15626 18760
rect 17420 18757 17448 18924
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18874 18912 18880 18964
rect 18932 18912 18938 18964
rect 19628 18924 23428 18952
rect 19628 18825 19656 18924
rect 23400 18884 23428 18924
rect 23474 18912 23480 18964
rect 23532 18912 23538 18964
rect 24762 18952 24768 18964
rect 23584 18924 24768 18952
rect 23584 18884 23612 18924
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 25501 18955 25559 18961
rect 25501 18952 25513 18955
rect 24912 18924 25513 18952
rect 24912 18912 24918 18924
rect 25501 18921 25513 18924
rect 25547 18921 25559 18955
rect 25501 18915 25559 18921
rect 20456 18856 21128 18884
rect 23400 18856 23612 18884
rect 24213 18887 24271 18893
rect 20456 18828 20484 18856
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 20438 18776 20444 18828
rect 20496 18776 20502 18828
rect 20898 18776 20904 18828
rect 20956 18776 20962 18828
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17586 18748 17592 18760
rect 17543 18720 17592 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 17764 18751 17822 18757
rect 17764 18717 17776 18751
rect 17810 18748 17822 18751
rect 18690 18748 18696 18760
rect 17810 18720 18696 18748
rect 17810 18717 17822 18720
rect 17764 18711 17822 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19444 18680 19472 18711
rect 20990 18708 20996 18760
rect 21048 18708 21054 18760
rect 21008 18680 21036 18708
rect 15396 18652 19380 18680
rect 19444 18652 21036 18680
rect 21100 18680 21128 18856
rect 24213 18853 24225 18887
rect 24259 18884 24271 18887
rect 25038 18884 25044 18896
rect 24259 18856 25044 18884
rect 24259 18853 24271 18856
rect 24213 18847 24271 18853
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 23569 18819 23627 18825
rect 23569 18816 23581 18819
rect 22388 18788 23581 18816
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18748 21419 18751
rect 21450 18748 21456 18760
rect 21407 18720 21456 18748
rect 21407 18717 21419 18720
rect 21361 18711 21419 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 22388 18748 22416 18788
rect 23569 18785 23581 18788
rect 23615 18785 23627 18819
rect 23569 18779 23627 18785
rect 24486 18776 24492 18828
rect 24544 18816 24550 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 24544 18788 25145 18816
rect 24544 18776 24550 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25516 18816 25544 18915
rect 26326 18912 26332 18964
rect 26384 18912 26390 18964
rect 26344 18884 26372 18912
rect 28353 18887 28411 18893
rect 28353 18884 28365 18887
rect 26344 18856 26648 18884
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 25516 18788 25881 18816
rect 25133 18779 25191 18785
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 25869 18779 25927 18785
rect 26053 18819 26111 18825
rect 26053 18785 26065 18819
rect 26099 18816 26111 18819
rect 26510 18816 26516 18828
rect 26099 18788 26516 18816
rect 26099 18785 26111 18788
rect 26053 18779 26111 18785
rect 26510 18776 26516 18788
rect 26568 18776 26574 18828
rect 26620 18825 26648 18856
rect 26804 18856 28365 18884
rect 26804 18825 26832 18856
rect 28353 18853 28365 18856
rect 28399 18853 28411 18887
rect 28353 18847 28411 18853
rect 26605 18819 26663 18825
rect 26605 18785 26617 18819
rect 26651 18785 26663 18819
rect 26605 18779 26663 18785
rect 26789 18819 26847 18825
rect 26789 18785 26801 18819
rect 26835 18785 26847 18819
rect 26789 18779 26847 18785
rect 27433 18819 27491 18825
rect 27433 18785 27445 18819
rect 27479 18816 27491 18819
rect 27522 18816 27528 18828
rect 27479 18788 27528 18816
rect 27479 18785 27491 18788
rect 27433 18779 27491 18785
rect 27522 18776 27528 18788
rect 27580 18776 27586 18828
rect 27617 18819 27675 18825
rect 27617 18785 27629 18819
rect 27663 18816 27675 18819
rect 27982 18816 27988 18828
rect 27663 18788 27988 18816
rect 27663 18785 27675 18788
rect 27617 18779 27675 18785
rect 27982 18776 27988 18788
rect 28040 18776 28046 18828
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 21560 18720 22416 18748
rect 22756 18720 22845 18748
rect 21560 18680 21588 18720
rect 21100 18652 21588 18680
rect 21628 18683 21686 18689
rect 11974 18612 11980 18624
rect 11112 18584 11980 18612
rect 11112 18572 11118 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 13648 18621 13676 18652
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 15286 18612 15292 18624
rect 13872 18584 15292 18612
rect 13872 18572 13878 18584
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 16022 18572 16028 18624
rect 16080 18572 16086 18624
rect 17218 18572 17224 18624
rect 17276 18572 17282 18624
rect 19352 18612 19380 18652
rect 21628 18649 21640 18683
rect 21674 18680 21686 18683
rect 22462 18680 22468 18692
rect 21674 18652 22468 18680
rect 21674 18649 21686 18652
rect 21628 18643 21686 18649
rect 22462 18640 22468 18652
rect 22520 18640 22526 18692
rect 22756 18624 22784 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23750 18708 23756 18760
rect 23808 18708 23814 18760
rect 24397 18751 24455 18757
rect 24397 18717 24409 18751
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24412 18680 24440 18711
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 25314 18708 25320 18760
rect 25372 18708 25378 18760
rect 28534 18708 28540 18760
rect 28592 18708 28598 18760
rect 22848 18652 24440 18680
rect 22848 18624 22876 18652
rect 21266 18612 21272 18624
rect 19352 18584 21272 18612
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 22830 18572 22836 18624
rect 22888 18572 22894 18624
rect 27246 18572 27252 18624
rect 27304 18572 27310 18624
rect 28074 18572 28080 18624
rect 28132 18572 28138 18624
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 2314 18368 2320 18420
rect 2372 18368 2378 18420
rect 2498 18368 2504 18420
rect 2556 18368 2562 18420
rect 2777 18411 2835 18417
rect 2777 18377 2789 18411
rect 2823 18408 2835 18411
rect 2866 18408 2872 18420
rect 2823 18380 2872 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 3970 18408 3976 18420
rect 3835 18380 3976 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4430 18368 4436 18420
rect 4488 18368 4494 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5718 18408 5724 18420
rect 5123 18380 5724 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 6696 18380 7052 18408
rect 6696 18368 6702 18380
rect 1664 18343 1722 18349
rect 1664 18309 1676 18343
rect 1710 18340 1722 18343
rect 2332 18340 2360 18368
rect 1710 18312 2360 18340
rect 1710 18309 1722 18312
rect 1664 18303 1722 18309
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 2516 18272 2544 18368
rect 3605 18343 3663 18349
rect 3605 18309 3617 18343
rect 3651 18340 3663 18343
rect 3651 18312 4016 18340
rect 3651 18309 3663 18312
rect 3605 18303 3663 18309
rect 2961 18275 3019 18281
rect 2961 18272 2973 18275
rect 2516 18244 2973 18272
rect 2961 18241 2973 18244
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 3988 18281 4016 18312
rect 3973 18275 4031 18281
rect 3973 18241 3985 18275
rect 4019 18272 4031 18275
rect 4448 18272 4476 18368
rect 4617 18343 4675 18349
rect 4617 18309 4629 18343
rect 4663 18340 4675 18343
rect 4798 18340 4804 18352
rect 4663 18312 4804 18340
rect 4663 18309 4675 18312
rect 4617 18303 4675 18309
rect 4798 18300 4804 18312
rect 4856 18340 4862 18352
rect 5166 18340 5172 18352
rect 4856 18312 5172 18340
rect 4856 18300 4862 18312
rect 5166 18300 5172 18312
rect 5224 18300 5230 18352
rect 7024 18340 7052 18380
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 7524 18380 8401 18408
rect 7524 18368 7530 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 8938 18368 8944 18420
rect 8996 18368 9002 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 9585 18411 9643 18417
rect 9585 18408 9597 18411
rect 9364 18380 9597 18408
rect 9364 18368 9370 18380
rect 9585 18377 9597 18380
rect 9631 18377 9643 18411
rect 9585 18371 9643 18377
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 10376 18380 10609 18408
rect 10376 18368 10382 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 10778 18368 10784 18420
rect 10836 18368 10842 18420
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 12066 18408 12072 18420
rect 11655 18380 12072 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12529 18411 12587 18417
rect 12529 18408 12541 18411
rect 12492 18380 12541 18408
rect 12492 18368 12498 18380
rect 12529 18377 12541 18380
rect 12575 18377 12587 18411
rect 12529 18371 12587 18377
rect 13170 18368 13176 18420
rect 13228 18368 13234 18420
rect 14921 18411 14979 18417
rect 14921 18377 14933 18411
rect 14967 18408 14979 18411
rect 15562 18408 15568 18420
rect 14967 18380 15568 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 16080 18380 16129 18408
rect 16080 18368 16086 18380
rect 16117 18377 16129 18380
rect 16163 18377 16175 18411
rect 16117 18371 16175 18377
rect 17218 18368 17224 18420
rect 17276 18368 17282 18420
rect 17310 18368 17316 18420
rect 17368 18368 17374 18420
rect 17862 18368 17868 18420
rect 17920 18368 17926 18420
rect 19886 18408 19892 18420
rect 17972 18380 19892 18408
rect 8662 18340 8668 18352
rect 7024 18312 7130 18340
rect 7944 18312 8668 18340
rect 4019 18244 4476 18272
rect 4709 18275 4767 18281
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4755 18244 4936 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 3142 18164 3148 18216
rect 3200 18164 3206 18216
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4801 18207 4859 18213
rect 4801 18204 4813 18207
rect 4203 18176 4813 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4801 18173 4813 18176
rect 4847 18173 4859 18207
rect 4801 18167 4859 18173
rect 3970 18096 3976 18148
rect 4028 18136 4034 18148
rect 4908 18136 4936 18244
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 5442 18232 5448 18284
rect 5500 18232 5506 18284
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6144 18244 6745 18272
rect 6144 18232 6150 18244
rect 6733 18241 6745 18244
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 7944 18272 7972 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 7708 18244 7972 18272
rect 8205 18275 8263 18281
rect 7708 18232 7714 18244
rect 8205 18241 8217 18275
rect 8251 18241 8263 18275
rect 8956 18272 8984 18368
rect 10796 18340 10824 18368
rect 10796 18312 12112 18340
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 8956 18244 9505 18272
rect 8205 18235 8263 18241
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18204 5595 18207
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5583 18176 6377 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 7190 18204 7196 18216
rect 6365 18167 6423 18173
rect 6472 18176 7196 18204
rect 4028 18108 4936 18136
rect 6089 18139 6147 18145
rect 4028 18096 4034 18108
rect 6089 18105 6101 18139
rect 6135 18136 6147 18139
rect 6472 18136 6500 18176
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 6135 18108 6500 18136
rect 6135 18105 6147 18108
rect 6089 18099 6147 18105
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 8220 18068 8248 18235
rect 9950 18232 9956 18284
rect 10008 18232 10014 18284
rect 10226 18272 10232 18284
rect 10060 18244 10232 18272
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 8772 18136 8800 18167
rect 8938 18164 8944 18216
rect 8996 18164 9002 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 9180 18176 9413 18204
rect 9180 18164 9186 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 9950 18136 9956 18148
rect 8772 18108 9956 18136
rect 9950 18096 9956 18108
rect 10008 18136 10014 18148
rect 10060 18136 10088 18244
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10652 18244 10701 18272
rect 10652 18232 10658 18244
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 12084 18281 12112 18312
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 13780 18312 15240 18340
rect 13780 18300 13786 18312
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11204 18244 11345 18272
rect 11204 18232 11210 18244
rect 11333 18241 11345 18244
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18241 11851 18275
rect 11793 18235 11851 18241
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18241 12127 18275
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12069 18235 12127 18241
rect 12452 18244 13093 18272
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10183 18176 10793 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 11808 18204 11836 18235
rect 12452 18216 12480 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 15212 18281 15240 18312
rect 14829 18275 14887 18281
rect 14829 18272 14841 18275
rect 13688 18244 14841 18272
rect 13688 18232 13694 18244
rect 14829 18241 14841 18244
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18272 15347 18275
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15335 18244 15669 18272
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 10781 18167 10839 18173
rect 11164 18176 11836 18204
rect 11164 18145 11192 18176
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 12158 18204 12164 18216
rect 11940 18176 12164 18204
rect 11940 18164 11946 18176
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 12434 18164 12440 18216
rect 12492 18164 12498 18216
rect 15120 18204 15148 18235
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16264 18244 16681 18272
rect 16264 18232 16270 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 17236 18272 17264 18368
rect 17589 18275 17647 18281
rect 17589 18272 17601 18275
rect 17236 18244 17601 18272
rect 16669 18235 16727 18241
rect 17589 18241 17601 18244
rect 17635 18241 17647 18275
rect 17589 18235 17647 18241
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18272 17739 18275
rect 17880 18272 17908 18368
rect 17727 18244 17908 18272
rect 17972 18272 18000 18380
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 21361 18411 21419 18417
rect 21048 18380 21312 18408
rect 21048 18368 21054 18380
rect 19334 18300 19340 18352
rect 19392 18300 19398 18352
rect 21177 18343 21235 18349
rect 21177 18340 21189 18343
rect 19812 18312 21189 18340
rect 19812 18281 19840 18312
rect 21177 18309 21189 18312
rect 21223 18309 21235 18343
rect 21284 18340 21312 18380
rect 21361 18377 21373 18411
rect 21407 18408 21419 18411
rect 22186 18408 22192 18420
rect 21407 18380 22192 18408
rect 21407 18377 21419 18380
rect 21361 18371 21419 18377
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 22278 18368 22284 18420
rect 22336 18368 22342 18420
rect 22462 18368 22468 18420
rect 22520 18368 22526 18420
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 23937 18411 23995 18417
rect 23937 18408 23949 18411
rect 23808 18380 23949 18408
rect 23808 18368 23814 18380
rect 23937 18377 23949 18380
rect 23983 18377 23995 18411
rect 23937 18371 23995 18377
rect 24213 18411 24271 18417
rect 24213 18377 24225 18411
rect 24259 18408 24271 18411
rect 24394 18408 24400 18420
rect 24259 18380 24400 18408
rect 24259 18377 24271 18380
rect 24213 18371 24271 18377
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 24636 18380 24869 18408
rect 24636 18368 24642 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 24946 18368 24952 18420
rect 25004 18368 25010 18420
rect 25133 18411 25191 18417
rect 25133 18377 25145 18411
rect 25179 18408 25191 18411
rect 25314 18408 25320 18420
rect 25179 18380 25320 18408
rect 25179 18377 25191 18380
rect 25133 18371 25191 18377
rect 25314 18368 25320 18380
rect 25372 18368 25378 18420
rect 25590 18368 25596 18420
rect 25648 18408 25654 18420
rect 25648 18380 25728 18408
rect 25648 18368 25654 18380
rect 22296 18340 22324 18368
rect 24302 18340 24308 18352
rect 21284 18312 22324 18340
rect 24136 18312 24308 18340
rect 21177 18303 21235 18309
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 17972 18244 18337 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18272 20591 18275
rect 20806 18272 20812 18284
rect 20579 18244 20812 18272
rect 20579 18241 20591 18244
rect 20533 18235 20591 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 20956 18244 21097 18272
rect 20956 18232 20962 18244
rect 21085 18241 21097 18244
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 21545 18275 21603 18281
rect 21545 18241 21557 18275
rect 21591 18272 21603 18275
rect 21634 18272 21640 18284
rect 21591 18244 21640 18272
rect 21591 18241 21603 18244
rect 21545 18235 21603 18241
rect 21634 18232 21640 18244
rect 21692 18272 21698 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21692 18244 21833 18272
rect 21692 18232 21698 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22738 18272 22744 18284
rect 22152 18244 22744 18272
rect 22152 18232 22158 18244
rect 22738 18232 22744 18244
rect 22796 18272 22802 18284
rect 24136 18281 24164 18312
rect 24302 18300 24308 18312
rect 24360 18300 24366 18352
rect 24964 18340 24992 18368
rect 25700 18349 25728 18380
rect 28074 18368 28080 18420
rect 28132 18408 28138 18420
rect 28353 18411 28411 18417
rect 28353 18408 28365 18411
rect 28132 18380 28365 18408
rect 28132 18368 28138 18380
rect 28353 18377 28365 18380
rect 28399 18377 28411 18411
rect 28353 18371 28411 18377
rect 24412 18312 24992 18340
rect 25676 18343 25734 18349
rect 24412 18281 24440 18312
rect 25676 18309 25688 18343
rect 25722 18309 25734 18343
rect 25676 18303 25734 18309
rect 22925 18275 22983 18281
rect 22925 18272 22937 18275
rect 22796 18244 22937 18272
rect 22796 18232 22802 18244
rect 22925 18241 22937 18244
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 24670 18232 24676 18284
rect 24728 18232 24734 18284
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18272 24823 18275
rect 24946 18272 24952 18284
rect 24811 18244 24952 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 24946 18232 24952 18244
rect 25004 18272 25010 18284
rect 25041 18275 25099 18281
rect 25041 18272 25053 18275
rect 25004 18244 25053 18272
rect 25004 18232 25010 18244
rect 25041 18241 25053 18244
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 27065 18275 27123 18281
rect 27065 18241 27077 18275
rect 27111 18272 27123 18275
rect 27154 18272 27160 18284
rect 27111 18244 27160 18272
rect 27111 18241 27123 18244
rect 27065 18235 27123 18241
rect 13004 18176 13860 18204
rect 10008 18108 10088 18136
rect 11149 18139 11207 18145
rect 10008 18096 10014 18108
rect 11149 18105 11161 18139
rect 11195 18105 11207 18139
rect 11149 18099 11207 18105
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 13004 18136 13032 18176
rect 13832 18148 13860 18176
rect 14660 18176 15148 18204
rect 15473 18207 15531 18213
rect 12032 18108 13032 18136
rect 13096 18108 13308 18136
rect 12032 18096 12038 18108
rect 6788 18040 8248 18068
rect 6788 18028 6794 18040
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 13096 18068 13124 18108
rect 9088 18040 13124 18068
rect 13280 18068 13308 18108
rect 13814 18096 13820 18148
rect 13872 18096 13878 18148
rect 14660 18145 14688 18176
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18105 14703 18139
rect 14645 18099 14703 18105
rect 15488 18068 15516 18167
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16224 18204 16252 18232
rect 15896 18176 16252 18204
rect 15896 18164 15902 18176
rect 17954 18164 17960 18216
rect 18012 18164 18018 18216
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 17405 18139 17463 18145
rect 17405 18105 17417 18139
rect 17451 18136 17463 18139
rect 18046 18136 18052 18148
rect 17451 18108 18052 18136
rect 17451 18105 17463 18108
rect 17405 18099 17463 18105
rect 18046 18096 18052 18108
rect 18104 18096 18110 18148
rect 19981 18139 20039 18145
rect 19981 18105 19993 18139
rect 20027 18136 20039 18139
rect 20364 18136 20392 18167
rect 23198 18164 23204 18216
rect 23256 18164 23262 18216
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 23750 18204 23756 18216
rect 23431 18176 23756 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 23934 18164 23940 18216
rect 23992 18204 23998 18216
rect 25130 18204 25136 18216
rect 23992 18176 25136 18204
rect 23992 18164 23998 18176
rect 25130 18164 25136 18176
rect 25188 18204 25194 18216
rect 25409 18207 25467 18213
rect 25409 18204 25421 18207
rect 25188 18176 25421 18204
rect 25188 18164 25194 18176
rect 25409 18173 25421 18176
rect 25455 18173 25467 18207
rect 25409 18167 25467 18173
rect 20027 18108 20392 18136
rect 26789 18139 26847 18145
rect 20027 18105 20039 18108
rect 19981 18099 20039 18105
rect 26789 18105 26801 18139
rect 26835 18136 26847 18139
rect 27080 18136 27108 18235
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27709 18275 27767 18281
rect 27709 18241 27721 18275
rect 27755 18272 27767 18275
rect 28350 18272 28356 18284
rect 27755 18244 28356 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 27890 18164 27896 18216
rect 27948 18164 27954 18216
rect 26835 18108 27108 18136
rect 26835 18105 26847 18108
rect 26789 18099 26847 18105
rect 13280 18040 15516 18068
rect 16301 18071 16359 18077
rect 9088 18028 9094 18040
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16482 18068 16488 18080
rect 16347 18040 16488 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 17770 18028 17776 18080
rect 17828 18028 17834 18080
rect 22741 18071 22799 18077
rect 22741 18037 22753 18071
rect 22787 18068 22799 18071
rect 23474 18068 23480 18080
rect 22787 18040 23480 18068
rect 22787 18037 22799 18040
rect 22741 18031 22799 18037
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 23842 18028 23848 18080
rect 23900 18028 23906 18080
rect 24486 18028 24492 18080
rect 24544 18028 24550 18080
rect 26878 18028 26884 18080
rect 26936 18068 26942 18080
rect 27617 18071 27675 18077
rect 27617 18068 27629 18071
rect 26936 18040 27629 18068
rect 26936 18028 26942 18040
rect 27617 18037 27629 18040
rect 27663 18037 27675 18071
rect 27617 18031 27675 18037
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 2774 17824 2780 17876
rect 2832 17824 2838 17876
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3142 17864 3148 17876
rect 3007 17836 3148 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 4798 17824 4804 17876
rect 4856 17824 4862 17876
rect 5994 17824 6000 17876
rect 6052 17824 6058 17876
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6638 17864 6644 17876
rect 6595 17836 6644 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 6788 17836 6837 17864
rect 6788 17824 6794 17836
rect 6825 17833 6837 17836
rect 6871 17833 6883 17867
rect 6825 17827 6883 17833
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7282 17864 7288 17876
rect 7055 17836 7288 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 8938 17864 8944 17876
rect 7423 17836 8944 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 8938 17824 8944 17836
rect 8996 17824 9002 17876
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 9309 17867 9367 17873
rect 9309 17864 9321 17867
rect 9180 17836 9321 17864
rect 9180 17824 9186 17836
rect 9309 17833 9321 17836
rect 9355 17833 9367 17867
rect 10042 17864 10048 17876
rect 9309 17827 9367 17833
rect 9416 17836 10048 17864
rect 4893 17799 4951 17805
rect 4893 17796 4905 17799
rect 4356 17768 4905 17796
rect 1394 17688 1400 17740
rect 1452 17688 1458 17740
rect 4356 17737 4384 17768
rect 4893 17765 4905 17768
rect 4939 17765 4951 17799
rect 6012 17796 6040 17824
rect 8478 17796 8484 17808
rect 6012 17768 8484 17796
rect 4893 17759 4951 17765
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17697 4399 17731
rect 4341 17691 4399 17697
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 3602 17660 3608 17672
rect 3191 17632 3608 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 4028 17632 4077 17660
rect 4028 17620 4034 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4246 17660 4252 17672
rect 4203 17632 4252 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 1664 17595 1722 17601
rect 1664 17561 1676 17595
rect 1710 17592 1722 17595
rect 2314 17592 2320 17604
rect 1710 17564 2320 17592
rect 1710 17561 1722 17564
rect 1664 17555 1722 17561
rect 2314 17552 2320 17564
rect 2372 17552 2378 17604
rect 5092 17592 5120 17623
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6328 17632 6469 17660
rect 6328 17620 6334 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 3896 17564 5120 17592
rect 6656 17592 6684 17623
rect 6730 17620 6736 17672
rect 6788 17620 6794 17672
rect 7006 17592 7012 17604
rect 6656 17564 7012 17592
rect 3896 17533 3924 17564
rect 7006 17552 7012 17564
rect 7064 17552 7070 17604
rect 7116 17592 7144 17768
rect 8478 17756 8484 17768
rect 8536 17756 8542 17808
rect 8754 17756 8760 17808
rect 8812 17756 8818 17808
rect 7208 17700 8248 17728
rect 7208 17669 7236 17700
rect 7760 17669 7788 17700
rect 8220 17672 8248 17700
rect 8294 17688 8300 17740
rect 8352 17688 8358 17740
rect 8386 17688 8392 17740
rect 8444 17728 8450 17740
rect 9125 17731 9183 17737
rect 9125 17728 9137 17731
rect 8444 17700 9137 17728
rect 8444 17688 8450 17700
rect 9125 17697 9137 17700
rect 9171 17697 9183 17731
rect 9125 17691 9183 17697
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17629 8079 17663
rect 8021 17623 8079 17629
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 7300 17592 7328 17623
rect 8036 17592 8064 17623
rect 7116 17564 7328 17592
rect 7576 17564 8064 17592
rect 8128 17592 8156 17623
rect 8202 17620 8208 17672
rect 8260 17620 8266 17672
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9416 17660 9444 17836
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 15654 17864 15660 17876
rect 10244 17836 15660 17864
rect 9953 17799 10011 17805
rect 9953 17765 9965 17799
rect 9999 17765 10011 17799
rect 9953 17759 10011 17765
rect 8987 17632 9444 17660
rect 9861 17663 9919 17669
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9861 17629 9873 17663
rect 9907 17660 9919 17663
rect 9968 17660 9996 17759
rect 9907 17632 9996 17660
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 10134 17620 10140 17672
rect 10192 17620 10198 17672
rect 10244 17604 10272 17836
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 19334 17824 19340 17876
rect 19392 17824 19398 17876
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 21542 17864 21548 17876
rect 21131 17836 21548 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24029 17867 24087 17873
rect 24029 17864 24041 17867
rect 23808 17836 24041 17864
rect 23808 17824 23814 17836
rect 24029 17833 24041 17836
rect 24075 17833 24087 17867
rect 24029 17827 24087 17833
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 24912 17836 25881 17864
rect 24912 17824 24918 17836
rect 25869 17833 25881 17836
rect 25915 17833 25927 17867
rect 25869 17827 25927 17833
rect 27246 17824 27252 17876
rect 27304 17824 27310 17876
rect 11330 17756 11336 17808
rect 11388 17796 11394 17808
rect 13998 17796 14004 17808
rect 11388 17768 14004 17796
rect 11388 17756 11394 17768
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 14737 17799 14795 17805
rect 14737 17765 14749 17799
rect 14783 17796 14795 17799
rect 15197 17799 15255 17805
rect 15197 17796 15209 17799
rect 14783 17768 15209 17796
rect 14783 17765 14795 17768
rect 14737 17759 14795 17765
rect 15197 17765 15209 17768
rect 15243 17765 15255 17799
rect 15197 17759 15255 17765
rect 16577 17799 16635 17805
rect 16577 17765 16589 17799
rect 16623 17796 16635 17799
rect 17037 17799 17095 17805
rect 17037 17796 17049 17799
rect 16623 17768 17049 17796
rect 16623 17765 16635 17768
rect 16577 17759 16635 17765
rect 17037 17765 17049 17768
rect 17083 17765 17095 17799
rect 17037 17759 17095 17765
rect 18049 17799 18107 17805
rect 18049 17765 18061 17799
rect 18095 17796 18107 17799
rect 18138 17796 18144 17808
rect 18095 17768 18144 17796
rect 18095 17765 18107 17768
rect 18049 17759 18107 17765
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17697 10379 17731
rect 12710 17728 12716 17740
rect 10321 17691 10379 17697
rect 11348 17700 12716 17728
rect 10336 17660 10364 17691
rect 11348 17660 11376 17700
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17728 13875 17731
rect 15013 17731 15071 17737
rect 15013 17728 15025 17731
rect 13863 17700 15025 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 15013 17697 15025 17700
rect 15059 17697 15071 17731
rect 15212 17728 15240 17759
rect 15933 17731 15991 17737
rect 15933 17728 15945 17731
rect 15212 17700 15945 17728
rect 15013 17691 15071 17697
rect 15933 17697 15945 17700
rect 15979 17697 15991 17731
rect 15933 17691 15991 17697
rect 16022 17688 16028 17740
rect 16080 17728 16086 17740
rect 16080 17700 16344 17728
rect 16080 17688 16086 17700
rect 10336 17632 11376 17660
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 12434 17660 12440 17672
rect 11664 17632 12440 17660
rect 11664 17620 11670 17632
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 13633 17639 13691 17645
rect 13633 17605 13645 17639
rect 13679 17605 13691 17639
rect 13722 17620 13728 17672
rect 13780 17620 13786 17672
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 14056 17632 14105 17660
rect 14056 17620 14062 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14274 17620 14280 17672
rect 14332 17620 14338 17672
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14792 17632 14841 17660
rect 14792 17620 14798 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16114 17620 16120 17672
rect 16172 17620 16178 17672
rect 16316 17660 16344 17700
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 16853 17731 16911 17737
rect 16853 17728 16865 17731
rect 16540 17700 16865 17728
rect 16540 17688 16546 17700
rect 16853 17697 16865 17700
rect 16899 17697 16911 17731
rect 17052 17728 17080 17759
rect 18138 17756 18144 17768
rect 18196 17796 18202 17808
rect 21637 17799 21695 17805
rect 18196 17768 18644 17796
rect 18196 17756 18202 17768
rect 18616 17737 18644 17768
rect 21637 17765 21649 17799
rect 21683 17765 21695 17799
rect 21637 17759 21695 17765
rect 21913 17799 21971 17805
rect 21913 17765 21925 17799
rect 21959 17796 21971 17799
rect 22833 17799 22891 17805
rect 21959 17768 22416 17796
rect 21959 17765 21971 17768
rect 21913 17759 21971 17765
rect 18325 17731 18383 17737
rect 18325 17728 18337 17731
rect 17052 17700 18337 17728
rect 16853 17691 16911 17697
rect 18325 17697 18337 17700
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17697 18659 17731
rect 21652 17728 21680 17759
rect 22388 17737 22416 17768
rect 22833 17765 22845 17799
rect 22879 17796 22891 17799
rect 23293 17799 23351 17805
rect 23293 17796 23305 17799
rect 22879 17768 23305 17796
rect 22879 17765 22891 17768
rect 22833 17759 22891 17765
rect 23293 17765 23305 17768
rect 23339 17796 23351 17799
rect 23566 17796 23572 17808
rect 23339 17768 23572 17796
rect 23339 17765 23351 17768
rect 23293 17759 23351 17765
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 23842 17756 23848 17808
rect 23900 17756 23906 17808
rect 25777 17799 25835 17805
rect 25777 17765 25789 17799
rect 25823 17796 25835 17799
rect 26326 17796 26332 17808
rect 25823 17768 26332 17796
rect 25823 17765 25835 17768
rect 25777 17759 25835 17765
rect 26326 17756 26332 17768
rect 26384 17796 26390 17808
rect 27264 17796 27292 17824
rect 26384 17768 27292 17796
rect 26384 17756 26390 17768
rect 22373 17731 22431 17737
rect 21652 17700 22140 17728
rect 18601 17691 18659 17697
rect 16669 17663 16727 17669
rect 16669 17660 16681 17663
rect 16316 17632 16681 17660
rect 16669 17629 16681 17632
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19475 17632 19564 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 10226 17592 10232 17604
rect 8128 17564 10232 17592
rect 7576 17533 7604 17564
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 10588 17595 10646 17601
rect 10588 17561 10600 17595
rect 10634 17592 10646 17595
rect 11882 17592 11888 17604
rect 10634 17564 11888 17592
rect 10634 17561 10646 17564
rect 10588 17555 10646 17561
rect 11882 17552 11888 17564
rect 11940 17552 11946 17604
rect 13633 17599 13691 17605
rect 13648 17536 13676 17599
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 15856 17592 15884 17620
rect 15528 17564 15884 17592
rect 15528 17552 15534 17564
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 17276 17564 17509 17592
rect 17276 17552 17282 17564
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 17589 17595 17647 17601
rect 17589 17561 17601 17595
rect 17635 17592 17647 17595
rect 17770 17592 17776 17604
rect 17635 17564 17776 17592
rect 17635 17561 17647 17564
rect 17589 17555 17647 17561
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 18417 17595 18475 17601
rect 18417 17561 18429 17595
rect 18463 17561 18475 17595
rect 18417 17555 18475 17561
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17493 3939 17527
rect 3881 17487 3939 17493
rect 7561 17527 7619 17533
rect 7561 17493 7573 17527
rect 7607 17493 7619 17527
rect 7561 17487 7619 17493
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7800 17496 7849 17524
rect 7800 17484 7806 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 9674 17484 9680 17536
rect 9732 17484 9738 17536
rect 11606 17484 11612 17536
rect 11664 17524 11670 17536
rect 11701 17527 11759 17533
rect 11701 17524 11713 17527
rect 11664 17496 11713 17524
rect 11664 17484 11670 17496
rect 11701 17493 11713 17496
rect 11747 17493 11759 17527
rect 11701 17487 11759 17493
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 13630 17484 13636 17536
rect 13688 17484 13694 17536
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 18432 17524 18460 17555
rect 19536 17536 19564 17632
rect 19610 17620 19616 17672
rect 19668 17660 19674 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19668 17632 19717 17660
rect 19668 17620 19674 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 19972 17663 20030 17669
rect 19972 17629 19984 17663
rect 20018 17660 20030 17663
rect 20530 17660 20536 17672
rect 20018 17632 20536 17660
rect 20018 17629 20030 17632
rect 19972 17623 20030 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 22002 17660 22008 17672
rect 21867 17632 22008 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 22112 17669 22140 17700
rect 22373 17697 22385 17731
rect 22419 17697 22431 17731
rect 23860 17728 23888 17756
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 23860 17700 24409 17728
rect 22373 17691 22431 17697
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 26237 17731 26295 17737
rect 26237 17728 26249 17731
rect 24627 17700 26249 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 26237 17697 26249 17700
rect 26283 17697 26295 17731
rect 26237 17691 26295 17697
rect 26786 17688 26792 17740
rect 26844 17728 26850 17740
rect 26881 17731 26939 17737
rect 26881 17728 26893 17731
rect 26844 17700 26893 17728
rect 26844 17688 26850 17700
rect 26881 17697 26893 17700
rect 26927 17697 26939 17731
rect 26881 17691 26939 17697
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17629 22155 17663
rect 22097 17623 22155 17629
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17629 22983 17663
rect 22925 17623 22983 17629
rect 20714 17552 20720 17604
rect 20772 17592 20778 17604
rect 22204 17592 22232 17623
rect 20772 17564 22232 17592
rect 20772 17552 20778 17564
rect 18104 17496 18460 17524
rect 18104 17484 18110 17496
rect 19518 17484 19524 17536
rect 19576 17484 19582 17536
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 22940 17524 22968 17623
rect 23106 17620 23112 17672
rect 23164 17620 23170 17672
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 23532 17632 23857 17660
rect 23532 17620 23538 17632
rect 23845 17629 23857 17632
rect 23891 17629 23903 17663
rect 23845 17623 23903 17629
rect 23937 17663 23995 17669
rect 23937 17629 23949 17663
rect 23983 17660 23995 17663
rect 24762 17660 24768 17672
rect 23983 17632 24768 17660
rect 23983 17629 23995 17632
rect 23937 17623 23995 17629
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 23952 17592 23980 17623
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25133 17663 25191 17669
rect 25133 17660 25145 17663
rect 25056 17632 25145 17660
rect 23348 17564 23980 17592
rect 23348 17552 23354 17564
rect 25056 17536 25084 17632
rect 25133 17629 25145 17632
rect 25179 17629 25191 17663
rect 25133 17623 25191 17629
rect 25317 17663 25375 17669
rect 25317 17629 25329 17663
rect 25363 17629 25375 17663
rect 25317 17623 25375 17629
rect 25332 17592 25360 17623
rect 26050 17620 26056 17672
rect 26108 17660 26114 17672
rect 26145 17663 26203 17669
rect 26145 17660 26157 17663
rect 26108 17632 26157 17660
rect 26108 17620 26114 17632
rect 26145 17629 26157 17632
rect 26191 17629 26203 17663
rect 26145 17623 26203 17629
rect 26418 17620 26424 17672
rect 26476 17620 26482 17672
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 26234 17592 26240 17604
rect 25332 17564 26240 17592
rect 26234 17552 26240 17564
rect 26292 17552 26298 17604
rect 26602 17552 26608 17604
rect 26660 17552 26666 17604
rect 27430 17552 27436 17604
rect 27488 17592 27494 17604
rect 28552 17592 28580 17623
rect 27488 17564 28580 17592
rect 27488 17552 27494 17564
rect 22244 17496 22968 17524
rect 22244 17484 22250 17496
rect 23658 17484 23664 17536
rect 23716 17484 23722 17536
rect 25038 17484 25044 17536
rect 25096 17484 25102 17536
rect 28350 17484 28356 17536
rect 28408 17484 28414 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 2314 17280 2320 17332
rect 2372 17280 2378 17332
rect 3694 17280 3700 17332
rect 3752 17280 3758 17332
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17289 4767 17323
rect 4709 17283 4767 17289
rect 5997 17323 6055 17329
rect 5997 17289 6009 17323
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 3712 17252 3740 17280
rect 2976 17224 3740 17252
rect 4724 17252 4752 17283
rect 6012 17252 6040 17283
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 6880 17292 9812 17320
rect 6880 17280 6886 17292
rect 4724 17224 5396 17252
rect 6012 17224 7328 17252
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 2976 17193 3004 17224
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 1360 17156 2513 17184
rect 1360 17144 1366 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17153 3019 17187
rect 2961 17147 3019 17153
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 3099 17156 3433 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3421 17153 3433 17156
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17184 4031 17187
rect 4338 17184 4344 17196
rect 4019 17156 4344 17184
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 5368 17193 5396 17224
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2866 17116 2872 17128
rect 1811 17088 2872 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3234 17076 3240 17128
rect 3292 17076 3298 17128
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 4908 17116 4936 17147
rect 6196 17116 6224 17147
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 7300 17193 7328 17224
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 7800 17224 8248 17252
rect 7800 17212 7806 17224
rect 7285 17187 7343 17193
rect 6472 17156 6684 17184
rect 6472 17128 6500 17156
rect 6454 17116 6460 17128
rect 4856 17088 6460 17116
rect 4856 17076 4862 17088
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6656 17116 6684 17156
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7484 17116 7512 17147
rect 7650 17144 7656 17196
rect 7708 17144 7714 17196
rect 8220 17193 8248 17224
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 9784 17252 9812 17292
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 9916 17292 10149 17320
rect 9916 17280 9922 17292
rect 10137 17289 10149 17292
rect 10183 17289 10195 17323
rect 12158 17320 12164 17332
rect 10137 17283 10195 17289
rect 10520 17292 12164 17320
rect 10520 17252 10548 17292
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12250 17280 12256 17332
rect 12308 17320 12314 17332
rect 12529 17323 12587 17329
rect 12308 17292 12434 17320
rect 12308 17280 12314 17292
rect 8444 17224 9628 17252
rect 9784 17224 10548 17252
rect 8444 17212 8450 17224
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8205 17187 8263 17193
rect 7975 17156 8156 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 6656 17088 7512 17116
rect 7668 17116 7696 17144
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7668 17088 8033 17116
rect 6549 17079 6607 17085
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8128 17116 8156 17156
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8352 17156 8892 17184
rect 8352 17144 8358 17156
rect 8312 17116 8340 17144
rect 8864 17128 8892 17156
rect 8128 17088 8340 17116
rect 8021 17079 8079 17085
rect 3881 17051 3939 17057
rect 3881 17017 3893 17051
rect 3927 17048 3939 17051
rect 4246 17048 4252 17060
rect 3927 17020 4252 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 4246 17008 4252 17020
rect 4304 17048 4310 17060
rect 4341 17051 4399 17057
rect 4341 17048 4353 17051
rect 4304 17020 4353 17048
rect 4304 17008 4310 17020
rect 4341 17017 4353 17020
rect 4387 17017 4399 17051
rect 4341 17011 4399 17017
rect 5169 17051 5227 17057
rect 5169 17017 5181 17051
rect 5215 17048 5227 17051
rect 6564 17048 6592 17079
rect 8570 17076 8576 17128
rect 8628 17076 8634 17128
rect 8754 17076 8760 17128
rect 8812 17076 8818 17128
rect 8846 17076 8852 17128
rect 8904 17076 8910 17128
rect 8938 17076 8944 17128
rect 8996 17076 9002 17128
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 7466 17048 7472 17060
rect 5215 17020 6592 17048
rect 6748 17020 7472 17048
rect 5215 17017 5227 17020
rect 5169 17011 5227 17017
rect 6748 16992 6776 17020
rect 7466 17008 7472 17020
rect 7524 17048 7530 17060
rect 7745 17051 7803 17057
rect 7524 17020 7696 17048
rect 7524 17008 7530 17020
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 6730 16980 6736 16992
rect 2823 16952 6736 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 6914 16940 6920 16992
rect 6972 16940 6978 16992
rect 7098 16940 7104 16992
rect 7156 16940 7162 16992
rect 7558 16940 7564 16992
rect 7616 16940 7622 16992
rect 7668 16980 7696 17020
rect 7745 17017 7757 17051
rect 7791 17048 7803 17051
rect 8588 17048 8616 17076
rect 7791 17020 8616 17048
rect 8665 17051 8723 17057
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 8665 17017 8677 17051
rect 8711 17048 8723 17051
rect 9125 17051 9183 17057
rect 9125 17048 9137 17051
rect 8711 17020 9137 17048
rect 8711 17017 8723 17020
rect 8665 17011 8723 17017
rect 9125 17017 9137 17020
rect 9171 17048 9183 17051
rect 9508 17048 9536 17079
rect 9171 17020 9536 17048
rect 9600 17048 9628 17224
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 11330 17252 11336 17264
rect 10652 17224 11336 17252
rect 10652 17212 10658 17224
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10229 17187 10287 17193
rect 10229 17184 10241 17187
rect 10192 17156 10241 17184
rect 10192 17144 10198 17156
rect 10229 17153 10241 17156
rect 10275 17184 10287 17187
rect 11606 17184 11612 17196
rect 10275 17156 11612 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17184 11759 17187
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11747 17156 12081 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12406 17184 12434 17292
rect 12529 17289 12541 17323
rect 12575 17320 12587 17323
rect 12618 17320 12624 17332
rect 12575 17292 12624 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 12618 17280 12624 17292
rect 12676 17320 12682 17332
rect 13265 17323 13323 17329
rect 13265 17320 13277 17323
rect 12676 17292 13277 17320
rect 12676 17280 12682 17292
rect 13265 17289 13277 17292
rect 13311 17289 13323 17323
rect 13265 17283 13323 17289
rect 13446 17280 13452 17332
rect 13504 17280 13510 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14274 17320 14280 17332
rect 14047 17292 14280 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 15654 17280 15660 17332
rect 15712 17280 15718 17332
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16172 17292 16681 17320
rect 16172 17280 16178 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 16669 17283 16727 17289
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17289 17003 17323
rect 16945 17283 17003 17289
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 17954 17320 17960 17332
rect 17911 17292 17960 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 13464 17252 13492 17280
rect 15672 17252 15700 17280
rect 16960 17252 16988 17283
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 20073 17323 20131 17329
rect 20073 17289 20085 17323
rect 20119 17320 20131 17323
rect 21082 17320 21088 17332
rect 20119 17292 21088 17320
rect 20119 17289 20131 17292
rect 20073 17283 20131 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 23106 17320 23112 17332
rect 22695 17292 23112 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23658 17280 23664 17332
rect 23716 17280 23722 17332
rect 23842 17280 23848 17332
rect 23900 17280 23906 17332
rect 26418 17280 26424 17332
rect 26476 17320 26482 17332
rect 27617 17323 27675 17329
rect 27617 17320 27629 17323
rect 26476 17292 27629 17320
rect 26476 17280 26482 17292
rect 27617 17289 27629 17292
rect 27663 17289 27675 17323
rect 27617 17283 27675 17289
rect 20898 17252 20904 17264
rect 13464 17224 14228 17252
rect 15672 17224 16896 17252
rect 16960 17224 17724 17252
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 12406 17156 13553 17184
rect 12069 17147 12127 17153
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 14200 17193 14228 17224
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 9723 17088 10333 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10652 17088 10701 17116
rect 10652 17076 10658 17088
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17116 11391 17119
rect 11790 17116 11796 17128
rect 11379 17088 11796 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 11790 17076 11796 17088
rect 11848 17116 11854 17128
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 11848 17088 11897 17116
rect 11848 17076 11854 17088
rect 11885 17085 11897 17088
rect 11931 17085 11943 17119
rect 11885 17079 11943 17085
rect 12618 17076 12624 17128
rect 12676 17076 12682 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 13648 17116 13676 17144
rect 15028 17116 15056 17147
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 16301 17187 16359 17193
rect 15528 17156 16252 17184
rect 15528 17144 15534 17156
rect 13648 17088 15056 17116
rect 12805 17079 12863 17085
rect 12820 17048 12848 17079
rect 15562 17076 15568 17128
rect 15620 17076 15626 17128
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 15712 17088 15761 17116
rect 15712 17076 15718 17088
rect 15749 17085 15761 17088
rect 15795 17085 15807 17119
rect 16224 17116 16252 17156
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16482 17184 16488 17196
rect 16347 17156 16488 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 16868 17193 16896 17224
rect 17696 17193 17724 17224
rect 19168 17224 20904 17252
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17175 17156 17233 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 17144 17116 17172 17147
rect 17770 17144 17776 17196
rect 17828 17144 17834 17196
rect 19168 17193 19196 17224
rect 20898 17212 20904 17224
rect 20956 17212 20962 17264
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 16224 17088 17172 17116
rect 15749 17079 15807 17085
rect 13357 17051 13415 17057
rect 13357 17048 13369 17051
rect 9600 17020 12434 17048
rect 12820 17020 13369 17048
rect 9171 17017 9183 17020
rect 9125 17011 9183 17017
rect 8202 16980 8208 16992
rect 7668 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 10594 16980 10600 16992
rect 8444 16952 10600 16980
rect 8444 16940 8450 16952
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 12406 16980 12434 17020
rect 13357 17017 13369 17020
rect 13403 17017 13415 17051
rect 19168 17048 19196 17147
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 19889 17187 19947 17193
rect 19889 17184 19901 17187
rect 19300 17156 19901 17184
rect 19300 17144 19306 17156
rect 19889 17153 19901 17156
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 13357 17011 13415 17017
rect 14752 17020 19196 17048
rect 20272 17048 20300 17147
rect 20438 17144 20444 17196
rect 20496 17144 20502 17196
rect 21358 17144 21364 17196
rect 21416 17184 21422 17196
rect 21637 17187 21695 17193
rect 21637 17184 21649 17187
rect 21416 17156 21649 17184
rect 21416 17144 21422 17156
rect 21637 17153 21649 17156
rect 21683 17153 21695 17187
rect 21637 17147 21695 17153
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 23290 17184 23296 17196
rect 22612 17156 23296 17184
rect 22612 17144 22618 17156
rect 23290 17144 23296 17156
rect 23348 17144 23354 17196
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17184 23443 17187
rect 23676 17184 23704 17280
rect 25308 17255 25366 17261
rect 25308 17221 25320 17255
rect 25354 17252 25366 17255
rect 26878 17252 26884 17264
rect 25354 17224 26884 17252
rect 25354 17221 25366 17224
rect 25308 17215 25366 17221
rect 26878 17212 26884 17224
rect 26936 17212 26942 17264
rect 23431 17156 23704 17184
rect 23431 17153 23443 17156
rect 23385 17147 23443 17153
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17184 25099 17187
rect 25130 17184 25136 17196
rect 25087 17156 25136 17184
rect 25087 17153 25099 17156
rect 25041 17147 25099 17153
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 26050 17144 26056 17196
rect 26108 17184 26114 17196
rect 26697 17187 26755 17193
rect 26697 17184 26709 17187
rect 26108 17156 26709 17184
rect 26108 17144 26114 17156
rect 26697 17153 26709 17156
rect 26743 17153 26755 17187
rect 26697 17147 26755 17153
rect 26970 17144 26976 17196
rect 27028 17144 27034 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27522 17184 27528 17196
rect 27203 17156 27528 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 20714 17116 20720 17128
rect 20671 17088 20720 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 20901 17119 20959 17125
rect 20901 17085 20913 17119
rect 20947 17085 20959 17119
rect 20901 17079 20959 17085
rect 23201 17119 23259 17125
rect 23201 17085 23213 17119
rect 23247 17116 23259 17119
rect 23474 17116 23480 17128
rect 23247 17088 23480 17116
rect 23247 17085 23259 17088
rect 23201 17079 23259 17085
rect 20806 17048 20812 17060
rect 20272 17020 20812 17048
rect 14752 16980 14780 17020
rect 20806 17008 20812 17020
rect 20864 17008 20870 17060
rect 20916 17048 20944 17079
rect 23474 17076 23480 17088
rect 23532 17116 23538 17128
rect 23768 17116 23796 17144
rect 23532 17088 23796 17116
rect 24213 17119 24271 17125
rect 23532 17076 23538 17088
rect 24213 17085 24225 17119
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 21453 17051 21511 17057
rect 21453 17048 21465 17051
rect 20916 17020 21465 17048
rect 21453 17017 21465 17020
rect 21499 17017 21511 17051
rect 24228 17048 24256 17079
rect 27632 17048 27660 17283
rect 28350 17280 28356 17332
rect 28408 17280 28414 17332
rect 27893 17187 27951 17193
rect 27893 17153 27905 17187
rect 27939 17184 27951 17187
rect 28368 17184 28396 17280
rect 27939 17156 28396 17184
rect 27939 17153 27951 17156
rect 27893 17147 27951 17153
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17116 27767 17119
rect 28074 17116 28080 17128
rect 27755 17088 28080 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 28074 17076 28080 17088
rect 28132 17076 28138 17128
rect 28169 17051 28227 17057
rect 28169 17048 28181 17051
rect 24228 17020 25084 17048
rect 21453 17011 21511 17017
rect 12406 16952 14780 16980
rect 14829 16983 14887 16989
rect 14829 16949 14841 16983
rect 14875 16980 14887 16983
rect 15194 16980 15200 16992
rect 14875 16952 15200 16980
rect 14875 16949 14887 16952
rect 14829 16943 14887 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16206 16940 16212 16992
rect 16264 16940 16270 16992
rect 16390 16940 16396 16992
rect 16448 16940 16454 16992
rect 17310 16940 17316 16992
rect 17368 16940 17374 16992
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 19337 16983 19395 16989
rect 19337 16949 19349 16983
rect 19383 16980 19395 16983
rect 19518 16980 19524 16992
rect 19383 16952 19524 16980
rect 19383 16949 19395 16952
rect 19337 16943 19395 16949
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 19702 16940 19708 16992
rect 19760 16940 19766 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20956 16952 21097 16980
rect 20956 16940 20962 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 24765 16983 24823 16989
rect 24765 16980 24777 16983
rect 23440 16952 24777 16980
rect 23440 16940 23446 16952
rect 24765 16949 24777 16952
rect 24811 16949 24823 16983
rect 25056 16980 25084 17020
rect 26436 17020 27568 17048
rect 27632 17020 28181 17048
rect 26436 16989 26464 17020
rect 26421 16983 26479 16989
rect 26421 16980 26433 16983
rect 25056 16952 26433 16980
rect 24765 16943 24823 16949
rect 26421 16949 26433 16952
rect 26467 16949 26479 16983
rect 26421 16943 26479 16949
rect 26510 16940 26516 16992
rect 26568 16940 26574 16992
rect 27540 16980 27568 17020
rect 28169 17017 28181 17020
rect 28215 17017 28227 17051
rect 28169 17011 28227 17017
rect 27614 16980 27620 16992
rect 27540 16952 27620 16980
rect 27614 16940 27620 16952
rect 27672 16940 27678 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2924 16748 3065 16776
rect 2924 16736 2930 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 3053 16739 3111 16745
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1452 16612 1685 16640
rect 1452 16600 1458 16612
rect 1673 16609 1685 16612
rect 1719 16609 1731 16643
rect 1673 16603 1731 16609
rect 3068 16572 3096 16739
rect 3234 16736 3240 16788
rect 3292 16736 3298 16788
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4396 16748 4629 16776
rect 4396 16736 4402 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 4617 16739 4675 16745
rect 7098 16736 7104 16788
rect 7156 16736 7162 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 7616 16748 7972 16776
rect 7616 16736 7622 16748
rect 6822 16708 6828 16720
rect 5736 16680 6828 16708
rect 5736 16649 5764 16680
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3344 16612 3801 16640
rect 3344 16584 3372 16612
rect 3789 16609 3801 16612
rect 3835 16640 3847 16643
rect 5721 16643 5779 16649
rect 3835 16612 4568 16640
rect 3835 16609 3847 16612
rect 3789 16603 3847 16609
rect 3145 16575 3203 16581
rect 3145 16572 3157 16575
rect 3068 16544 3157 16572
rect 3145 16541 3157 16544
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 3326 16532 3332 16584
rect 3384 16532 3390 16584
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 4540 16581 4568 16612
rect 5721 16609 5733 16643
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6549 16643 6607 16649
rect 6549 16640 6561 16643
rect 5951 16612 6561 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6549 16609 6561 16612
rect 6595 16609 6607 16643
rect 7116 16640 7144 16736
rect 7469 16643 7527 16649
rect 7469 16640 7481 16643
rect 7116 16612 7481 16640
rect 6549 16603 6607 16609
rect 7469 16609 7481 16612
rect 7515 16609 7527 16643
rect 7944 16640 7972 16748
rect 8938 16736 8944 16788
rect 8996 16776 9002 16788
rect 9033 16779 9091 16785
rect 9033 16776 9045 16779
rect 8996 16748 9045 16776
rect 8996 16736 9002 16748
rect 9033 16745 9045 16748
rect 9079 16745 9091 16779
rect 9033 16739 9091 16745
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9732 16748 9812 16776
rect 9732 16736 9738 16748
rect 8205 16643 8263 16649
rect 8205 16640 8217 16643
rect 7944 16612 8217 16640
rect 7469 16603 7527 16609
rect 8205 16609 8217 16612
rect 8251 16609 8263 16643
rect 8386 16640 8392 16652
rect 8205 16603 8263 16609
rect 8312 16612 8392 16640
rect 3605 16575 3663 16581
rect 3605 16572 3617 16575
rect 3568 16544 3617 16572
rect 3568 16532 3574 16544
rect 3605 16541 3617 16544
rect 3651 16541 3663 16575
rect 3605 16535 3663 16541
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16541 4583 16575
rect 4525 16535 4583 16541
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16541 7343 16575
rect 7285 16535 7343 16541
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16572 8079 16575
rect 8312 16572 8340 16612
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 8478 16600 8484 16652
rect 8536 16600 8542 16652
rect 9784 16640 9812 16748
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 9916 16748 10057 16776
rect 9916 16736 9922 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10045 16739 10103 16745
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10928 16748 10977 16776
rect 10928 16736 10934 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 11940 16748 12725 16776
rect 11940 16736 11946 16748
rect 12713 16745 12725 16748
rect 12759 16745 12771 16779
rect 12713 16739 12771 16745
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 14516 16748 15424 16776
rect 14516 16736 14522 16748
rect 11054 16708 11060 16720
rect 9959 16680 11060 16708
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9784 16612 9873 16640
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 8067 16544 8340 16572
rect 8496 16572 8524 16600
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8496 16544 8953 16572
rect 8067 16541 8079 16544
rect 8021 16535 8079 16541
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 1940 16507 1998 16513
rect 1940 16473 1952 16507
rect 1986 16504 1998 16507
rect 4433 16507 4491 16513
rect 4433 16504 4445 16507
rect 1986 16476 4445 16504
rect 1986 16473 1998 16476
rect 1940 16467 1998 16473
rect 4433 16473 4445 16476
rect 4479 16473 4491 16507
rect 4433 16467 4491 16473
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 6932 16504 6960 16532
rect 6411 16476 6960 16504
rect 7300 16504 7328 16535
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 9959 16504 9987 16680
rect 11054 16668 11060 16680
rect 11112 16708 11118 16720
rect 11112 16680 11192 16708
rect 11112 16668 11118 16680
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10778 16640 10784 16652
rect 10100 16612 10784 16640
rect 10100 16600 10106 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 11164 16649 11192 16680
rect 11149 16643 11207 16649
rect 11149 16609 11161 16643
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 12768 16612 14105 16640
rect 12768 16600 12774 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 15396 16640 15424 16748
rect 15470 16736 15476 16788
rect 15528 16736 15534 16788
rect 16206 16736 16212 16788
rect 16264 16736 16270 16788
rect 16390 16736 16396 16788
rect 16448 16736 16454 16788
rect 17218 16736 17224 16788
rect 17276 16736 17282 16788
rect 17310 16736 17316 16788
rect 17368 16736 17374 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 19610 16776 19616 16788
rect 17644 16748 19616 16776
rect 17644 16736 17650 16748
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 19702 16736 19708 16788
rect 19760 16736 19766 16788
rect 22186 16776 22192 16788
rect 20824 16748 22192 16776
rect 15746 16640 15752 16652
rect 15396 16612 15752 16640
rect 14093 16603 14151 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16408 16640 16436 16736
rect 15979 16612 16436 16640
rect 16853 16643 16911 16649
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 17328 16640 17356 16736
rect 17604 16649 17632 16736
rect 16899 16612 17356 16640
rect 17589 16643 17647 16649
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 19720 16640 19748 16736
rect 19567 16612 19748 16640
rect 20073 16643 20131 16649
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20622 16640 20628 16652
rect 20119 16612 20628 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16541 10931 16575
rect 10873 16535 10931 16541
rect 7300 16476 9987 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 10888 16504 10916 16535
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 11296 16544 11345 16572
rect 11296 16532 11302 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16572 13323 16575
rect 13630 16572 13636 16584
rect 13311 16544 13636 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 13722 16532 13728 16584
rect 13780 16532 13786 16584
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14349 16575 14407 16581
rect 14349 16572 14361 16575
rect 14240 16544 14361 16572
rect 14240 16532 14246 16544
rect 14349 16541 14361 16544
rect 14395 16541 14407 16575
rect 14349 16535 14407 16541
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 19334 16532 19340 16584
rect 19392 16532 19398 16584
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 20088 16572 20116 16603
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 20824 16649 20852 16748
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 26234 16736 26240 16788
rect 26292 16776 26298 16788
rect 27065 16779 27123 16785
rect 27065 16776 27077 16779
rect 26292 16748 27077 16776
rect 26292 16736 26298 16748
rect 27065 16745 27077 16748
rect 27111 16745 27123 16779
rect 27065 16739 27123 16745
rect 27709 16779 27767 16785
rect 27709 16745 27721 16779
rect 27755 16776 27767 16779
rect 27798 16776 27804 16788
rect 27755 16748 27804 16776
rect 27755 16745 27767 16748
rect 27709 16739 27767 16745
rect 27798 16736 27804 16748
rect 27856 16736 27862 16788
rect 23661 16711 23719 16717
rect 23661 16708 23673 16711
rect 23584 16680 23673 16708
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 21450 16600 21456 16652
rect 21508 16640 21514 16652
rect 21508 16612 21956 16640
rect 21508 16600 21514 16612
rect 19484 16544 20116 16572
rect 19484 16532 19490 16544
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20588 16544 21005 16572
rect 20588 16532 20594 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21542 16532 21548 16584
rect 21600 16532 21606 16584
rect 21928 16581 21956 16612
rect 23584 16597 23612 16680
rect 23661 16677 23673 16680
rect 23707 16677 23719 16711
rect 23661 16671 23719 16677
rect 26326 16668 26332 16720
rect 26384 16668 26390 16720
rect 25041 16643 25099 16649
rect 25041 16609 25053 16643
rect 25087 16640 25099 16643
rect 26344 16640 26372 16668
rect 25087 16612 26372 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 27985 16643 28043 16649
rect 27985 16609 27997 16643
rect 28031 16640 28043 16643
rect 28626 16640 28632 16652
rect 28031 16612 28632 16640
rect 28031 16609 28043 16612
rect 27985 16603 28043 16609
rect 28626 16600 28632 16612
rect 28684 16600 28690 16652
rect 23569 16591 23627 16597
rect 21913 16575 21971 16581
rect 21913 16541 21925 16575
rect 21959 16572 21971 16575
rect 22180 16575 22238 16581
rect 21959 16544 22140 16572
rect 21959 16541 21971 16544
rect 21913 16535 21971 16541
rect 11146 16504 11152 16516
rect 10100 16476 11152 16504
rect 10100 16464 10106 16476
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 11422 16464 11428 16516
rect 11480 16504 11486 16516
rect 11882 16504 11888 16516
rect 11480 16476 11888 16504
rect 11480 16464 11486 16476
rect 11882 16464 11888 16476
rect 11940 16504 11946 16516
rect 13740 16504 13768 16532
rect 15286 16504 15292 16516
rect 11940 16476 12434 16504
rect 13740 16476 15292 16504
rect 11940 16464 11946 16476
rect 3418 16396 3424 16448
rect 3476 16396 3482 16448
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 7929 16439 7987 16445
rect 7929 16436 7941 16439
rect 7800 16408 7941 16436
rect 7800 16396 7806 16408
rect 7929 16405 7941 16408
rect 7975 16436 7987 16439
rect 8665 16439 8723 16445
rect 8665 16436 8677 16439
rect 7975 16408 8677 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8665 16405 8677 16408
rect 8711 16405 8723 16439
rect 8665 16399 8723 16405
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 11698 16436 11704 16448
rect 9824 16408 11704 16436
rect 9824 16396 9830 16408
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 12406 16436 12434 16476
rect 15286 16464 15292 16476
rect 15344 16504 15350 16516
rect 16482 16504 16488 16516
rect 15344 16476 16488 16504
rect 15344 16464 15350 16476
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 17856 16507 17914 16513
rect 17856 16473 17868 16507
rect 17902 16504 17914 16507
rect 22112 16504 22140 16544
rect 22180 16541 22192 16575
rect 22226 16572 22238 16575
rect 23382 16572 23388 16584
rect 22226 16544 23388 16572
rect 22226 16541 22238 16544
rect 22180 16535 22238 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23569 16557 23581 16591
rect 23615 16557 23627 16591
rect 23569 16551 23627 16557
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16541 23903 16575
rect 23845 16535 23903 16541
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16572 24823 16575
rect 26973 16575 27031 16581
rect 24811 16544 24992 16572
rect 24811 16541 24823 16544
rect 24765 16535 24823 16541
rect 22370 16504 22376 16516
rect 17902 16476 22048 16504
rect 22112 16476 22376 16504
rect 17902 16473 17914 16476
rect 17856 16467 17914 16473
rect 14734 16436 14740 16448
rect 12406 16408 14740 16436
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 18966 16396 18972 16448
rect 19024 16396 19030 16448
rect 19981 16439 20039 16445
rect 19981 16405 19993 16439
rect 20027 16436 20039 16439
rect 20346 16436 20352 16448
rect 20027 16408 20352 16436
rect 20027 16405 20039 16408
rect 19981 16399 20039 16405
rect 20346 16396 20352 16408
rect 20404 16436 20410 16448
rect 20717 16439 20775 16445
rect 20717 16436 20729 16439
rect 20404 16408 20729 16436
rect 20404 16396 20410 16408
rect 20717 16405 20729 16408
rect 20763 16405 20775 16439
rect 20717 16399 20775 16405
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 20956 16408 21465 16436
rect 20956 16396 20962 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21453 16399 21511 16405
rect 21634 16396 21640 16448
rect 21692 16396 21698 16448
rect 22020 16436 22048 16476
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 23860 16504 23888 16535
rect 23308 16476 23888 16504
rect 22278 16436 22284 16448
rect 22020 16408 22284 16436
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 23014 16396 23020 16448
rect 23072 16436 23078 16448
rect 23308 16445 23336 16476
rect 24964 16448 24992 16544
rect 26973 16541 26985 16575
rect 27019 16572 27031 16575
rect 27172 16572 27200 16600
rect 27019 16544 27200 16572
rect 27019 16541 27031 16544
rect 26973 16535 27031 16541
rect 25225 16507 25283 16513
rect 25225 16473 25237 16507
rect 25271 16473 25283 16507
rect 25225 16467 25283 16473
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 23072 16408 23305 16436
rect 23072 16396 23078 16408
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 23382 16396 23388 16448
rect 23440 16396 23446 16448
rect 24578 16396 24584 16448
rect 24636 16396 24642 16448
rect 24946 16396 24952 16448
rect 25004 16396 25010 16448
rect 25240 16436 25268 16467
rect 26878 16464 26884 16516
rect 26936 16464 26942 16516
rect 27433 16507 27491 16513
rect 27433 16473 27445 16507
rect 27479 16504 27491 16507
rect 28350 16504 28356 16516
rect 27479 16476 28356 16504
rect 27479 16473 27491 16476
rect 27433 16467 27491 16473
rect 28350 16464 28356 16476
rect 28408 16464 28414 16516
rect 27798 16436 27804 16448
rect 25240 16408 27804 16436
rect 27798 16396 27804 16408
rect 27856 16396 27862 16448
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 28316 16408 28549 16436
rect 28316 16396 28322 16408
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 2777 16235 2835 16241
rect 2777 16201 2789 16235
rect 2823 16232 2835 16235
rect 3326 16232 3332 16244
rect 2823 16204 3332 16232
rect 2823 16201 2835 16204
rect 2777 16195 2835 16201
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3418 16192 3424 16244
rect 3476 16192 3482 16244
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16201 4031 16235
rect 3973 16195 4031 16201
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 1664 16099 1722 16105
rect 1664 16065 1676 16099
rect 1710 16096 1722 16099
rect 2222 16096 2228 16108
rect 1710 16068 2228 16096
rect 1710 16065 1722 16068
rect 1664 16059 1722 16065
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 3436 16096 3464 16192
rect 3513 16167 3571 16173
rect 3513 16133 3525 16167
rect 3559 16164 3571 16167
rect 3694 16164 3700 16176
rect 3559 16136 3700 16164
rect 3559 16133 3571 16136
rect 3513 16127 3571 16133
rect 3694 16124 3700 16136
rect 3752 16124 3758 16176
rect 3988 16164 4016 16195
rect 7742 16192 7748 16244
rect 7800 16192 7806 16244
rect 8478 16192 8484 16244
rect 8536 16192 8542 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9732 16204 9873 16232
rect 9732 16192 9738 16204
rect 9861 16201 9873 16204
rect 9907 16232 9919 16235
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 9907 16204 10609 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 12805 16235 12863 16241
rect 12805 16232 12817 16235
rect 12676 16204 12817 16232
rect 12676 16192 12682 16204
rect 12805 16201 12817 16204
rect 12851 16232 12863 16235
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 12851 16204 13553 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 13541 16195 13599 16201
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 14645 16235 14703 16241
rect 14645 16201 14657 16235
rect 14691 16201 14703 16235
rect 14645 16195 14703 16201
rect 7098 16164 7104 16176
rect 3988 16136 4568 16164
rect 4540 16105 4568 16136
rect 4632 16136 7104 16164
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3436 16068 3893 16096
rect 2961 16059 3019 16065
rect 3881 16065 3893 16068
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16096 4215 16099
rect 4525 16099 4583 16105
rect 4203 16068 4292 16096
rect 4203 16065 4215 16068
rect 4157 16059 4215 16065
rect 2976 16028 3004 16059
rect 3418 16028 3424 16040
rect 2976 16000 3424 16028
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3697 15963 3755 15969
rect 3697 15929 3709 15963
rect 3743 15960 3755 15963
rect 4154 15960 4160 15972
rect 3743 15932 4160 15960
rect 3743 15929 3755 15932
rect 3697 15923 3755 15929
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 4264 15892 4292 16068
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 4632 16037 4660 16136
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16096 6423 16099
rect 6914 16096 6920 16108
rect 6411 16068 6920 16096
rect 6411 16065 6423 16068
rect 6365 16059 6423 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 7760 16096 7788 16192
rect 8496 16164 8524 16192
rect 10042 16164 10048 16176
rect 8496 16136 10048 16164
rect 7607 16068 7788 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 8956 16105 8984 16136
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 14108 16164 14136 16195
rect 14660 16164 14688 16195
rect 15194 16192 15200 16244
rect 15252 16192 15258 16244
rect 15286 16192 15292 16244
rect 15344 16192 15350 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17276 16204 17417 16232
rect 17276 16192 17282 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 19061 16235 19119 16241
rect 19061 16201 19073 16235
rect 19107 16232 19119 16235
rect 19242 16232 19248 16244
rect 19107 16204 19248 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19521 16235 19579 16241
rect 19521 16201 19533 16235
rect 19567 16232 19579 16235
rect 20254 16232 20260 16244
rect 19567 16204 20260 16232
rect 19567 16201 19579 16204
rect 19521 16195 19579 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 20346 16192 20352 16244
rect 20404 16192 20410 16244
rect 20530 16232 20536 16244
rect 20456 16204 20536 16232
rect 11348 16136 11928 16164
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9079 16068 9413 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9824 16068 9965 16096
rect 9824 16056 9830 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 10060 16096 10088 16124
rect 11348 16105 11376 16136
rect 11900 16105 11928 16136
rect 12176 16136 13584 16164
rect 14108 16136 14412 16164
rect 14660 16136 15148 16164
rect 12176 16105 12204 16136
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10060 16068 11069 16096
rect 9953 16059 10011 16065
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11103 16068 11345 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11333 16065 11345 16068
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 12986 16096 12992 16108
rect 12943 16068 12992 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 4341 15963 4399 15969
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 4816 15960 4844 15991
rect 6546 15988 6552 16040
rect 6604 15988 6610 16040
rect 7742 15988 7748 16040
rect 7800 15988 7806 16040
rect 4387 15932 4844 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 4798 15892 4804 15904
rect 4264 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5166 15852 5172 15904
rect 5224 15852 5230 15904
rect 6730 15852 6736 15904
rect 6788 15852 6794 15904
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 7929 15895 7987 15901
rect 7929 15892 7941 15895
rect 7708 15864 7941 15892
rect 7708 15852 7714 15864
rect 7929 15861 7941 15864
rect 7975 15861 7987 15895
rect 7929 15855 7987 15861
rect 8662 15852 8668 15904
rect 8720 15852 8726 15904
rect 8864 15892 8892 16056
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 10134 15988 10140 16040
rect 10192 15988 10198 16040
rect 11808 16028 11836 16059
rect 12986 16056 12992 16068
rect 13044 16096 13050 16108
rect 13262 16096 13268 16108
rect 13044 16068 13268 16096
rect 13044 16056 13050 16068
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 12345 16031 12403 16037
rect 12345 16028 12357 16031
rect 11164 16000 11836 16028
rect 11992 16000 12357 16028
rect 9232 15960 9260 15988
rect 11164 15969 11192 16000
rect 11992 15969 12020 16000
rect 12345 15997 12357 16000
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 11149 15963 11207 15969
rect 9232 15932 11100 15960
rect 9582 15892 9588 15904
rect 8864 15864 9588 15892
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 10870 15852 10876 15904
rect 10928 15852 10934 15904
rect 11072 15892 11100 15932
rect 11149 15929 11161 15963
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 11977 15963 12035 15969
rect 11977 15929 11989 15963
rect 12023 15929 12035 15963
rect 11977 15923 12035 15929
rect 11422 15892 11428 15904
rect 11072 15864 11428 15892
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11609 15895 11667 15901
rect 11609 15861 11621 15895
rect 11655 15892 11667 15895
rect 13096 15892 13124 15991
rect 13556 15960 13584 16136
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16096 13875 16099
rect 14090 16096 14096 16108
rect 13863 16068 14096 16096
rect 13863 16065 13875 16068
rect 13817 16059 13875 16065
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 14274 16056 14280 16108
rect 14332 16056 14338 16108
rect 14384 16096 14412 16136
rect 15120 16105 15148 16136
rect 14529 16099 14587 16105
rect 14529 16096 14541 16099
rect 14384 16068 14541 16096
rect 14529 16065 14541 16068
rect 14575 16065 14587 16099
rect 14529 16059 14587 16065
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16065 15163 16099
rect 15212 16096 15240 16192
rect 15304 16164 15332 16192
rect 15304 16136 15516 16164
rect 15488 16105 15516 16136
rect 15381 16099 15439 16105
rect 15381 16096 15393 16099
rect 15212 16068 15393 16096
rect 15105 16059 15163 16065
rect 15381 16065 15393 16068
rect 15427 16065 15439 16099
rect 15381 16059 15439 16065
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16096 15623 16099
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15611 16068 15945 16096
rect 15611 16065 15623 16068
rect 15565 16059 15623 16065
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 14844 16028 14872 16059
rect 16206 16056 16212 16108
rect 16264 16096 16270 16108
rect 16761 16099 16819 16105
rect 16761 16096 16773 16099
rect 16264 16068 16773 16096
rect 16264 16056 16270 16068
rect 16761 16065 16773 16068
rect 16807 16065 16819 16099
rect 16761 16059 16819 16065
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17494 16096 17500 16108
rect 16991 16068 17500 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 18138 16096 18144 16108
rect 17727 16068 18144 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 18138 16056 18144 16068
rect 18196 16096 18202 16108
rect 20364 16105 20392 16192
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 18196 16068 19257 16096
rect 18196 16056 18202 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16096 19487 16099
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19475 16068 19993 16096
rect 19475 16065 19487 16068
rect 19429 16059 19487 16065
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 13688 16000 14872 16028
rect 13688 15988 13694 16000
rect 15654 15988 15660 16040
rect 15712 15988 15718 16040
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 16028 18291 16031
rect 19150 16028 19156 16040
rect 18279 16000 19156 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 14550 15960 14556 15972
rect 13556 15932 14556 15960
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 15197 15963 15255 15969
rect 14844 15932 15148 15960
rect 11655 15864 13124 15892
rect 13909 15895 13967 15901
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 14182 15892 14188 15904
rect 13955 15864 14188 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 14182 15852 14188 15864
rect 14240 15852 14246 15904
rect 14369 15895 14427 15901
rect 14369 15861 14381 15895
rect 14415 15892 14427 15895
rect 14844 15892 14872 15932
rect 14415 15864 14872 15892
rect 14415 15861 14427 15864
rect 14369 15855 14427 15861
rect 14918 15852 14924 15904
rect 14976 15852 14982 15904
rect 15120 15892 15148 15932
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 15672 15960 15700 15988
rect 15243 15932 15700 15960
rect 15764 15960 15792 15991
rect 19150 15988 19156 16000
rect 19208 16028 19214 16040
rect 19444 16028 19472 16059
rect 19208 16000 19472 16028
rect 19208 15988 19214 16000
rect 19426 15960 19432 15972
rect 15764 15932 19432 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 19996 15960 20024 16059
rect 20073 16031 20131 16037
rect 20073 15997 20085 16031
rect 20119 16028 20131 16031
rect 20456 16028 20484 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20806 16192 20812 16244
rect 20864 16232 20870 16244
rect 21361 16235 21419 16241
rect 21361 16232 21373 16235
rect 20864 16204 21373 16232
rect 20864 16192 20870 16204
rect 21361 16201 21373 16204
rect 21407 16201 21419 16235
rect 21361 16195 21419 16201
rect 21634 16192 21640 16244
rect 21692 16192 21698 16244
rect 25038 16192 25044 16244
rect 25096 16192 25102 16244
rect 26237 16235 26295 16241
rect 26237 16201 26249 16235
rect 26283 16232 26295 16235
rect 26602 16232 26608 16244
rect 26283 16204 26608 16232
rect 26283 16201 26295 16204
rect 26237 16195 26295 16201
rect 26602 16192 26608 16204
rect 26660 16192 26666 16244
rect 26973 16235 27031 16241
rect 26973 16201 26985 16235
rect 27019 16232 27031 16235
rect 28534 16232 28540 16244
rect 27019 16204 28540 16232
rect 27019 16201 27031 16204
rect 26973 16195 27031 16201
rect 28534 16192 28540 16204
rect 28592 16192 28598 16244
rect 21652 16164 21680 16192
rect 20548 16136 21680 16164
rect 22557 16167 22615 16173
rect 20548 16105 20576 16136
rect 22557 16133 22569 16167
rect 22603 16164 22615 16167
rect 22646 16164 22652 16176
rect 22603 16136 22652 16164
rect 22603 16133 22615 16136
rect 22557 16127 22615 16133
rect 22646 16124 22652 16136
rect 22704 16164 22710 16176
rect 24946 16164 24952 16176
rect 22704 16136 24952 16164
rect 22704 16124 22710 16136
rect 24946 16124 24952 16136
rect 25004 16164 25010 16176
rect 25004 16136 26372 16164
rect 25004 16124 25010 16136
rect 26344 16108 26372 16136
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16065 20591 16099
rect 21077 16089 21135 16095
rect 21077 16086 21089 16089
rect 20533 16059 20591 16065
rect 21008 16058 21089 16086
rect 21008 16028 21036 16058
rect 21077 16055 21089 16058
rect 21123 16055 21135 16089
rect 21266 16056 21272 16108
rect 21324 16056 21330 16108
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21508 16068 21557 16096
rect 21508 16056 21514 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 21077 16049 21135 16055
rect 20119 16000 20484 16028
rect 20539 16000 21036 16028
rect 21284 16028 21312 16056
rect 21818 16028 21824 16040
rect 21284 16000 21824 16028
rect 20119 15997 20131 16000
rect 20073 15991 20131 15997
rect 20539 15960 20567 16000
rect 21818 15988 21824 16000
rect 21876 15988 21882 16040
rect 22020 16028 22048 16059
rect 23382 16056 23388 16108
rect 23440 16096 23446 16108
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23440 16068 23673 16096
rect 23440 16056 23446 16068
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 24486 16056 24492 16108
rect 24544 16096 24550 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24544 16068 24593 16096
rect 24544 16056 24550 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16096 25191 16099
rect 25682 16096 25688 16108
rect 25179 16068 25688 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22020 16000 22845 16028
rect 22833 15997 22845 16000
rect 22879 16028 22891 16031
rect 23014 16028 23020 16040
rect 22879 16000 23020 16028
rect 22879 15997 22891 16000
rect 22833 15991 22891 15997
rect 23014 15988 23020 16000
rect 23072 15988 23078 16040
rect 23474 15988 23480 16040
rect 23532 15988 23538 16040
rect 23566 15988 23572 16040
rect 23624 16028 23630 16040
rect 24397 16031 24455 16037
rect 24397 16028 24409 16031
rect 23624 16000 24409 16028
rect 23624 15988 23630 16000
rect 24397 15997 24409 16000
rect 24443 15997 24455 16031
rect 25148 16028 25176 16059
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 24397 15991 24455 15997
rect 24504 16000 25176 16028
rect 25317 16031 25375 16037
rect 19996 15932 20567 15960
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 20680 15932 20729 15960
rect 20680 15920 20686 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 20806 15920 20812 15972
rect 20864 15960 20870 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20864 15932 21189 15960
rect 20864 15920 20870 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 23492 15960 23520 15988
rect 24504 15960 24532 16000
rect 25317 15997 25329 16031
rect 25363 15997 25375 16031
rect 26068 16028 26096 16059
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 26605 16099 26663 16105
rect 26605 16096 26617 16099
rect 26384 16068 26617 16096
rect 26384 16056 26390 16068
rect 26605 16065 26617 16068
rect 26651 16096 26663 16099
rect 26970 16096 26976 16108
rect 26651 16068 26976 16096
rect 26651 16065 26663 16068
rect 26605 16059 26663 16065
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 27154 16056 27160 16108
rect 27212 16105 27218 16108
rect 27212 16096 27223 16105
rect 27212 16068 27257 16096
rect 27212 16059 27223 16068
rect 27212 16056 27218 16059
rect 27338 16056 27344 16108
rect 27396 16056 27402 16108
rect 27430 16056 27436 16108
rect 27488 16096 27494 16108
rect 27893 16099 27951 16105
rect 27893 16096 27905 16099
rect 27488 16068 27905 16096
rect 27488 16056 27494 16068
rect 27893 16065 27905 16068
rect 27939 16065 27951 16099
rect 27893 16059 27951 16065
rect 27062 16028 27068 16040
rect 26068 16000 27068 16028
rect 25317 15991 25375 15997
rect 21177 15923 21235 15929
rect 22066 15932 23520 15960
rect 23584 15932 24532 15960
rect 15286 15892 15292 15904
rect 15120 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 16393 15895 16451 15901
rect 16393 15861 16405 15895
rect 16439 15892 16451 15895
rect 16666 15892 16672 15904
rect 16439 15864 16672 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 16666 15852 16672 15864
rect 16724 15892 16730 15904
rect 17218 15892 17224 15904
rect 16724 15864 17224 15892
rect 16724 15852 16730 15864
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 22066 15892 22094 15932
rect 23584 15904 23612 15932
rect 24854 15920 24860 15972
rect 24912 15960 24918 15972
rect 25332 15960 25360 15991
rect 27062 15988 27068 16000
rect 27120 15988 27126 16040
rect 27706 16028 27712 16040
rect 27540 16000 27712 16028
rect 24912 15932 25360 15960
rect 24912 15920 24918 15932
rect 25958 15920 25964 15972
rect 26016 15960 26022 15972
rect 26697 15963 26755 15969
rect 26697 15960 26709 15963
rect 26016 15932 26709 15960
rect 26016 15920 26022 15932
rect 26697 15929 26709 15932
rect 26743 15929 26755 15963
rect 26697 15923 26755 15929
rect 19392 15864 22094 15892
rect 19392 15852 19398 15864
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 23566 15852 23572 15904
rect 23624 15852 23630 15904
rect 24026 15852 24032 15904
rect 24084 15852 24090 15904
rect 25774 15852 25780 15904
rect 25832 15852 25838 15904
rect 26418 15852 26424 15904
rect 26476 15852 26482 15904
rect 26786 15852 26792 15904
rect 26844 15892 26850 15904
rect 27540 15901 27568 16000
rect 27706 15988 27712 16000
rect 27764 15988 27770 16040
rect 27525 15895 27583 15901
rect 27525 15892 27537 15895
rect 26844 15864 27537 15892
rect 26844 15852 26850 15864
rect 27525 15861 27537 15864
rect 27571 15861 27583 15895
rect 27525 15855 27583 15861
rect 28074 15852 28080 15904
rect 28132 15852 28138 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 2222 15648 2228 15700
rect 2280 15648 2286 15700
rect 5166 15648 5172 15700
rect 5224 15648 5230 15700
rect 6641 15691 6699 15697
rect 6641 15657 6653 15691
rect 6687 15688 6699 15691
rect 6730 15688 6736 15700
rect 6687 15660 6736 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 7800 15660 8493 15688
rect 7800 15648 7806 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 8662 15648 8668 15700
rect 8720 15648 8726 15700
rect 9309 15691 9367 15697
rect 9309 15657 9321 15691
rect 9355 15688 9367 15691
rect 10134 15688 10140 15700
rect 9355 15660 10140 15688
rect 9355 15657 9367 15660
rect 9309 15651 9367 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10870 15648 10876 15700
rect 10928 15648 10934 15700
rect 12710 15688 12716 15700
rect 12544 15660 12716 15688
rect 3421 15623 3479 15629
rect 3421 15589 3433 15623
rect 3467 15620 3479 15623
rect 4154 15620 4160 15632
rect 3467 15592 4160 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 5184 15552 5212 15648
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 3752 15524 4016 15552
rect 5184 15524 5273 15552
rect 3752 15512 3758 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 2222 15484 2228 15496
rect 1719 15456 2228 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2314 15444 2320 15496
rect 2372 15444 2378 15496
rect 3326 15444 3332 15496
rect 3384 15444 3390 15496
rect 3988 15493 4016 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6362 15552 6368 15564
rect 6043 15524 6368 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 6748 15552 6776 15648
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6748 15524 6837 15552
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7515 15524 7941 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 7929 15521 7941 15524
rect 7975 15552 7987 15555
rect 8294 15552 8300 15564
rect 7975 15524 8300 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4433 15487 4491 15493
rect 4433 15453 4445 15487
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 3620 15416 3648 15447
rect 4448 15416 4476 15447
rect 4522 15444 4528 15496
rect 4580 15444 4586 15496
rect 4706 15444 4712 15496
rect 4764 15444 4770 15496
rect 5442 15444 5448 15496
rect 5500 15444 5506 15496
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 6178 15444 6184 15496
rect 6236 15444 6242 15496
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8478 15484 8484 15496
rect 8435 15456 8484 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 8680 15484 8708 15648
rect 10042 15512 10048 15564
rect 10100 15512 10106 15564
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 8680 15456 9505 15484
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9640 15456 9781 15484
rect 9640 15444 9646 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 10888 15484 10916 15648
rect 12544 15561 12572 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 14918 15648 14924 15700
rect 14976 15648 14982 15700
rect 17218 15648 17224 15700
rect 17276 15648 17282 15700
rect 20530 15688 20536 15700
rect 18156 15660 20536 15688
rect 13909 15623 13967 15629
rect 13909 15589 13921 15623
rect 13955 15589 13967 15623
rect 13909 15583 13967 15589
rect 12529 15555 12587 15561
rect 11072 15524 12204 15552
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10888 15456 10977 15484
rect 9769 15447 9827 15453
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 5920 15416 5948 15444
rect 3620 15388 4016 15416
rect 4448 15388 5948 15416
rect 3988 15360 4016 15388
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 7650 15376 7656 15428
rect 7708 15376 7714 15428
rect 7742 15376 7748 15428
rect 7800 15376 7806 15428
rect 9784 15416 9812 15447
rect 11072 15416 11100 15524
rect 12176 15496 12204 15524
rect 12529 15521 12541 15555
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 11238 15444 11244 15496
rect 11296 15444 11302 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 13924 15484 13952 15583
rect 14936 15552 14964 15648
rect 15010 15580 15016 15632
rect 15068 15620 15074 15632
rect 15068 15592 17908 15620
rect 15068 15580 15074 15592
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 14936 15524 17049 15552
rect 17037 15521 17049 15524
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 12216 15456 13952 15484
rect 12216 15444 12222 15456
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 9784 15388 11100 15416
rect 2958 15308 2964 15360
rect 3016 15308 3022 15360
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 3145 15351 3203 15357
rect 3145 15348 3157 15351
rect 3108 15320 3157 15348
rect 3108 15308 3114 15320
rect 3145 15317 3157 15320
rect 3191 15317 3203 15351
rect 3145 15311 3203 15317
rect 3970 15308 3976 15360
rect 4028 15308 4034 15360
rect 4062 15308 4068 15360
rect 4120 15308 4126 15360
rect 4246 15308 4252 15360
rect 4304 15308 4310 15360
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 7668 15348 7696 15376
rect 5951 15320 7696 15348
rect 10781 15351 10839 15357
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 10781 15317 10793 15351
rect 10827 15348 10839 15351
rect 11256 15348 11284 15444
rect 12796 15419 12854 15425
rect 12796 15385 12808 15419
rect 12842 15416 12854 15419
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 12842 15388 14749 15416
rect 12842 15385 12854 15388
rect 12796 15379 12854 15385
rect 14737 15385 14749 15388
rect 14783 15385 14795 15419
rect 14737 15379 14795 15385
rect 14826 15376 14832 15428
rect 14884 15416 14890 15428
rect 15013 15419 15071 15425
rect 15013 15416 15025 15419
rect 14884 15388 15025 15416
rect 14884 15376 14890 15388
rect 15013 15385 15025 15388
rect 15059 15385 15071 15419
rect 16868 15416 16896 15447
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17276 15456 17785 15484
rect 17276 15444 17282 15456
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17880 15484 17908 15592
rect 18156 15561 18184 15660
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 21266 15688 21272 15700
rect 20916 15660 21272 15688
rect 18248 15592 20208 15620
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15521 18199 15555
rect 18141 15515 18199 15521
rect 18248 15484 18276 15592
rect 18325 15555 18383 15561
rect 18325 15521 18337 15555
rect 18371 15552 18383 15555
rect 18969 15555 19027 15561
rect 18969 15552 18981 15555
rect 18371 15524 18981 15552
rect 18371 15521 18383 15524
rect 18325 15515 18383 15521
rect 18969 15521 18981 15524
rect 19015 15521 19027 15555
rect 18969 15515 19027 15521
rect 19150 15512 19156 15564
rect 19208 15512 19214 15564
rect 19242 15512 19248 15564
rect 19300 15552 19306 15564
rect 20180 15561 20208 15592
rect 20622 15580 20628 15632
rect 20680 15620 20686 15632
rect 20916 15620 20944 15660
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 22278 15648 22284 15700
rect 22336 15648 22342 15700
rect 24026 15648 24032 15700
rect 24084 15648 24090 15700
rect 24854 15648 24860 15700
rect 24912 15648 24918 15700
rect 25774 15648 25780 15700
rect 25832 15648 25838 15700
rect 25958 15648 25964 15700
rect 26016 15648 26022 15700
rect 26418 15648 26424 15700
rect 26476 15648 26482 15700
rect 26881 15691 26939 15697
rect 26881 15657 26893 15691
rect 26927 15688 26939 15691
rect 28074 15688 28080 15700
rect 26927 15660 28080 15688
rect 26927 15657 26939 15660
rect 26881 15651 26939 15657
rect 25590 15620 25596 15632
rect 20680 15592 20944 15620
rect 21468 15592 25596 15620
rect 20680 15580 20686 15592
rect 20165 15555 20223 15561
rect 19300 15524 20116 15552
rect 19300 15512 19306 15524
rect 17880 15456 18276 15484
rect 17773 15447 17831 15453
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19168 15484 19196 15512
rect 18932 15456 19196 15484
rect 19429 15487 19487 15493
rect 18932 15444 18938 15456
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 20088 15484 20116 15524
rect 20165 15521 20177 15555
rect 20211 15521 20223 15555
rect 20165 15515 20223 15521
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20806 15552 20812 15564
rect 20395 15524 20812 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 20898 15512 20904 15564
rect 20956 15512 20962 15564
rect 21082 15512 21088 15564
rect 21140 15512 21146 15564
rect 21468 15484 21496 15592
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 23385 15555 23443 15561
rect 23385 15552 23397 15555
rect 23256 15524 23397 15552
rect 23256 15512 23262 15524
rect 23385 15521 23397 15524
rect 23431 15521 23443 15555
rect 23385 15515 23443 15521
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 25148 15561 25176 15592
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 25133 15555 25191 15561
rect 25133 15521 25145 15555
rect 25179 15521 25191 15555
rect 25133 15515 25191 15521
rect 25317 15555 25375 15561
rect 25317 15521 25329 15555
rect 25363 15552 25375 15555
rect 25976 15552 26004 15648
rect 26326 15552 26332 15564
rect 25363 15524 26004 15552
rect 26068 15524 26332 15552
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 20088 15456 21496 15484
rect 19429 15447 19487 15453
rect 19334 15416 19340 15428
rect 16868 15388 19340 15416
rect 15013 15379 15071 15385
rect 19334 15376 19340 15388
rect 19392 15376 19398 15428
rect 19444 15416 19472 15447
rect 21634 15444 21640 15496
rect 21692 15444 21698 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22373 15487 22431 15493
rect 22373 15484 22385 15487
rect 22244 15456 22385 15484
rect 22244 15444 22250 15456
rect 22373 15453 22385 15456
rect 22419 15484 22431 15487
rect 22462 15484 22468 15496
rect 22419 15456 22468 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 22554 15444 22560 15496
rect 22612 15444 22618 15496
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23293 15487 23351 15493
rect 23293 15484 23305 15487
rect 23072 15456 23305 15484
rect 23072 15444 23078 15456
rect 23293 15453 23305 15456
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15453 23627 15487
rect 23569 15447 23627 15453
rect 21450 15416 21456 15428
rect 19444 15388 21456 15416
rect 10827 15320 11284 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12066 15348 12072 15360
rect 11756 15320 12072 15348
rect 11756 15308 11762 15320
rect 12066 15308 12072 15320
rect 12124 15348 12130 15360
rect 13998 15348 14004 15360
rect 12124 15320 14004 15348
rect 12124 15308 12130 15320
rect 13998 15308 14004 15320
rect 14056 15348 14062 15360
rect 16114 15348 16120 15360
rect 14056 15320 16120 15348
rect 14056 15308 14062 15320
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16298 15308 16304 15360
rect 16356 15308 16362 15360
rect 17586 15308 17592 15360
rect 17644 15308 17650 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 18564 15320 18797 15348
rect 18564 15308 18570 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 18966 15308 18972 15360
rect 19024 15348 19030 15360
rect 19444 15348 19472 15388
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 21818 15376 21824 15428
rect 21876 15416 21882 15428
rect 23198 15416 23204 15428
rect 21876 15388 23204 15416
rect 21876 15376 21882 15388
rect 23198 15376 23204 15388
rect 23256 15376 23262 15428
rect 23584 15416 23612 15447
rect 23934 15444 23940 15496
rect 23992 15484 23998 15496
rect 24489 15487 24547 15493
rect 24489 15484 24501 15487
rect 23992 15456 24501 15484
rect 23992 15444 23998 15456
rect 24489 15453 24501 15456
rect 24535 15453 24547 15487
rect 24596 15484 24624 15512
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 24596 15456 25053 15484
rect 24489 15447 24547 15453
rect 25041 15453 25053 15456
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 25869 15487 25927 15493
rect 25869 15453 25881 15487
rect 25915 15484 25927 15487
rect 26068 15484 26096 15524
rect 26326 15512 26332 15524
rect 26384 15512 26390 15564
rect 26436 15561 26464 15648
rect 26421 15555 26479 15561
rect 26421 15521 26433 15555
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 26694 15512 26700 15564
rect 26752 15512 26758 15564
rect 26988 15561 27016 15660
rect 28074 15648 28080 15660
rect 28132 15648 28138 15700
rect 28350 15648 28356 15700
rect 28408 15648 28414 15700
rect 27062 15580 27068 15632
rect 27120 15620 27126 15632
rect 27985 15623 28043 15629
rect 27985 15620 27997 15623
rect 27120 15592 27997 15620
rect 27120 15580 27126 15592
rect 27985 15589 27997 15592
rect 28031 15589 28043 15623
rect 27985 15583 28043 15589
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 27614 15512 27620 15564
rect 27672 15512 27678 15564
rect 27798 15512 27804 15564
rect 27856 15512 27862 15564
rect 26237 15487 26295 15493
rect 26237 15484 26249 15487
rect 25915 15456 26096 15484
rect 26160 15456 26249 15484
rect 25915 15453 25927 15456
rect 25869 15447 25927 15453
rect 25961 15419 26019 15425
rect 25961 15416 25973 15419
rect 23584 15388 25973 15416
rect 25961 15385 25973 15388
rect 26007 15385 26019 15419
rect 25961 15379 26019 15385
rect 19024 15320 19472 15348
rect 19024 15308 19030 15320
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 20073 15351 20131 15357
rect 20073 15348 20085 15351
rect 20036 15320 20085 15348
rect 20036 15308 20042 15320
rect 20073 15317 20085 15320
rect 20119 15317 20131 15351
rect 20073 15311 20131 15317
rect 20806 15308 20812 15360
rect 20864 15308 20870 15360
rect 22922 15308 22928 15360
rect 22980 15348 22986 15360
rect 23017 15351 23075 15357
rect 23017 15348 23029 15351
rect 22980 15320 23029 15348
rect 22980 15308 22986 15320
rect 23017 15317 23029 15320
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 23106 15308 23112 15360
rect 23164 15308 23170 15360
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 24581 15351 24639 15357
rect 24581 15348 24593 15351
rect 23532 15320 24593 15348
rect 23532 15308 23538 15320
rect 24581 15317 24593 15320
rect 24627 15317 24639 15351
rect 24581 15311 24639 15317
rect 24762 15308 24768 15360
rect 24820 15348 24826 15360
rect 26160 15348 26188 15456
rect 26237 15453 26249 15456
rect 26283 15484 26295 15487
rect 26712 15484 26740 15512
rect 26283 15456 26740 15484
rect 27157 15487 27215 15493
rect 26283 15453 26295 15456
rect 26237 15447 26295 15453
rect 27157 15453 27169 15487
rect 27203 15453 27215 15487
rect 27632 15484 27660 15512
rect 27709 15487 27767 15493
rect 27709 15484 27721 15487
rect 27632 15456 27721 15484
rect 27157 15447 27215 15453
rect 27709 15453 27721 15456
rect 27755 15484 27767 15487
rect 28169 15487 28227 15493
rect 28169 15484 28181 15487
rect 27755 15456 28181 15484
rect 27755 15453 27767 15456
rect 27709 15447 27767 15453
rect 28169 15453 28181 15456
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15484 28319 15487
rect 28307 15456 28488 15484
rect 28307 15453 28319 15456
rect 28261 15447 28319 15453
rect 27172 15416 27200 15447
rect 28350 15416 28356 15428
rect 27172 15388 28356 15416
rect 28350 15376 28356 15388
rect 28408 15376 28414 15428
rect 24820 15320 26188 15348
rect 24820 15308 24826 15320
rect 26234 15308 26240 15360
rect 26292 15348 26298 15360
rect 27338 15348 27344 15360
rect 26292 15320 27344 15348
rect 26292 15308 26298 15320
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27617 15351 27675 15357
rect 27617 15317 27629 15351
rect 27663 15348 27675 15351
rect 27706 15348 27712 15360
rect 27663 15320 27712 15348
rect 27663 15317 27675 15320
rect 27617 15311 27675 15317
rect 27706 15308 27712 15320
rect 27764 15308 27770 15360
rect 27798 15308 27804 15360
rect 27856 15348 27862 15360
rect 28166 15348 28172 15360
rect 27856 15320 28172 15348
rect 27856 15308 27862 15320
rect 28166 15308 28172 15320
rect 28224 15348 28230 15360
rect 28460 15348 28488 15456
rect 28224 15320 28488 15348
rect 28224 15308 28230 15320
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 2777 15147 2835 15153
rect 2777 15144 2789 15147
rect 2280 15116 2789 15144
rect 2280 15104 2286 15116
rect 2777 15113 2789 15116
rect 2823 15113 2835 15147
rect 2777 15107 2835 15113
rect 4246 15104 4252 15156
rect 4304 15104 4310 15156
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4764 15116 4813 15144
rect 4764 15104 4770 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 5261 15147 5319 15153
rect 5261 15113 5273 15147
rect 5307 15144 5319 15147
rect 5442 15144 5448 15156
rect 5307 15116 5448 15144
rect 5307 15113 5319 15116
rect 5261 15107 5319 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 6178 15144 6184 15156
rect 6043 15116 6184 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 6362 15104 6368 15156
rect 6420 15104 6426 15156
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 6604 15116 6745 15144
rect 6604 15104 6610 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15113 7067 15147
rect 7009 15107 7067 15113
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 7742 15144 7748 15156
rect 7515 15116 7748 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 1664 15079 1722 15085
rect 1664 15045 1676 15079
rect 1710 15076 1722 15079
rect 2958 15076 2964 15088
rect 1710 15048 2964 15076
rect 1710 15045 1722 15048
rect 1664 15039 1722 15045
rect 2958 15036 2964 15048
rect 3016 15036 3022 15088
rect 3970 15036 3976 15088
rect 4028 15076 4034 15088
rect 4264 15076 4292 15104
rect 7024 15076 7052 15107
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15113 10471 15147
rect 13906 15144 13912 15156
rect 10413 15107 10471 15113
rect 13004 15116 13912 15144
rect 10428 15076 10456 15107
rect 12710 15076 12716 15088
rect 4028 15048 4200 15076
rect 4264 15048 5488 15076
rect 4028 15036 4034 15048
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 4062 15008 4068 15020
rect 3099 14980 4068 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4172 15008 4200 15048
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4172 14980 4445 15008
rect 4433 14977 4445 14980
rect 4479 15008 4491 15011
rect 4709 15011 4767 15017
rect 4479 14980 4660 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 1394 14900 1400 14952
rect 1452 14900 1458 14952
rect 2866 14900 2872 14952
rect 2924 14900 2930 14952
rect 3697 14943 3755 14949
rect 3697 14940 3709 14943
rect 3252 14912 3709 14940
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3252 14813 3280 14912
rect 3697 14909 3709 14912
rect 3743 14909 3755 14943
rect 3697 14903 3755 14909
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4525 14943 4583 14949
rect 4525 14940 4537 14943
rect 3927 14912 4537 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4525 14909 4537 14912
rect 4571 14909 4583 14943
rect 4632 14940 4660 14980
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 4798 15008 4804 15020
rect 4755 14980 4804 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 5460 15017 5488 15048
rect 5920 15048 6684 15076
rect 7024 15048 7880 15076
rect 10428 15048 10916 15076
rect 5920 15020 5948 15048
rect 5445 15011 5503 15017
rect 5445 14977 5457 15011
rect 5491 14977 5503 15011
rect 5445 14971 5503 14977
rect 5902 14968 5908 15020
rect 5960 14968 5966 15020
rect 6656 15017 6684 15048
rect 7852 15017 7880 15048
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 6641 14971 6699 14977
rect 6748 14980 7205 15008
rect 6196 14940 6224 14971
rect 4632 14912 5028 14940
rect 4525 14903 4583 14909
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 3200 14776 3249 14804
rect 3200 14764 3206 14776
rect 3237 14773 3249 14776
rect 3283 14773 3295 14807
rect 3237 14767 3295 14773
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 4890 14804 4896 14816
rect 4396 14776 4896 14804
rect 4396 14764 4402 14776
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5000 14804 5028 14912
rect 5736 14912 6224 14940
rect 5736 14881 5764 14912
rect 5721 14875 5779 14881
rect 5721 14841 5733 14875
rect 5767 14841 5779 14875
rect 5721 14835 5779 14841
rect 6362 14804 6368 14816
rect 5000 14776 6368 14804
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6656 14804 6684 14971
rect 6748 14884 6776 14980
rect 7193 14977 7205 14980
rect 7239 15008 7251 15011
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7239 14980 7389 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8018 14968 8024 15020
rect 8076 14968 8082 15020
rect 8294 14968 8300 15020
rect 8352 14968 8358 15020
rect 10888 15017 10916 15048
rect 12084 15048 12716 15076
rect 12084 15017 12112 15048
rect 12710 15036 12716 15048
rect 12768 15036 12774 15088
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 9968 14980 10272 15008
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 6730 14832 6736 14884
rect 6788 14832 6794 14884
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 6972 14844 7665 14872
rect 6972 14832 6978 14844
rect 7653 14841 7665 14844
rect 7699 14841 7711 14875
rect 7653 14835 7711 14841
rect 8205 14875 8263 14881
rect 8205 14841 8217 14875
rect 8251 14872 8263 14875
rect 8496 14872 8524 14903
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 9968 14940 9996 14980
rect 9548 14912 9996 14940
rect 10045 14943 10103 14949
rect 9548 14900 9554 14912
rect 10045 14909 10057 14943
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 8251 14844 8524 14872
rect 8251 14841 8263 14844
rect 8205 14835 8263 14841
rect 10060 14816 10088 14903
rect 10244 14872 10272 14980
rect 10336 14980 10609 15008
rect 10336 14952 10364 14980
rect 10597 14977 10609 14980
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12336 15011 12394 15017
rect 12336 14977 12348 15011
rect 12382 15008 12394 15011
rect 13004 15008 13032 15116
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 15470 15144 15476 15156
rect 14608 15116 15476 15144
rect 14608 15104 14614 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15144 16727 15147
rect 17218 15144 17224 15156
rect 16715 15116 17224 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 18874 15144 18880 15156
rect 17328 15116 18880 15144
rect 14458 15076 14464 15088
rect 12382 14980 13032 15008
rect 13096 15048 14464 15076
rect 12382 14977 12394 14980
rect 12336 14971 12394 14977
rect 10318 14900 10324 14952
rect 10376 14900 10382 14952
rect 10244 14844 10824 14872
rect 8478 14804 8484 14816
rect 6656 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 10686 14764 10692 14816
rect 10744 14764 10750 14816
rect 10796 14804 10824 14844
rect 13096 14804 13124 15048
rect 14458 15036 14464 15048
rect 14516 15036 14522 15088
rect 17328 15076 17356 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20806 15144 20812 15156
rect 20579 15116 20812 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 16868 15048 17356 15076
rect 18156 15048 20208 15076
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15746 15008 15752 15020
rect 15436 14980 15752 15008
rect 15436 14968 15442 14980
rect 15746 14968 15752 14980
rect 15804 15008 15810 15020
rect 16868 15017 16896 15048
rect 16853 15011 16911 15017
rect 15804 14980 16068 15008
rect 15804 14968 15810 14980
rect 13998 14900 14004 14952
rect 14056 14900 14062 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 13909 14875 13967 14881
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 14200 14872 14228 14903
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 15470 14900 15476 14952
rect 15528 14900 15534 14952
rect 15930 14900 15936 14952
rect 15988 14900 15994 14952
rect 16040 14940 16068 14980
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 15008 17003 15011
rect 17497 15011 17555 15017
rect 16991 14980 17448 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 16040 14912 17325 14940
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 13955 14844 14228 14872
rect 15488 14872 15516 14900
rect 17126 14872 17132 14884
rect 15488 14844 17132 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 17420 14872 17448 14980
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 17586 15008 17592 15020
rect 17543 14980 17592 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 18156 15017 18184 15048
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 14977 19027 15011
rect 19794 15008 19800 15020
rect 18969 14971 19027 14977
rect 19076 14980 19800 15008
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18288 14912 18337 14940
rect 18288 14900 18294 14912
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 18325 14903 18383 14909
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 18984 14940 19012 14971
rect 18564 14912 19012 14940
rect 18564 14900 18570 14912
rect 19076 14872 19104 14980
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 20180 14952 20208 15048
rect 20640 15017 20668 15116
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 21358 15104 21364 15156
rect 21416 15104 21422 15156
rect 26697 15147 26755 15153
rect 22296 15116 26648 15144
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 21174 15076 21180 15088
rect 20772 15048 21180 15076
rect 20772 15036 20778 15048
rect 21174 15036 21180 15048
rect 21232 15076 21238 15088
rect 21232 15048 21864 15076
rect 21232 15036 21238 15048
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 14977 20683 15011
rect 21082 15008 21088 15020
rect 20625 14971 20683 14977
rect 20732 14980 21088 15008
rect 19150 14900 19156 14952
rect 19208 14900 19214 14952
rect 19242 14900 19248 14952
rect 19300 14900 19306 14952
rect 19886 14900 19892 14952
rect 19944 14900 19950 14952
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20162 14900 20168 14952
rect 20220 14940 20226 14952
rect 20732 14940 20760 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21836 15017 21864 15048
rect 21545 15011 21603 15017
rect 21545 14977 21557 15011
rect 21591 14977 21603 15011
rect 21545 14971 21603 14977
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 14977 21879 15011
rect 22296 15008 22324 15116
rect 22370 15036 22376 15088
rect 22428 15076 22434 15088
rect 25130 15076 25136 15088
rect 22428 15048 25136 15076
rect 22428 15036 22434 15048
rect 22572 15017 22600 15048
rect 25130 15036 25136 15048
rect 25188 15036 25194 15088
rect 26620 15020 26648 15116
rect 26697 15113 26709 15147
rect 26743 15144 26755 15147
rect 27706 15144 27712 15156
rect 26743 15116 27712 15144
rect 26743 15113 26755 15116
rect 26697 15107 26755 15113
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 27948 15116 28365 15144
rect 27948 15104 27954 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 28353 15107 28411 15113
rect 28442 15104 28448 15156
rect 28500 15104 28506 15156
rect 26970 15036 26976 15088
rect 27028 15076 27034 15088
rect 27028 15048 28304 15076
rect 27028 15036 27034 15048
rect 21821 14971 21879 14977
rect 21928 14980 22324 15008
rect 22557 15011 22615 15017
rect 20220 14912 20760 14940
rect 20220 14900 20226 14912
rect 20806 14900 20812 14952
rect 20864 14900 20870 14952
rect 21560 14940 21588 14971
rect 21634 14940 21640 14952
rect 21560 14912 21640 14940
rect 17420 14844 19104 14872
rect 19260 14872 19288 14900
rect 21560 14872 21588 14912
rect 21634 14900 21640 14912
rect 21692 14940 21698 14952
rect 21928 14940 21956 14980
rect 22557 14977 22569 15011
rect 22603 14977 22615 15011
rect 22557 14971 22615 14977
rect 22824 15011 22882 15017
rect 22824 14977 22836 15011
rect 22870 15008 22882 15011
rect 23382 15008 23388 15020
rect 22870 14980 23388 15008
rect 22870 14977 22882 14980
rect 22824 14971 22882 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 24026 14968 24032 15020
rect 24084 15008 24090 15020
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 24084 14980 24225 15008
rect 24084 14968 24090 14980
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 25774 14968 25780 15020
rect 25832 14968 25838 15020
rect 25866 14968 25872 15020
rect 25924 14968 25930 15020
rect 26602 14968 26608 15020
rect 26660 14968 26666 15020
rect 27172 15017 27200 15048
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27246 14968 27252 15020
rect 27304 15008 27310 15020
rect 27433 15011 27491 15017
rect 27433 15008 27445 15011
rect 27304 14980 27445 15008
rect 27304 14968 27310 14980
rect 27433 14977 27445 14980
rect 27479 14977 27491 15011
rect 27433 14971 27491 14977
rect 27522 14968 27528 15020
rect 27580 14968 27586 15020
rect 28276 15017 28304 15048
rect 27709 15011 27767 15017
rect 27709 15008 27721 15011
rect 27632 14980 27721 15008
rect 21692 14912 21956 14940
rect 21692 14900 21698 14912
rect 22002 14900 22008 14952
rect 22060 14900 22066 14952
rect 24394 14900 24400 14952
rect 24452 14900 24458 14952
rect 24949 14943 25007 14949
rect 24949 14909 24961 14943
rect 24995 14909 25007 14943
rect 24949 14903 25007 14909
rect 25133 14943 25191 14949
rect 25133 14909 25145 14943
rect 25179 14940 25191 14943
rect 25792 14940 25820 14968
rect 26053 14943 26111 14949
rect 26053 14940 26065 14943
rect 25179 14912 25728 14940
rect 25792 14912 26065 14940
rect 25179 14909 25191 14912
rect 25133 14903 25191 14909
rect 24964 14872 24992 14903
rect 25700 14881 25728 14912
rect 26053 14909 26065 14912
rect 26099 14909 26111 14943
rect 26053 14903 26111 14909
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14940 26295 14943
rect 27540 14940 27568 14968
rect 27632 14952 27660 14980
rect 27709 14977 27721 14980
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 28261 15011 28319 15017
rect 28261 14977 28273 15011
rect 28307 14977 28319 15011
rect 28460 15008 28488 15104
rect 28537 15011 28595 15017
rect 28537 15008 28549 15011
rect 28460 14980 28549 15008
rect 28261 14971 28319 14977
rect 28537 14977 28549 14980
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 26283 14912 27108 14940
rect 26283 14909 26295 14912
rect 26237 14903 26295 14909
rect 19260 14844 21588 14872
rect 23492 14844 24992 14872
rect 25685 14875 25743 14881
rect 10796 14776 13124 14804
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 14090 14804 14096 14816
rect 13504 14776 14096 14804
rect 13504 14764 13510 14776
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 17954 14764 17960 14816
rect 18012 14764 18018 14816
rect 18506 14764 18512 14816
rect 18564 14764 18570 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 20990 14804 20996 14816
rect 19659 14776 20996 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 22465 14807 22523 14813
rect 22465 14773 22477 14807
rect 22511 14804 22523 14807
rect 22922 14804 22928 14816
rect 22511 14776 22928 14804
rect 22511 14773 22523 14776
rect 22465 14767 22523 14773
rect 22922 14764 22928 14776
rect 22980 14804 22986 14816
rect 23492 14804 23520 14844
rect 25685 14841 25697 14875
rect 25731 14841 25743 14875
rect 25685 14835 25743 14841
rect 22980 14776 23520 14804
rect 23937 14807 23995 14813
rect 22980 14764 22986 14776
rect 23937 14773 23949 14807
rect 23983 14804 23995 14807
rect 24026 14804 24032 14816
rect 23983 14776 24032 14804
rect 23983 14773 23995 14776
rect 23937 14767 23995 14773
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24857 14807 24915 14813
rect 24857 14773 24869 14807
rect 24903 14804 24915 14807
rect 24946 14804 24952 14816
rect 24903 14776 24952 14804
rect 24903 14773 24915 14776
rect 24857 14767 24915 14773
rect 24946 14764 24952 14776
rect 25004 14804 25010 14816
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 25004 14776 25329 14804
rect 25004 14764 25010 14776
rect 25317 14773 25329 14776
rect 25363 14773 25375 14807
rect 25317 14767 25375 14773
rect 26970 14764 26976 14816
rect 27028 14764 27034 14816
rect 27080 14804 27108 14912
rect 27264 14912 27568 14940
rect 27264 14881 27292 14912
rect 27614 14900 27620 14952
rect 27672 14900 27678 14952
rect 28000 14940 28028 14971
rect 27724 14912 28028 14940
rect 28276 14940 28304 14971
rect 28276 14912 28580 14940
rect 27249 14875 27307 14881
rect 27249 14841 27261 14875
rect 27295 14841 27307 14875
rect 27249 14835 27307 14841
rect 27525 14875 27583 14881
rect 27525 14841 27537 14875
rect 27571 14872 27583 14875
rect 27724 14872 27752 14912
rect 27571 14844 27752 14872
rect 27571 14841 27583 14844
rect 27525 14835 27583 14841
rect 28552 14816 28580 14912
rect 27801 14807 27859 14813
rect 27801 14804 27813 14807
rect 27080 14776 27813 14804
rect 27801 14773 27813 14776
rect 27847 14773 27859 14807
rect 27801 14767 27859 14773
rect 28074 14764 28080 14816
rect 28132 14764 28138 14816
rect 28534 14764 28540 14816
rect 28592 14764 28598 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 2866 14600 2872 14612
rect 2363 14572 2872 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3142 14560 3148 14612
rect 3200 14560 3206 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3326 14600 3332 14612
rect 3283 14572 3332 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 4338 14560 4344 14612
rect 4396 14560 4402 14612
rect 4816 14572 7880 14600
rect 2958 14532 2964 14544
rect 1688 14504 2964 14532
rect 1688 14405 1716 14504
rect 2958 14492 2964 14504
rect 3016 14492 3022 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 3988 14504 4537 14532
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2501 14467 2559 14473
rect 2501 14464 2513 14467
rect 2087 14436 2513 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2501 14433 2513 14436
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 3050 14464 3056 14476
rect 2731 14436 3056 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3988 14473 4016 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 3789 14467 3847 14473
rect 3789 14464 3801 14467
rect 3252 14436 3801 14464
rect 3252 14408 3280 14436
rect 3789 14433 3801 14436
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 1964 14328 1992 14359
rect 2222 14356 2228 14408
rect 2280 14356 2286 14408
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 3418 14356 3424 14408
rect 3476 14356 3482 14408
rect 4172 14396 4200 14424
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4172 14368 4721 14396
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 2314 14328 2320 14340
rect 1964 14300 2320 14328
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 3436 14328 3464 14356
rect 4062 14328 4068 14340
rect 3436 14300 4068 14328
rect 4062 14288 4068 14300
rect 4120 14328 4126 14340
rect 4816 14328 4844 14572
rect 7852 14532 7880 14572
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8076 14572 8401 14600
rect 8076 14560 8082 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 10042 14600 10048 14612
rect 8389 14563 8447 14569
rect 8496 14572 10048 14600
rect 8496 14532 8524 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10686 14560 10692 14612
rect 10744 14560 10750 14612
rect 12069 14603 12127 14609
rect 12069 14569 12081 14603
rect 12115 14600 12127 14603
rect 12342 14600 12348 14612
rect 12115 14572 12348 14600
rect 12115 14569 12127 14572
rect 12069 14563 12127 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14600 13047 14603
rect 13722 14600 13728 14612
rect 13035 14572 13728 14600
rect 13035 14569 13047 14572
rect 12989 14563 13047 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 13906 14560 13912 14612
rect 13964 14560 13970 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 16577 14603 16635 14609
rect 16577 14600 16589 14603
rect 14056 14572 16589 14600
rect 14056 14560 14062 14572
rect 16577 14569 16589 14572
rect 16623 14600 16635 14603
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 16623 14572 17141 14600
rect 16623 14569 16635 14572
rect 16577 14563 16635 14569
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17129 14563 17187 14569
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 18288 14572 18521 14600
rect 18288 14560 18294 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19337 14603 19395 14609
rect 19337 14600 19349 14603
rect 19208 14572 19349 14600
rect 19208 14560 19214 14572
rect 19337 14569 19349 14572
rect 19383 14569 19395 14603
rect 19337 14563 19395 14569
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 20070 14600 20076 14612
rect 19935 14572 20076 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20165 14603 20223 14609
rect 20165 14569 20177 14603
rect 20211 14569 20223 14603
rect 20165 14563 20223 14569
rect 20441 14603 20499 14609
rect 20441 14569 20453 14603
rect 20487 14600 20499 14603
rect 20806 14600 20812 14612
rect 20487 14572 20812 14600
rect 20487 14569 20499 14572
rect 20441 14563 20499 14569
rect 7852 14504 8524 14532
rect 6362 14424 6368 14476
rect 6420 14464 6426 14476
rect 6420 14436 7052 14464
rect 6420 14424 6426 14436
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 4120 14300 4844 14328
rect 5092 14328 5120 14359
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 5316 14368 6929 14396
rect 5316 14356 5322 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 7024 14396 7052 14436
rect 7944 14436 8708 14464
rect 7944 14396 7972 14436
rect 7024 14368 7972 14396
rect 8573 14399 8631 14405
rect 6917 14359 6975 14365
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 5350 14328 5356 14340
rect 5092 14300 5356 14328
rect 4120 14288 4126 14300
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 5525 14337 5531 14340
rect 5517 14331 5531 14337
rect 5517 14297 5529 14331
rect 5517 14291 5531 14297
rect 5525 14288 5531 14291
rect 5583 14288 5589 14340
rect 7184 14331 7242 14337
rect 7184 14297 7196 14331
rect 7230 14328 7242 14331
rect 7558 14328 7564 14340
rect 7230 14300 7564 14328
rect 7230 14297 7242 14300
rect 7184 14291 7242 14297
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 8588 14272 8616 14359
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14260 1823 14263
rect 2038 14260 2044 14272
rect 1811 14232 2044 14260
rect 1811 14229 1823 14232
rect 1765 14223 1823 14229
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5810 14260 5816 14272
rect 4939 14232 5816 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 6730 14260 6736 14272
rect 6687 14232 6736 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8570 14260 8576 14272
rect 8343 14232 8576 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 8680 14260 8708 14436
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10284 14436 10425 14464
rect 10284 14424 10290 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10704 14464 10732 14560
rect 13446 14532 13452 14544
rect 13188 14504 13452 14532
rect 10643 14436 10732 14464
rect 11808 14436 12112 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 10134 14396 10140 14408
rect 8987 14368 10140 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 11808 14405 11836 14436
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 11072 14368 11161 14396
rect 9208 14331 9266 14337
rect 9208 14297 9220 14331
rect 9254 14328 9266 14331
rect 9950 14328 9956 14340
rect 9254 14300 9956 14328
rect 9254 14297 9266 14300
rect 9208 14291 9266 14297
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 10226 14260 10232 14272
rect 8680 14232 10232 14260
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 10318 14220 10324 14272
rect 10376 14220 10382 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11072 14269 11100 14368
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11985 14399 12043 14405
rect 11985 14365 11997 14399
rect 12031 14365 12043 14399
rect 12084 14396 12112 14436
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 12437 14467 12495 14473
rect 12437 14464 12449 14467
rect 12400 14436 12449 14464
rect 12400 14424 12406 14436
rect 12437 14433 12449 14436
rect 12483 14433 12495 14467
rect 12437 14427 12495 14433
rect 12158 14396 12164 14408
rect 12084 14368 12164 14396
rect 11985 14359 12043 14365
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10928 14232 11069 14260
rect 10928 14220 10934 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11348 14260 11376 14359
rect 11992 14328 12020 14359
rect 12158 14356 12164 14368
rect 12216 14396 12222 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12216 14368 12265 14396
rect 12216 14356 12222 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 13078 14396 13084 14408
rect 12253 14359 12311 14365
rect 12406 14368 13084 14396
rect 12406 14328 12434 14368
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13188 14405 13216 14504
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 16114 14492 16120 14544
rect 16172 14532 16178 14544
rect 19426 14532 19432 14544
rect 16172 14504 19432 14532
rect 16172 14492 16178 14504
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 19613 14535 19671 14541
rect 19613 14501 19625 14535
rect 19659 14501 19671 14535
rect 19613 14495 19671 14501
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 15286 14424 15292 14476
rect 15344 14464 15350 14476
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15344 14436 16221 14464
rect 15344 14424 15350 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17184 14436 17509 14464
rect 17184 14424 17190 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 17497 14427 17555 14433
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 19150 14464 19156 14476
rect 18196 14436 19156 14464
rect 18196 14424 18202 14436
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14108 14328 14136 14359
rect 16022 14356 16028 14408
rect 16080 14356 16086 14408
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 11992 14300 12434 14328
rect 12912 14300 14136 14328
rect 14277 14331 14335 14337
rect 12912 14272 12940 14300
rect 14277 14297 14289 14331
rect 14323 14297 14335 14331
rect 16960 14328 16988 14359
rect 17678 14356 17684 14408
rect 17736 14356 17742 14408
rect 18432 14405 18460 14436
rect 19150 14424 19156 14436
rect 19208 14464 19214 14476
rect 19628 14464 19656 14495
rect 20180 14464 20208 14563
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 22002 14560 22008 14612
rect 22060 14600 22066 14612
rect 22465 14603 22523 14609
rect 22465 14600 22477 14603
rect 22060 14572 22477 14600
rect 22060 14560 22066 14572
rect 22465 14569 22477 14572
rect 22511 14569 22523 14603
rect 22465 14563 22523 14569
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22612 14572 22845 14600
rect 22612 14560 22618 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 24394 14560 24400 14612
rect 24452 14600 24458 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 24452 14572 25053 14600
rect 24452 14560 24458 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25866 14600 25872 14612
rect 25041 14563 25099 14569
rect 25148 14572 25872 14600
rect 20717 14535 20775 14541
rect 20717 14501 20729 14535
rect 20763 14501 20775 14535
rect 20717 14495 20775 14501
rect 20732 14464 20760 14495
rect 22646 14492 22652 14544
rect 22704 14492 22710 14544
rect 24029 14535 24087 14541
rect 24029 14501 24041 14535
rect 24075 14532 24087 14535
rect 25148 14532 25176 14572
rect 25866 14560 25872 14572
rect 25924 14560 25930 14612
rect 26602 14560 26608 14612
rect 26660 14560 26666 14612
rect 26970 14560 26976 14612
rect 27028 14560 27034 14612
rect 27430 14560 27436 14612
rect 27488 14560 27494 14612
rect 24075 14504 25176 14532
rect 24075 14501 24087 14504
rect 24029 14495 24087 14501
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 19208 14436 19564 14464
rect 19628 14436 20116 14464
rect 20180 14436 20668 14464
rect 20732 14436 21189 14464
rect 19208 14424 19214 14436
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 18708 14328 18736 14359
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 18966 14396 18972 14408
rect 18840 14368 18972 14396
rect 18840 14356 18846 14368
rect 18966 14356 18972 14368
rect 19024 14396 19030 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19024 14368 19257 14396
rect 19024 14356 19030 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19536 14396 19564 14436
rect 20088 14405 20116 14436
rect 20640 14405 20668 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 21266 14424 21272 14476
rect 21324 14464 21330 14476
rect 21729 14467 21787 14473
rect 21729 14464 21741 14467
rect 21324 14436 21741 14464
rect 21324 14424 21330 14436
rect 21729 14433 21741 14436
rect 21775 14433 21787 14467
rect 22278 14464 22284 14476
rect 21729 14427 21787 14433
rect 21836 14436 22284 14464
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19536 14368 19809 14396
rect 19245 14359 19303 14365
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 20625 14399 20683 14405
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 14277 14291 14335 14297
rect 16040 14300 16988 14328
rect 18248 14300 18736 14328
rect 19260 14328 19288 14359
rect 20364 14328 20392 14359
rect 20898 14356 20904 14408
rect 20956 14356 20962 14408
rect 20990 14356 20996 14408
rect 21048 14356 21054 14408
rect 21836 14396 21864 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 22664 14464 22692 14492
rect 22664 14436 22784 14464
rect 22756 14405 22784 14436
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 25225 14467 25283 14473
rect 25225 14464 25237 14467
rect 25188 14436 25237 14464
rect 25188 14424 25194 14436
rect 25225 14433 25237 14436
rect 25271 14433 25283 14467
rect 25225 14427 25283 14433
rect 21100 14368 21864 14396
rect 21913 14399 21971 14405
rect 19260 14300 20392 14328
rect 12250 14260 12256 14272
rect 11348 14232 12256 14260
rect 11057 14223 11115 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12894 14220 12900 14272
rect 12952 14220 12958 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14292 14260 14320 14291
rect 14240 14232 14320 14260
rect 14240 14220 14246 14232
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16040 14260 16068 14300
rect 18248 14269 18276 14300
rect 15896 14232 16068 14260
rect 18233 14263 18291 14269
rect 15896 14220 15902 14232
rect 18233 14229 18245 14263
rect 18279 14229 18291 14263
rect 18233 14223 18291 14229
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 21100 14260 21128 14368
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14396 22799 14399
rect 23014 14396 23020 14408
rect 22787 14368 23020 14396
rect 22787 14365 22799 14368
rect 22741 14359 22799 14365
rect 21450 14288 21456 14340
rect 21508 14328 21514 14340
rect 21928 14328 21956 14359
rect 21508 14300 21956 14328
rect 22664 14328 22692 14359
rect 23014 14356 23020 14368
rect 23072 14356 23078 14408
rect 23106 14356 23112 14408
rect 23164 14356 23170 14408
rect 23198 14356 23204 14408
rect 23256 14356 23262 14408
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24213 14399 24271 14405
rect 24213 14396 24225 14399
rect 24084 14368 24225 14396
rect 24084 14356 24090 14368
rect 24213 14365 24225 14368
rect 24259 14396 24271 14399
rect 24949 14399 25007 14405
rect 24949 14396 24961 14399
rect 24259 14368 24961 14396
rect 24259 14365 24271 14368
rect 24213 14359 24271 14365
rect 24949 14365 24961 14368
rect 24995 14396 25007 14399
rect 24995 14368 25268 14396
rect 24995 14365 25007 14368
rect 24949 14359 25007 14365
rect 23124 14328 23152 14356
rect 22664 14300 23152 14328
rect 21508 14288 21514 14300
rect 19484 14232 21128 14260
rect 19484 14220 19490 14232
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 22373 14263 22431 14269
rect 22373 14260 22385 14263
rect 21692 14232 22385 14260
rect 21692 14220 21698 14232
rect 22373 14229 22385 14232
rect 22419 14229 22431 14263
rect 23216 14260 23244 14356
rect 25240 14340 25268 14368
rect 25314 14356 25320 14408
rect 25372 14396 25378 14408
rect 26697 14399 26755 14405
rect 26697 14396 26709 14399
rect 25372 14368 26709 14396
rect 25372 14356 25378 14368
rect 26697 14365 26709 14368
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 26881 14399 26939 14405
rect 26881 14365 26893 14399
rect 26927 14365 26939 14399
rect 26988 14396 27016 14560
rect 27338 14492 27344 14544
rect 27396 14532 27402 14544
rect 28077 14535 28135 14541
rect 28077 14532 28089 14535
rect 27396 14504 28089 14532
rect 27396 14492 27402 14504
rect 28077 14501 28089 14504
rect 28123 14501 28135 14535
rect 28077 14495 28135 14501
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 27709 14467 27767 14473
rect 27709 14464 27721 14467
rect 27580 14436 27721 14464
rect 27580 14424 27586 14436
rect 27709 14433 27721 14436
rect 27755 14464 27767 14467
rect 27798 14464 27804 14476
rect 27755 14436 27804 14464
rect 27755 14433 27767 14436
rect 27709 14427 27767 14433
rect 27798 14424 27804 14436
rect 27856 14424 27862 14476
rect 27617 14399 27675 14405
rect 27617 14396 27629 14399
rect 26988 14368 27629 14396
rect 26881 14359 26939 14365
rect 27617 14365 27629 14368
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 27893 14399 27951 14405
rect 27893 14365 27905 14399
rect 27939 14396 27951 14399
rect 28166 14396 28172 14408
rect 27939 14368 28172 14396
rect 27939 14365 27951 14368
rect 27893 14359 27951 14365
rect 24486 14288 24492 14340
rect 24544 14288 24550 14340
rect 25222 14288 25228 14340
rect 25280 14288 25286 14340
rect 25492 14331 25550 14337
rect 25492 14297 25504 14331
rect 25538 14328 25550 14331
rect 26418 14328 26424 14340
rect 25538 14300 26424 14328
rect 25538 14297 25550 14300
rect 25492 14291 25550 14297
rect 26418 14288 26424 14300
rect 26476 14288 26482 14340
rect 26896 14328 26924 14359
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 28442 14328 28448 14340
rect 26896 14300 28448 14328
rect 28442 14288 28448 14300
rect 28500 14288 28506 14340
rect 23290 14260 23296 14272
rect 23216 14232 23296 14260
rect 22373 14223 22431 14229
rect 23290 14220 23296 14232
rect 23348 14260 23354 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 23348 14232 24593 14260
rect 23348 14220 23354 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2372 14028 2789 14056
rect 2372 14016 2378 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 2777 14019 2835 14025
rect 3694 14016 3700 14068
rect 3752 14016 3758 14068
rect 4062 14016 4068 14068
rect 4120 14016 4126 14068
rect 4798 14016 4804 14068
rect 4856 14016 4862 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 7190 14056 7196 14068
rect 6687 14028 7196 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 7558 14016 7564 14068
rect 7616 14016 7622 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8386 14056 8392 14068
rect 8159 14028 8392 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 10870 14016 10876 14068
rect 10928 14016 10934 14068
rect 12158 14016 12164 14068
rect 12216 14016 12222 14068
rect 12250 14016 12256 14068
rect 12308 14016 12314 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 12952 14028 13185 14056
rect 12952 14016 12958 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 13173 14019 13231 14025
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14274 14056 14280 14068
rect 13412 14028 14280 14056
rect 13412 14016 13418 14028
rect 14274 14016 14280 14028
rect 14332 14056 14338 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 14332 14028 14657 14056
rect 14332 14016 14338 14028
rect 14645 14025 14657 14028
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15838 14056 15844 14068
rect 15151 14028 15844 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 1664 13923 1722 13929
rect 1664 13889 1676 13923
rect 1710 13920 1722 13923
rect 2774 13920 2780 13932
rect 1710 13892 2780 13920
rect 1710 13889 1722 13892
rect 1664 13883 1722 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3712 13920 3740 14016
rect 4080 13929 4108 14016
rect 4246 13948 4252 14000
rect 4304 13988 4310 14000
rect 4816 13988 4844 14016
rect 6457 13991 6515 13997
rect 4304 13960 6408 13988
rect 4304 13948 4310 13960
rect 6380 13932 6408 13960
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 6914 13988 6920 14000
rect 6503 13960 6920 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 9490 13988 9496 14000
rect 7432 13960 9496 13988
rect 7432 13948 7438 13960
rect 9490 13948 9496 13960
rect 9548 13988 9554 14000
rect 9548 13960 9720 13988
rect 9548 13948 9554 13960
rect 3651 13892 3740 13920
rect 4065 13923 4123 13929
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4212 13892 4445 13920
rect 4212 13880 4218 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4982 13920 4988 13932
rect 4433 13883 4491 13889
rect 4724 13892 4988 13920
rect 1394 13812 1400 13864
rect 1452 13812 1458 13864
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13852 3111 13855
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3099 13824 3709 13852
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4724 13852 4752 13892
rect 4982 13880 4988 13892
rect 5040 13920 5046 13932
rect 5040 13892 5212 13920
rect 5040 13880 5046 13892
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4295 13824 4752 13852
rect 4816 13824 5089 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4816 13728 4844 13824
rect 5077 13821 5089 13824
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 5184 13784 5212 13892
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5902 13920 5908 13932
rect 5408 13892 5908 13920
rect 5408 13880 5414 13892
rect 5902 13880 5908 13892
rect 5960 13920 5966 13932
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5960 13892 6009 13920
rect 5960 13880 5966 13892
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6362 13880 6368 13932
rect 6420 13880 6426 13932
rect 6822 13880 6828 13932
rect 6880 13880 6886 13932
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 7883 13892 7972 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5626 13852 5632 13864
rect 5307 13824 5632 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6788 13824 7021 13852
rect 6788 13812 6794 13824
rect 7009 13821 7021 13824
rect 7055 13852 7067 13855
rect 7944 13852 7972 13892
rect 8018 13880 8024 13932
rect 8076 13880 8082 13932
rect 9692 13920 9720 13960
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 10192 13960 13308 13988
rect 10192 13948 10198 13960
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9692 13892 10241 13920
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 13280 13929 13308 13960
rect 14182 13948 14188 14000
rect 14240 13948 14246 14000
rect 14660 13988 14688 14019
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16022 14016 16028 14068
rect 16080 14056 16086 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 16080 14028 16129 14056
rect 16080 14016 16086 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 15948 13988 15976 14016
rect 14660 13960 15056 13988
rect 13538 13929 13544 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 11020 13892 11345 13920
rect 11020 13880 11026 13892
rect 11333 13889 11345 13892
rect 11379 13889 11391 13923
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 11333 13883 11391 13889
rect 11440 13892 12449 13920
rect 8110 13852 8116 13864
rect 7055 13824 7880 13852
rect 7944 13824 8116 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 7374 13784 7380 13796
rect 5184 13756 7380 13784
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 7852 13728 7880 13824
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8312 13784 8340 13815
rect 8478 13812 8484 13864
rect 8536 13812 8542 13864
rect 10042 13812 10048 13864
rect 10100 13812 10106 13864
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11440 13852 11468 13892
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13532 13883 13544 13929
rect 13538 13880 13544 13883
rect 13596 13880 13602 13932
rect 14200 13920 14228 13948
rect 15028 13929 15056 13960
rect 15488 13960 15976 13988
rect 15488 13929 15516 13960
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14200 13892 14933 13920
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 16224 13920 16252 14019
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17402 14056 17408 14068
rect 16632 14028 17408 14056
rect 16632 14016 16638 14028
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 17589 14059 17647 14065
rect 17589 14056 17601 14059
rect 17460 14028 17601 14056
rect 17460 14016 17466 14028
rect 17589 14025 17601 14028
rect 17635 14025 17647 14059
rect 17589 14019 17647 14025
rect 17678 14016 17684 14068
rect 17736 14056 17742 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 17736 14028 18061 14056
rect 17736 14016 17742 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18432 14028 20852 14056
rect 17497 13991 17555 13997
rect 17497 13957 17509 13991
rect 17543 13988 17555 13991
rect 18432 13988 18460 14028
rect 17543 13960 18460 13988
rect 17543 13957 17555 13960
rect 17497 13951 17555 13957
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19880 13991 19938 13997
rect 19024 13960 19564 13988
rect 19024 13948 19030 13960
rect 15703 13892 16252 13920
rect 16393 13923 16451 13929
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 16393 13889 16405 13923
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 11164 13824 11468 13852
rect 11517 13855 11575 13861
rect 7944 13756 8340 13784
rect 7944 13728 7972 13756
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 10502 13784 10508 13796
rect 9088 13756 10508 13784
rect 9088 13744 9094 13756
rect 10502 13744 10508 13756
rect 10560 13744 10566 13796
rect 11164 13793 11192 13824
rect 11517 13821 11529 13855
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 11701 13855 11759 13861
rect 11701 13821 11713 13855
rect 11747 13852 11759 13855
rect 11790 13852 11796 13864
rect 11747 13824 11796 13852
rect 11747 13821 11759 13824
rect 11701 13815 11759 13821
rect 11149 13787 11207 13793
rect 11149 13753 11161 13787
rect 11195 13753 11207 13787
rect 11149 13747 11207 13753
rect 3234 13676 3240 13728
rect 3292 13676 3298 13728
rect 3602 13676 3608 13728
rect 3660 13716 3666 13728
rect 3881 13719 3939 13725
rect 3881 13716 3893 13719
rect 3660 13688 3893 13716
rect 3660 13676 3666 13688
rect 3881 13685 3893 13688
rect 3927 13685 3939 13719
rect 3881 13679 3939 13685
rect 4798 13676 4804 13728
rect 4856 13676 4862 13728
rect 5718 13676 5724 13728
rect 5776 13676 5782 13728
rect 6086 13676 6092 13728
rect 6144 13676 6150 13728
rect 7650 13676 7656 13728
rect 7708 13676 7714 13728
rect 7834 13676 7840 13728
rect 7892 13676 7898 13728
rect 7926 13676 7932 13728
rect 7984 13676 7990 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11532 13716 11560 13815
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12526 13812 12532 13864
rect 12584 13812 12590 13864
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 16408 13852 16436 13883
rect 14752 13824 16436 13852
rect 14752 13793 14780 13824
rect 17972 13796 18000 13883
rect 18532 13852 18560 13883
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 19536 13929 19564 13960
rect 19880 13957 19892 13991
rect 19926 13988 19938 13991
rect 19978 13988 19984 14000
rect 19926 13960 19984 13988
rect 19926 13957 19938 13960
rect 19880 13951 19938 13957
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20824 13988 20852 14028
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 20956 14028 21097 14056
rect 20956 14016 20962 14028
rect 21085 14025 21097 14028
rect 21131 14025 21143 14059
rect 21085 14019 21143 14025
rect 21450 14016 21456 14068
rect 21508 14016 21514 14068
rect 27798 14056 27804 14068
rect 24136 14028 27804 14056
rect 24136 13997 24164 14028
rect 27798 14016 27804 14028
rect 27856 14016 27862 14068
rect 28350 14016 28356 14068
rect 28408 14056 28414 14068
rect 28445 14059 28503 14065
rect 28445 14056 28457 14059
rect 28408 14028 28457 14056
rect 28408 14016 28414 14028
rect 28445 14025 28457 14028
rect 28491 14025 28503 14059
rect 28445 14019 28503 14025
rect 24121 13991 24179 13997
rect 20824 13960 24072 13988
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19521 13923 19579 13929
rect 18831 13892 19380 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 18708 13852 18736 13880
rect 18532 13824 18736 13852
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 14737 13787 14795 13793
rect 14737 13753 14749 13787
rect 14783 13753 14795 13787
rect 14737 13747 14795 13753
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18892 13784 18920 13812
rect 19352 13793 19380 13892
rect 19521 13889 19533 13923
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19610 13880 19616 13932
rect 19668 13880 19674 13932
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13920 21327 13923
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 21315 13892 21373 13920
rect 21315 13889 21327 13892
rect 21269 13883 21327 13889
rect 21361 13889 21373 13892
rect 21407 13920 21419 13923
rect 21450 13920 21456 13932
rect 21407 13892 21456 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 18012 13756 18920 13784
rect 19337 13787 19395 13793
rect 18012 13744 18018 13756
rect 19337 13753 19349 13787
rect 19383 13753 19395 13787
rect 19337 13747 19395 13753
rect 20993 13787 21051 13793
rect 20993 13753 21005 13787
rect 21039 13784 21051 13787
rect 21284 13784 21312 13883
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 22922 13920 22928 13932
rect 22235 13892 22928 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 23014 13880 23020 13932
rect 23072 13880 23078 13932
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13920 23167 13923
rect 23477 13923 23535 13929
rect 23477 13920 23489 13923
rect 23155 13892 23489 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 23477 13889 23489 13892
rect 23523 13889 23535 13923
rect 24044 13920 24072 13960
rect 24121 13957 24133 13991
rect 24167 13957 24179 13991
rect 27614 13988 27620 14000
rect 24121 13951 24179 13957
rect 26252 13960 26464 13988
rect 26252 13932 26280 13960
rect 24044 13892 24532 13920
rect 23477 13883 23535 13889
rect 21542 13812 21548 13864
rect 21600 13852 21606 13864
rect 23293 13855 23351 13861
rect 23293 13852 23305 13855
rect 21600 13824 23305 13852
rect 21600 13812 21606 13824
rect 23293 13821 23305 13824
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 24504 13852 24532 13892
rect 24578 13880 24584 13932
rect 24636 13880 24642 13932
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25774 13880 25780 13932
rect 25832 13880 25838 13932
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13920 25927 13923
rect 26234 13920 26240 13932
rect 25915 13892 26240 13920
rect 25915 13889 25927 13892
rect 25869 13883 25927 13889
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 26326 13880 26332 13932
rect 26384 13880 26390 13932
rect 26436 13929 26464 13960
rect 27080 13960 27620 13988
rect 27080 13932 27108 13960
rect 27614 13948 27620 13960
rect 27672 13988 27678 14000
rect 27672 13960 28396 13988
rect 27672 13948 27678 13960
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 27062 13880 27068 13932
rect 27120 13880 27126 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27525 13923 27583 13929
rect 27525 13920 27537 13923
rect 27203 13892 27537 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 27525 13889 27537 13892
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 28368 13929 28396 13960
rect 28261 13923 28319 13929
rect 28261 13920 28273 13923
rect 28132 13892 28273 13920
rect 28132 13880 28138 13892
rect 28261 13889 28273 13892
rect 28307 13889 28319 13923
rect 28261 13883 28319 13889
rect 28353 13923 28411 13929
rect 28353 13889 28365 13923
rect 28399 13889 28411 13923
rect 28353 13883 28411 13889
rect 25792 13852 25820 13880
rect 24504 13824 25820 13852
rect 27338 13812 27344 13864
rect 27396 13812 27402 13864
rect 27982 13812 27988 13864
rect 28040 13812 28046 13864
rect 28166 13852 28172 13864
rect 28092 13824 28172 13852
rect 21039 13756 21312 13784
rect 21039 13753 21051 13756
rect 20993 13747 21051 13753
rect 11112 13688 11560 13716
rect 11112 13676 11118 13688
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 16574 13716 16580 13728
rect 12492 13688 16580 13716
rect 12492 13676 12498 13688
rect 16574 13676 16580 13688
rect 16632 13676 16638 13728
rect 18325 13719 18383 13725
rect 18325 13685 18337 13719
rect 18371 13716 18383 13719
rect 18966 13716 18972 13728
rect 18371 13688 18972 13716
rect 18371 13685 18383 13688
rect 18325 13679 18383 13685
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19245 13719 19303 13725
rect 19245 13685 19257 13719
rect 19291 13716 19303 13719
rect 19610 13716 19616 13728
rect 19291 13688 19616 13716
rect 19291 13685 19303 13688
rect 19245 13679 19303 13685
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 21560 13716 21588 13812
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 22830 13784 22836 13796
rect 22244 13756 22836 13784
rect 22244 13744 22250 13756
rect 22830 13744 22836 13756
rect 22888 13784 22894 13796
rect 28092 13793 28120 13824
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 28077 13787 28135 13793
rect 22888 13756 25360 13784
rect 22888 13744 22894 13756
rect 25332 13728 25360 13756
rect 28077 13753 28089 13787
rect 28123 13753 28135 13787
rect 28077 13747 28135 13753
rect 20588 13688 21588 13716
rect 22005 13719 22063 13725
rect 20588 13676 20594 13688
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 22554 13716 22560 13728
rect 22051 13688 22560 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 23658 13676 23664 13728
rect 23716 13676 23722 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 25314 13676 25320 13728
rect 25372 13676 25378 13728
rect 25774 13676 25780 13728
rect 25832 13676 25838 13728
rect 25958 13676 25964 13728
rect 26016 13676 26022 13728
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 26513 13719 26571 13725
rect 26513 13685 26525 13719
rect 26559 13716 26571 13719
rect 26602 13716 26608 13728
rect 26559 13688 26608 13716
rect 26559 13685 26571 13688
rect 26513 13679 26571 13685
rect 26602 13676 26608 13688
rect 26660 13676 26666 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 2774 13472 2780 13524
rect 2832 13472 2838 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 2924 13484 3893 13512
rect 2924 13472 2930 13484
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 3881 13475 3939 13481
rect 4798 13472 4804 13524
rect 4856 13472 4862 13524
rect 5534 13472 5540 13524
rect 5592 13472 5598 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5776 13484 6009 13512
rect 5776 13472 5782 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7926 13512 7932 13524
rect 7147 13484 7932 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13413 1823 13447
rect 2792 13444 2820 13472
rect 3421 13447 3479 13453
rect 3421 13444 3433 13447
rect 2792 13416 3433 13444
rect 1765 13407 1823 13413
rect 3421 13413 3433 13416
rect 3467 13413 3479 13447
rect 6012 13444 6040 13475
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 8168 13484 8309 13512
rect 8168 13472 8174 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 8297 13475 8355 13481
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 9950 13472 9956 13524
rect 10008 13472 10014 13524
rect 10410 13472 10416 13524
rect 10468 13472 10474 13524
rect 10502 13472 10508 13524
rect 10560 13472 10566 13524
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12584 13484 12725 13512
rect 12584 13472 12590 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13596 13484 13737 13512
rect 13596 13472 13602 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 16022 13472 16028 13524
rect 16080 13472 16086 13524
rect 19610 13472 19616 13524
rect 19668 13472 19674 13524
rect 19886 13472 19892 13524
rect 19944 13512 19950 13524
rect 20438 13512 20444 13524
rect 19944 13484 20444 13512
rect 19944 13472 19950 13484
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 22066 13484 23980 13512
rect 7377 13447 7435 13453
rect 3421 13407 3479 13413
rect 4172 13416 5212 13444
rect 6012 13416 6500 13444
rect 1780 13376 1808 13407
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 1780 13348 2237 13376
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 3234 13376 3240 13388
rect 2731 13348 3240 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 4172 13385 4200 13416
rect 5184 13388 5212 13416
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 5166 13336 5172 13388
rect 5224 13336 5230 13388
rect 5350 13336 5356 13388
rect 5408 13336 5414 13388
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 6086 13376 6092 13388
rect 5859 13348 6092 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6472 13385 6500 13416
rect 7377 13413 7389 13447
rect 7423 13444 7435 13447
rect 8496 13444 8524 13472
rect 7423 13416 8524 13444
rect 9125 13447 9183 13453
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 9125 13413 9137 13447
rect 9171 13444 9183 13447
rect 10428 13444 10456 13472
rect 9171 13416 10456 13444
rect 10520 13444 10548 13472
rect 10520 13416 11652 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 7708 13348 7757 13376
rect 7708 13336 7714 13348
rect 7745 13345 7757 13348
rect 7791 13345 7803 13379
rect 9309 13379 9367 13385
rect 9309 13376 9321 13379
rect 7745 13339 7803 13345
rect 8588 13348 9321 13376
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 992 13212 1501 13240
rect 992 13200 998 13212
rect 1489 13209 1501 13212
rect 1535 13209 1547 13243
rect 1964 13240 1992 13271
rect 2038 13268 2044 13320
rect 2096 13268 2102 13320
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 2958 13308 2964 13320
rect 2915 13280 2964 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 2958 13268 2964 13280
rect 3016 13308 3022 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3016 13280 3801 13308
rect 3016 13268 3022 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4338 13268 4344 13320
rect 4396 13268 4402 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5368 13308 5396 13336
rect 8588 13320 8616 13348
rect 9309 13345 9321 13348
rect 9355 13345 9367 13379
rect 9309 13339 9367 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10318 13376 10324 13388
rect 10183 13348 10324 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 4939 13280 5396 13308
rect 5552 13280 5641 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5552 13252 5580 13280
rect 5629 13277 5641 13280
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 6638 13268 6644 13320
rect 6696 13268 6702 13320
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 3602 13240 3608 13252
rect 1964 13212 3608 13240
rect 1489 13203 1547 13209
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 5534 13200 5540 13252
rect 5592 13200 5598 13252
rect 7300 13240 7328 13271
rect 7558 13268 7564 13320
rect 7616 13268 7622 13320
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 8481 13311 8539 13317
rect 8481 13308 8493 13311
rect 7892 13280 8493 13308
rect 7892 13268 7898 13280
rect 8481 13277 8493 13280
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9033 13311 9091 13317
rect 9033 13277 9045 13311
rect 9079 13308 9091 13311
rect 9079 13280 9168 13308
rect 9079 13277 9091 13280
rect 9033 13271 9091 13277
rect 8588 13240 8616 13268
rect 7300 13212 8616 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 6270 13172 6276 13184
rect 1627 13144 6276 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 8772 13172 8800 13271
rect 9140 13240 9168 13280
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 10152 13308 10180 13339
rect 10318 13336 10324 13348
rect 10376 13376 10382 13388
rect 11624 13385 11652 13416
rect 12342 13404 12348 13456
rect 12400 13444 12406 13456
rect 14642 13444 14648 13456
rect 12400 13416 13124 13444
rect 12400 13404 12406 13416
rect 11609 13379 11667 13385
rect 10376 13348 10916 13376
rect 10376 13336 10382 13348
rect 10888 13320 10916 13348
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13376 11851 13379
rect 12894 13376 12900 13388
rect 11839 13348 12900 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 9272 13280 10180 13308
rect 9272 13268 9278 13280
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 10778 13308 10784 13320
rect 10560 13280 10784 13308
rect 10560 13268 10566 13280
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13277 11023 13311
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 10965 13271 11023 13277
rect 12268 13280 12357 13308
rect 9674 13240 9680 13252
rect 9140 13212 9680 13240
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10980 13240 11008 13271
rect 10008 13212 11008 13240
rect 10008 13200 10014 13212
rect 9214 13172 9220 13184
rect 8772 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10689 13175 10747 13181
rect 10689 13172 10701 13175
rect 10100 13144 10701 13172
rect 10100 13132 10106 13144
rect 10689 13141 10701 13144
rect 10735 13141 10747 13175
rect 10689 13135 10747 13141
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 11054 13172 11060 13184
rect 10836 13144 11060 13172
rect 10836 13132 10842 13144
rect 11054 13132 11060 13144
rect 11112 13172 11118 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 11112 13144 11437 13172
rect 11112 13132 11118 13144
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 11425 13135 11483 13141
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12268 13181 12296 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 13096 13308 13124 13416
rect 14384 13416 14648 13444
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 14384 13376 14412 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 16669 13447 16727 13453
rect 16669 13413 16681 13447
rect 16715 13413 16727 13447
rect 16669 13407 16727 13413
rect 16945 13447 17003 13453
rect 16945 13413 16957 13447
rect 16991 13444 17003 13447
rect 18049 13447 18107 13453
rect 16991 13416 17632 13444
rect 16991 13413 17003 13416
rect 16945 13407 17003 13413
rect 13556 13348 14412 13376
rect 14461 13379 14519 13385
rect 13556 13308 13584 13348
rect 14461 13345 14473 13379
rect 14507 13376 14519 13379
rect 14829 13379 14887 13385
rect 14829 13376 14841 13379
rect 14507 13348 14841 13376
rect 14507 13345 14519 13348
rect 14461 13339 14519 13345
rect 14829 13345 14841 13348
rect 14875 13345 14887 13379
rect 14829 13339 14887 13345
rect 15565 13379 15623 13385
rect 15565 13345 15577 13379
rect 15611 13376 15623 13379
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 15611 13348 16221 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 16209 13345 16221 13348
rect 16255 13345 16267 13379
rect 16684 13376 16712 13407
rect 16684 13348 17172 13376
rect 16209 13339 16267 13345
rect 13096 13280 13584 13308
rect 12529 13271 12587 13277
rect 12544 13240 12572 13271
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13688 13280 14289 13308
rect 13688 13268 13694 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 13446 13240 13452 13252
rect 12544 13212 13452 13240
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 14384 13240 14412 13271
rect 14292 13212 14412 13240
rect 14660 13240 14688 13271
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 17144 13317 17172 13348
rect 17402 13336 17408 13388
rect 17460 13336 17466 13388
rect 17604 13385 17632 13416
rect 18049 13413 18061 13447
rect 18095 13444 18107 13447
rect 18509 13447 18567 13453
rect 18509 13444 18521 13447
rect 18095 13416 18521 13444
rect 18095 13413 18107 13416
rect 18049 13407 18107 13413
rect 18509 13413 18521 13416
rect 18555 13413 18567 13447
rect 18509 13407 18567 13413
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15344 13280 15393 13308
rect 15344 13268 15350 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 15562 13240 15568 13252
rect 14660 13212 15568 13240
rect 14292 13184 14320 13212
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 15746 13200 15752 13252
rect 15804 13240 15810 13252
rect 16132 13240 16160 13271
rect 15804 13212 16160 13240
rect 16868 13240 16896 13271
rect 17954 13268 17960 13320
rect 18012 13268 18018 13320
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18230 13308 18236 13320
rect 18187 13280 18236 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 17972 13240 18000 13268
rect 16868 13212 18000 13240
rect 18524 13240 18552 13407
rect 18969 13379 19027 13385
rect 18969 13345 18981 13379
rect 19015 13376 19027 13379
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 19015 13348 19441 13376
rect 19015 13345 19027 13348
rect 18969 13339 19027 13345
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 19628 13376 19656 13472
rect 20990 13404 20996 13456
rect 21048 13444 21054 13456
rect 22066 13444 22094 13484
rect 23952 13456 23980 13484
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24452 13484 24777 13512
rect 24452 13472 24458 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 25038 13472 25044 13524
rect 25096 13512 25102 13524
rect 25498 13512 25504 13524
rect 25096 13484 25504 13512
rect 25096 13472 25102 13484
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 27246 13512 27252 13524
rect 26476 13484 27252 13512
rect 26476 13472 26482 13484
rect 27246 13472 27252 13484
rect 27304 13472 27310 13524
rect 21048 13416 22094 13444
rect 22925 13447 22983 13453
rect 21048 13404 21054 13416
rect 22925 13413 22937 13447
rect 22971 13444 22983 13447
rect 23385 13447 23443 13453
rect 23385 13444 23397 13447
rect 22971 13416 23397 13444
rect 22971 13413 22983 13416
rect 22925 13407 22983 13413
rect 23385 13413 23397 13416
rect 23431 13444 23443 13447
rect 23842 13444 23848 13456
rect 23431 13416 23848 13444
rect 23431 13413 23443 13416
rect 23385 13407 23443 13413
rect 23842 13404 23848 13416
rect 23900 13404 23906 13456
rect 23934 13404 23940 13456
rect 23992 13404 23998 13456
rect 24670 13404 24676 13456
rect 24728 13444 24734 13456
rect 28626 13444 28632 13456
rect 24728 13416 28632 13444
rect 24728 13404 24734 13416
rect 28626 13404 28632 13416
rect 28684 13404 28690 13456
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 19628 13348 20729 13376
rect 19429 13339 19487 13345
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 22278 13336 22284 13388
rect 22336 13336 22342 13388
rect 24121 13379 24179 13385
rect 24121 13345 24133 13379
rect 24167 13376 24179 13379
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24167 13348 24593 13376
rect 24167 13345 24179 13348
rect 24121 13339 24179 13345
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 24946 13336 24952 13388
rect 25004 13376 25010 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 25004 13348 25145 13376
rect 25004 13336 25010 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13376 25375 13379
rect 25958 13376 25964 13388
rect 25363 13348 25964 13376
rect 25363 13345 25375 13348
rect 25317 13339 25375 13345
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 26970 13336 26976 13388
rect 27028 13376 27034 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 27028 13348 27169 13376
rect 27028 13336 27034 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 27157 13339 27215 13345
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18840 13280 18889 13308
rect 18840 13268 18846 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19260 13240 19288 13271
rect 20898 13268 20904 13320
rect 20956 13268 20962 13320
rect 21450 13268 21456 13320
rect 21508 13268 21514 13320
rect 22462 13268 22468 13320
rect 22520 13268 22526 13320
rect 22738 13268 22744 13320
rect 22796 13308 22802 13320
rect 23014 13308 23020 13320
rect 22796 13280 23020 13308
rect 22796 13268 22802 13280
rect 23014 13268 23020 13280
rect 23072 13268 23078 13320
rect 23198 13268 23204 13320
rect 23256 13268 23262 13320
rect 23658 13268 23664 13320
rect 23716 13268 23722 13320
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 24026 13268 24032 13320
rect 24084 13268 24090 13320
rect 24397 13311 24455 13317
rect 24397 13277 24409 13311
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 25869 13311 25927 13317
rect 25869 13277 25881 13311
rect 25915 13308 25927 13311
rect 26234 13308 26240 13320
rect 25915 13280 26240 13308
rect 25915 13277 25927 13280
rect 25869 13271 25927 13277
rect 18524 13212 19288 13240
rect 15804 13200 15810 13212
rect 21266 13200 21272 13252
rect 21324 13240 21330 13252
rect 22097 13243 22155 13249
rect 22097 13240 22109 13243
rect 21324 13212 22109 13240
rect 21324 13200 21330 13212
rect 22097 13209 22109 13212
rect 22143 13209 22155 13243
rect 23676 13240 23704 13268
rect 24412 13240 24440 13271
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 23676 13212 24440 13240
rect 22097 13203 22155 13209
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 12216 13144 12265 13172
rect 12216 13132 12222 13144
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 12253 13135 12311 13141
rect 14090 13132 14096 13184
rect 14148 13132 14154 13184
rect 14274 13132 14280 13184
rect 14332 13132 14338 13184
rect 15580 13172 15608 13200
rect 17402 13172 17408 13184
rect 15580 13144 17408 13172
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20254 13172 20260 13184
rect 20027 13144 20260 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 21358 13132 21364 13184
rect 21416 13132 21422 13184
rect 23750 13132 23756 13184
rect 23808 13132 23814 13184
rect 26510 13132 26516 13184
rect 26568 13132 26574 13184
rect 26712 13172 26740 13271
rect 26881 13243 26939 13249
rect 26881 13209 26893 13243
rect 26927 13240 26939 13243
rect 27890 13240 27896 13252
rect 26927 13212 27896 13240
rect 26927 13209 26939 13212
rect 26881 13203 26939 13209
rect 27890 13200 27896 13212
rect 27948 13200 27954 13252
rect 28074 13172 28080 13184
rect 26712 13144 28080 13172
rect 28074 13132 28080 13144
rect 28132 13132 28138 13184
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 2958 12928 2964 12980
rect 3016 12928 3022 12980
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4154 12968 4160 12980
rect 4019 12940 4160 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4246 12928 4252 12980
rect 4304 12928 4310 12980
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5684 12940 6009 12968
rect 5684 12928 5690 12940
rect 5997 12937 6009 12940
rect 6043 12937 6055 12971
rect 5997 12931 6055 12937
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6638 12968 6644 12980
rect 6595 12940 6644 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7616 12940 8125 12968
rect 7616 12928 7622 12940
rect 8113 12937 8125 12940
rect 8159 12968 8171 12971
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 8159 12940 8953 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 8941 12931 8999 12937
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9950 12968 9956 12980
rect 9263 12940 9956 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12937 10839 12971
rect 10781 12931 10839 12937
rect 1848 12835 1906 12841
rect 1848 12801 1860 12835
rect 1894 12832 1906 12835
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 1894 12804 3709 12832
rect 1894 12801 1906 12804
rect 1848 12795 1906 12801
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4264 12841 4292 12928
rect 5810 12860 5816 12912
rect 5868 12900 5874 12912
rect 8018 12900 8024 12912
rect 5868 12872 6224 12900
rect 5868 12860 5874 12872
rect 6196 12841 6224 12872
rect 6748 12872 8024 12900
rect 4249 12835 4307 12841
rect 4249 12832 4261 12835
rect 3936 12804 4261 12832
rect 3936 12792 3942 12804
rect 4249 12801 4261 12804
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4387 12804 4721 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6638 12832 6644 12844
rect 6503 12804 6644 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 1394 12724 1400 12776
rect 1452 12764 1458 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1452 12736 1593 12764
rect 1452 12724 1458 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 3050 12724 3056 12776
rect 3108 12724 3114 12776
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5074 12764 5080 12776
rect 4571 12736 5080 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 5626 12764 5632 12776
rect 5491 12736 5632 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5276 12696 5304 12727
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 6748 12773 6776 12872
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 10502 12900 10508 12912
rect 8312 12872 10508 12900
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7248 12804 7665 12832
rect 7248 12792 7254 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 8312 12832 8340 12872
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 10796 12900 10824 12931
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11020 12940 12112 12968
rect 11020 12928 11026 12940
rect 10796 12872 11376 12900
rect 7653 12795 7711 12801
rect 8220 12804 8340 12832
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7432 12736 7481 12764
rect 7432 12724 7438 12736
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 5276 12668 5764 12696
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5534 12628 5540 12640
rect 5215 12600 5540 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5534 12588 5540 12600
rect 5592 12628 5598 12640
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5592 12600 5641 12628
rect 5592 12588 5598 12600
rect 5629 12597 5641 12600
rect 5675 12597 5687 12631
rect 5736 12628 5764 12668
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 7190 12696 7196 12708
rect 6328 12668 7196 12696
rect 6328 12656 6334 12668
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 8220 12696 8248 12804
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8444 12804 8493 12832
rect 8444 12792 8450 12804
rect 8481 12801 8493 12804
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8628 12804 9413 12832
rect 8628 12792 8634 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9674 12832 9680 12844
rect 9539 12804 9680 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 10689 12835 10747 12841
rect 9815 12804 10640 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 7300 12668 8248 12696
rect 8312 12696 8340 12727
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9916 12736 10057 12764
rect 9916 12724 9922 12736
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10229 12767 10287 12773
rect 10229 12733 10241 12767
rect 10275 12733 10287 12767
rect 10229 12727 10287 12733
rect 8570 12696 8576 12708
rect 8312 12668 8576 12696
rect 7300 12628 7328 12668
rect 8570 12656 8576 12668
rect 8628 12656 8634 12708
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10244 12696 10272 12727
rect 9631 12668 10272 12696
rect 10612 12696 10640 12804
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 10778 12832 10784 12844
rect 10735 12804 10784 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11348 12841 11376 12872
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10928 12804 10977 12832
rect 10928 12792 10934 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 10962 12696 10968 12708
rect 10612 12668 10968 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11149 12699 11207 12705
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 11716 12696 11744 12727
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 12084 12764 12112 12940
rect 12158 12928 12164 12980
rect 12216 12928 12222 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12710 12968 12716 12980
rect 12299 12940 12716 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 12894 12928 12900 12980
rect 12952 12928 12958 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 13096 12900 13124 12931
rect 13354 12928 13360 12980
rect 13412 12928 13418 12980
rect 13446 12928 13452 12980
rect 13504 12928 13510 12980
rect 13630 12928 13636 12980
rect 13688 12928 13694 12980
rect 14090 12928 14096 12980
rect 14148 12928 14154 12980
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 15473 12971 15531 12977
rect 15473 12937 15485 12971
rect 15519 12937 15531 12971
rect 15473 12931 15531 12937
rect 13372 12900 13400 12928
rect 12452 12872 13124 12900
rect 13280 12872 13400 12900
rect 12452 12841 12480 12872
rect 13280 12841 13308 12872
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 12805 12835 12863 12841
rect 12805 12801 12817 12835
rect 12851 12832 12863 12835
rect 13265 12835 13323 12841
rect 12851 12804 12940 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 12728 12764 12756 12795
rect 12912 12776 12940 12804
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13354 12792 13360 12844
rect 13412 12792 13418 12844
rect 13825 12835 13883 12841
rect 13825 12801 13837 12835
rect 13871 12832 13883 12835
rect 14108 12832 14136 12928
rect 14182 12860 14188 12912
rect 14240 12900 14246 12912
rect 15488 12900 15516 12931
rect 16574 12928 16580 12980
rect 16632 12928 16638 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 16816 12940 17325 12968
rect 16816 12928 16822 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 18322 12968 18328 12980
rect 17635 12940 18328 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21545 12971 21603 12977
rect 21545 12968 21557 12971
rect 20956 12940 21557 12968
rect 20956 12928 20962 12940
rect 21545 12937 21557 12940
rect 21591 12937 21603 12971
rect 22186 12968 22192 12980
rect 21545 12931 21603 12937
rect 21744 12940 22192 12968
rect 16592 12900 16620 12928
rect 21744 12900 21772 12940
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 22462 12968 22468 12980
rect 22419 12940 22468 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 22646 12928 22652 12980
rect 22704 12928 22710 12980
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23198 12968 23204 12980
rect 22787 12940 23204 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 23750 12928 23756 12980
rect 23808 12928 23814 12980
rect 23842 12928 23848 12980
rect 23900 12928 23906 12980
rect 24394 12928 24400 12980
rect 24452 12968 24458 12980
rect 24581 12971 24639 12977
rect 24581 12968 24593 12971
rect 24452 12940 24593 12968
rect 24452 12928 24458 12940
rect 24581 12937 24593 12940
rect 24627 12937 24639 12971
rect 24581 12931 24639 12937
rect 26602 12928 26608 12980
rect 26660 12928 26666 12980
rect 27246 12928 27252 12980
rect 27304 12968 27310 12980
rect 27617 12971 27675 12977
rect 27617 12968 27629 12971
rect 27304 12940 27629 12968
rect 27304 12928 27310 12940
rect 27617 12937 27629 12940
rect 27663 12937 27675 12971
rect 27617 12931 27675 12937
rect 28074 12928 28080 12980
rect 28132 12968 28138 12980
rect 28353 12971 28411 12977
rect 28353 12968 28365 12971
rect 28132 12940 28365 12968
rect 28132 12928 28138 12940
rect 28353 12937 28365 12940
rect 28399 12937 28411 12971
rect 28353 12931 28411 12937
rect 14240 12872 14964 12900
rect 15488 12872 16068 12900
rect 16592 12872 21772 12900
rect 14240 12860 14246 12872
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 13871 12804 13952 12832
rect 14108 12804 14841 12832
rect 13871 12801 13883 12804
rect 13825 12795 13883 12801
rect 12084 12736 12756 12764
rect 11195 12668 11744 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 5736 12600 7328 12628
rect 5629 12591 5687 12597
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12628 9919 12631
rect 11808 12628 11836 12724
rect 12728 12696 12756 12736
rect 12894 12724 12900 12776
rect 12952 12724 12958 12776
rect 13924 12764 13952 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14936 12832 14964 12872
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 14936 12804 15669 12832
rect 14829 12795 14887 12801
rect 15657 12801 15669 12804
rect 15703 12832 15715 12835
rect 15746 12832 15752 12844
rect 15703 12804 15752 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 16040 12841 16068 12872
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 17954 12832 17960 12844
rect 17543 12804 17960 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18874 12832 18880 12844
rect 18340 12804 18880 12832
rect 14274 12764 14280 12776
rect 13924 12736 14280 12764
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 13170 12696 13176 12708
rect 12728 12668 13176 12696
rect 13170 12656 13176 12668
rect 13228 12696 13234 12708
rect 14090 12696 14096 12708
rect 13228 12668 14096 12696
rect 13228 12656 13234 12668
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 9907 12600 11836 12628
rect 9907 12597 9919 12600
rect 9861 12591 9919 12597
rect 12526 12588 12532 12640
rect 12584 12588 12590 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14660 12628 14688 12727
rect 16666 12724 16672 12776
rect 16724 12724 16730 12776
rect 18340 12773 18368 12804
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19076 12841 19104 12872
rect 21818 12860 21824 12912
rect 21876 12900 21882 12912
rect 21876 12872 22324 12900
rect 21876 12860 21882 12872
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 20254 12792 20260 12844
rect 20312 12832 20318 12844
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 20312 12804 20545 12832
rect 20312 12792 20318 12804
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 21450 12792 21456 12844
rect 21508 12832 21514 12844
rect 22296 12841 22324 12872
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21508 12804 22017 12832
rect 21508 12792 21514 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 22664 12841 22692 12928
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 22922 12792 22928 12844
rect 22980 12832 22986 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22980 12804 23121 12832
rect 22980 12792 22986 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 23290 12832 23296 12844
rect 23247 12804 23296 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 23385 12835 23443 12841
rect 23385 12801 23397 12835
rect 23431 12832 23443 12835
rect 23768 12832 23796 12928
rect 23431 12804 23796 12832
rect 23860 12832 23888 12928
rect 25400 12903 25458 12909
rect 25400 12869 25412 12903
rect 25446 12900 25458 12903
rect 25774 12900 25780 12912
rect 25446 12872 25780 12900
rect 25446 12869 25458 12872
rect 25400 12863 25458 12869
rect 25774 12860 25780 12872
rect 25832 12860 25838 12912
rect 26620 12900 26648 12928
rect 26620 12872 27936 12900
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23860 12804 23949 12832
rect 23431 12801 23443 12804
rect 23385 12795 23443 12801
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 27908 12841 27936 12872
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 24360 12804 24869 12832
rect 24360 12792 24366 12804
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 27893 12835 27951 12841
rect 26651 12804 27108 12832
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 27080 12776 27108 12804
rect 27893 12801 27905 12835
rect 27939 12801 27951 12835
rect 27893 12795 27951 12801
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 15841 12699 15899 12705
rect 15841 12665 15853 12699
rect 15887 12696 15899 12699
rect 16868 12696 16896 12727
rect 15887 12668 16896 12696
rect 15887 12665 15899 12668
rect 15841 12659 15899 12665
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18524 12696 18552 12727
rect 19242 12724 19248 12776
rect 19300 12724 19306 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12733 19855 12767
rect 19797 12727 19855 12733
rect 18196 12668 18552 12696
rect 18969 12699 19027 12705
rect 18196 12656 18202 12668
rect 18969 12665 18981 12699
rect 19015 12696 19027 12699
rect 19429 12699 19487 12705
rect 19429 12696 19441 12699
rect 19015 12668 19441 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 19429 12665 19441 12668
rect 19475 12696 19487 12699
rect 19812 12696 19840 12727
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 20714 12724 20720 12776
rect 20772 12724 20778 12776
rect 24121 12767 24179 12773
rect 20824 12736 24072 12764
rect 20824 12696 20852 12736
rect 19475 12668 19840 12696
rect 20364 12668 20852 12696
rect 19475 12665 19487 12668
rect 19429 12659 19487 12665
rect 13964 12600 14688 12628
rect 17773 12631 17831 12637
rect 13964 12588 13970 12600
rect 17773 12597 17785 12631
rect 17819 12628 17831 12631
rect 17954 12628 17960 12640
rect 17819 12600 17960 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18230 12588 18236 12640
rect 18288 12628 18294 12640
rect 20364 12628 20392 12668
rect 23658 12656 23664 12708
rect 23716 12656 23722 12708
rect 23934 12656 23940 12708
rect 23992 12656 23998 12708
rect 18288 12600 20392 12628
rect 20441 12631 20499 12637
rect 18288 12588 18294 12600
rect 20441 12597 20453 12631
rect 20487 12628 20499 12631
rect 20806 12628 20812 12640
rect 20487 12600 20812 12628
rect 20487 12597 20499 12600
rect 20441 12591 20499 12597
rect 20806 12588 20812 12600
rect 20864 12628 20870 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20864 12600 20913 12628
rect 20864 12588 20870 12600
rect 20901 12597 20913 12600
rect 20947 12597 20959 12631
rect 20901 12591 20959 12597
rect 21818 12588 21824 12640
rect 21876 12588 21882 12640
rect 22094 12588 22100 12640
rect 22152 12588 22158 12640
rect 22925 12631 22983 12637
rect 22925 12597 22937 12631
rect 22971 12628 22983 12631
rect 23952 12628 23980 12656
rect 22971 12600 23980 12628
rect 24044 12628 24072 12736
rect 24121 12733 24133 12767
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 24136 12696 24164 12727
rect 24946 12724 24952 12776
rect 25004 12764 25010 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 25004 12736 25145 12764
rect 25004 12724 25010 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 27062 12724 27068 12776
rect 27120 12724 27126 12776
rect 27706 12724 27712 12776
rect 27764 12724 27770 12776
rect 24673 12699 24731 12705
rect 24673 12696 24685 12699
rect 24136 12668 24685 12696
rect 24673 12665 24685 12668
rect 24719 12665 24731 12699
rect 24673 12659 24731 12665
rect 26234 12656 26240 12708
rect 26292 12696 26298 12708
rect 26513 12699 26571 12705
rect 26513 12696 26525 12699
rect 26292 12668 26525 12696
rect 26292 12656 26298 12668
rect 26513 12665 26525 12668
rect 26559 12696 26571 12699
rect 26559 12668 27476 12696
rect 26559 12665 26571 12668
rect 26513 12659 26571 12665
rect 27448 12640 27476 12668
rect 24762 12628 24768 12640
rect 24044 12600 24768 12628
rect 22971 12597 22983 12600
rect 22925 12591 22983 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 26694 12588 26700 12640
rect 26752 12588 26758 12640
rect 27430 12588 27436 12640
rect 27488 12588 27494 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 3050 12424 3056 12436
rect 2823 12396 3056 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 5169 12427 5227 12433
rect 3804 12396 4936 12424
rect 3804 12356 3832 12396
rect 2516 12328 3832 12356
rect 4908 12356 4936 12396
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5350 12424 5356 12436
rect 5215 12396 5356 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5350 12384 5356 12396
rect 5408 12424 5414 12436
rect 6089 12427 6147 12433
rect 5408 12396 6040 12424
rect 5408 12384 5414 12396
rect 4908 12328 5396 12356
rect 2516 12300 2544 12328
rect 2498 12248 2504 12300
rect 2556 12248 2562 12300
rect 2746 12260 3832 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 2746 12220 2774 12260
rect 1452 12192 2774 12220
rect 2961 12223 3019 12229
rect 1452 12180 1458 12192
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3418 12220 3424 12232
rect 3007 12192 3424 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12220 3571 12223
rect 3694 12220 3700 12232
rect 3559 12192 3700 12220
rect 3559 12189 3571 12192
rect 3513 12183 3571 12189
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 3804 12229 3832 12260
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 4798 12220 4804 12232
rect 3835 12192 4804 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 4798 12180 4804 12192
rect 4856 12220 4862 12232
rect 5258 12220 5264 12232
rect 4856 12192 5264 12220
rect 4856 12180 4862 12192
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 5368 12229 5396 12328
rect 6012 12288 6040 12396
rect 6089 12393 6101 12427
rect 6135 12424 6147 12427
rect 6822 12424 6828 12436
rect 6135 12396 6828 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 8628 12396 9321 12424
rect 8628 12384 8634 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 9692 12396 11008 12424
rect 6457 12359 6515 12365
rect 6457 12325 6469 12359
rect 6503 12325 6515 12359
rect 6457 12319 6515 12325
rect 7561 12359 7619 12365
rect 7561 12325 7573 12359
rect 7607 12325 7619 12359
rect 7561 12319 7619 12325
rect 6472 12288 6500 12319
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6012 12260 6316 12288
rect 6472 12260 6929 12288
rect 6288 12229 6316 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 7576 12288 7604 12319
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 9692 12356 9720 12396
rect 7800 12328 9720 12356
rect 10980 12356 11008 12396
rect 11054 12384 11060 12436
rect 11112 12384 11118 12436
rect 11698 12424 11704 12436
rect 11164 12396 11704 12424
rect 11164 12356 11192 12396
rect 11698 12384 11704 12396
rect 11756 12424 11762 12436
rect 12342 12424 12348 12436
rect 11756 12396 12348 12424
rect 11756 12384 11762 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 12802 12384 12808 12436
rect 12860 12384 12866 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 15289 12427 15347 12433
rect 13044 12396 14964 12424
rect 13044 12384 13050 12396
rect 10980 12328 11192 12356
rect 7800 12316 7806 12328
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7576 12260 8309 12288
rect 6917 12251 6975 12257
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 6273 12223 6331 12229
rect 5399 12192 6224 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 1664 12155 1722 12161
rect 1664 12121 1676 12155
rect 1710 12152 1722 12155
rect 4056 12155 4114 12161
rect 1710 12124 2774 12152
rect 1710 12121 1722 12124
rect 1664 12115 1722 12121
rect 2746 12084 2774 12124
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4706 12152 4712 12164
rect 4102 12124 4712 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 4816 12124 6009 12152
rect 4816 12084 4844 12124
rect 5997 12121 6009 12124
rect 6043 12121 6055 12155
rect 5997 12115 6055 12121
rect 2746 12056 4844 12084
rect 6196 12084 6224 12192
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 6822 12220 6828 12232
rect 6779 12192 6828 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8404 12220 8432 12328
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11296 12328 13308 12356
rect 11296 12316 11302 12328
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12288 8999 12291
rect 9030 12288 9036 12300
rect 8987 12260 9036 12288
rect 8987 12257 8999 12260
rect 8941 12251 8999 12257
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12288 11943 12291
rect 12802 12288 12808 12300
rect 11931 12260 12808 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 8159 12192 8432 12220
rect 9125 12223 9183 12229
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 9766 12220 9772 12232
rect 9723 12192 9772 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 7852 12152 7880 12183
rect 6420 12124 7880 12152
rect 7929 12155 7987 12161
rect 6420 12112 6426 12124
rect 7929 12121 7941 12155
rect 7975 12152 7987 12155
rect 9140 12152 9168 12183
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 9950 12229 9956 12232
rect 9944 12183 9956 12229
rect 9950 12180 9956 12183
rect 10008 12180 10014 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 10744 12192 11437 12220
rect 10744 12180 10750 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 11974 12220 11980 12232
rect 11747 12192 11980 12220
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 11716 12152 11744 12183
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 13280 12229 13308 12328
rect 14090 12316 14096 12368
rect 14148 12316 14154 12368
rect 14108 12288 14136 12316
rect 14461 12291 14519 12297
rect 14108 12260 14412 12288
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12360 12192 12449 12220
rect 7975 12124 9168 12152
rect 11072 12124 11744 12152
rect 7975 12121 7987 12124
rect 7929 12115 7987 12121
rect 6914 12084 6920 12096
rect 6196 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 11072 12084 11100 12124
rect 8168 12056 11100 12084
rect 8168 12044 8174 12056
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12360 12093 12388 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 12216 12056 12357 12084
rect 12216 12044 12222 12056
rect 12345 12053 12357 12056
rect 12391 12053 12403 12087
rect 12345 12047 12403 12053
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12636 12084 12664 12183
rect 12492 12056 12664 12084
rect 13280 12084 13308 12183
rect 13446 12180 13452 12232
rect 13504 12180 13510 12232
rect 13538 12180 13544 12232
rect 13596 12220 13602 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13596 12192 14105 12220
rect 13596 12180 13602 12192
rect 14093 12189 14105 12192
rect 14139 12220 14151 12223
rect 14274 12220 14280 12232
rect 14139 12192 14280 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14384 12229 14412 12260
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14507 12260 14841 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 14936 12288 14964 12396
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 16758 12424 16764 12436
rect 15335 12396 16764 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17773 12427 17831 12433
rect 17773 12393 17785 12427
rect 17819 12424 17831 12427
rect 18138 12424 18144 12436
rect 17819 12396 18144 12424
rect 17819 12393 17831 12396
rect 17773 12387 17831 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18785 12427 18843 12433
rect 18785 12393 18797 12427
rect 18831 12424 18843 12427
rect 19242 12424 19248 12436
rect 18831 12396 19248 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 19978 12424 19984 12436
rect 19659 12396 19984 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20714 12424 20720 12436
rect 20119 12396 20720 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 22094 12424 22100 12436
rect 21008 12396 22100 12424
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16485 12359 16543 12365
rect 16485 12356 16497 12359
rect 16071 12328 16497 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16485 12325 16497 12328
rect 16531 12356 16543 12359
rect 16666 12356 16672 12368
rect 16531 12328 16672 12356
rect 16531 12325 16543 12328
rect 16485 12319 16543 12325
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 14936 12260 16129 12288
rect 14829 12251 14887 12257
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 18782 12248 18788 12300
rect 18840 12288 18846 12300
rect 18840 12260 19564 12288
rect 18840 12248 18846 12260
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 13909 12155 13967 12161
rect 13909 12121 13921 12155
rect 13955 12152 13967 12155
rect 14458 12152 14464 12164
rect 13955 12124 14464 12152
rect 13955 12121 13967 12124
rect 13909 12115 13967 12121
rect 14458 12112 14464 12124
rect 14516 12152 14522 12164
rect 14660 12152 14688 12183
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15344 12192 15393 12220
rect 15344 12180 15350 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 16264 12192 16313 12220
rect 16264 12180 16270 12192
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 17954 12180 17960 12232
rect 18012 12180 18018 12232
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 19536 12229 19564 12260
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 21008 12297 21036 12396
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 23845 12427 23903 12433
rect 23845 12393 23857 12427
rect 23891 12424 23903 12427
rect 24302 12424 24308 12436
rect 23891 12396 24308 12424
rect 23891 12393 23903 12396
rect 23845 12387 23903 12393
rect 24302 12384 24308 12396
rect 24360 12384 24366 12436
rect 25041 12427 25099 12433
rect 25041 12393 25053 12427
rect 25087 12424 25099 12427
rect 26326 12424 26332 12436
rect 25087 12396 26332 12424
rect 25087 12393 25099 12396
rect 25041 12387 25099 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 21358 12316 21364 12368
rect 21416 12316 21422 12368
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 25317 12359 25375 12365
rect 21508 12328 22876 12356
rect 21508 12316 21514 12328
rect 20993 12291 21051 12297
rect 20993 12257 21005 12291
rect 21039 12257 21051 12291
rect 21376 12288 21404 12316
rect 21729 12291 21787 12297
rect 21729 12288 21741 12291
rect 21376 12260 21741 12288
rect 20993 12251 21051 12257
rect 21729 12257 21741 12260
rect 21775 12257 21787 12291
rect 21729 12251 21787 12257
rect 22848 12229 22876 12328
rect 25317 12325 25329 12359
rect 25363 12356 25375 12359
rect 25363 12328 27936 12356
rect 25363 12325 25375 12328
rect 25317 12319 25375 12325
rect 24118 12288 24124 12300
rect 23584 12260 24124 12288
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18104 12192 18705 12220
rect 18104 12180 18110 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19567 12192 19993 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 20272 12152 20300 12183
rect 23290 12180 23296 12232
rect 23348 12180 23354 12232
rect 23584 12229 23612 12260
rect 24118 12248 24124 12260
rect 24176 12288 24182 12300
rect 24176 12260 24808 12288
rect 24176 12248 24182 12260
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 24026 12180 24032 12232
rect 24084 12180 24090 12232
rect 24780 12229 24808 12260
rect 25590 12248 25596 12300
rect 25648 12248 25654 12300
rect 25777 12291 25835 12297
rect 25777 12257 25789 12291
rect 25823 12288 25835 12291
rect 26694 12288 26700 12300
rect 25823 12260 26700 12288
rect 25823 12257 25835 12260
rect 25777 12251 25835 12257
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 26786 12248 26792 12300
rect 26844 12248 26850 12300
rect 27706 12248 27712 12300
rect 27764 12248 27770 12300
rect 27908 12297 27936 12328
rect 27982 12316 27988 12368
rect 28040 12356 28046 12368
rect 28077 12359 28135 12365
rect 28077 12356 28089 12359
rect 28040 12328 28089 12356
rect 28040 12316 28046 12328
rect 28077 12325 28089 12328
rect 28123 12325 28135 12359
rect 28077 12319 28135 12325
rect 27893 12291 27951 12297
rect 27893 12257 27905 12291
rect 27939 12257 27951 12291
rect 27893 12251 27951 12257
rect 24489 12223 24547 12229
rect 24489 12189 24501 12223
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 14516 12124 14688 12152
rect 19812 12124 20300 12152
rect 21821 12155 21879 12161
rect 14516 12112 14522 12124
rect 14090 12084 14096 12096
rect 13280 12056 14096 12084
rect 12492 12044 12498 12056
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14182 12044 14188 12096
rect 14240 12044 14246 12096
rect 19812 12093 19840 12124
rect 21821 12121 21833 12155
rect 21867 12152 21879 12155
rect 21867 12124 22094 12152
rect 21867 12121 21879 12124
rect 21821 12115 21879 12121
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12053 19855 12087
rect 22066 12084 22094 12124
rect 22738 12112 22744 12164
rect 22796 12112 22802 12164
rect 24504 12152 24532 12183
rect 25130 12152 25136 12164
rect 24504 12124 25136 12152
rect 25130 12112 25136 12124
rect 25188 12112 25194 12164
rect 25240 12152 25268 12183
rect 25498 12180 25504 12232
rect 25556 12180 25562 12232
rect 26234 12152 26240 12164
rect 25240 12124 26240 12152
rect 26234 12112 26240 12124
rect 26292 12112 26298 12164
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 22066 12056 23029 12084
rect 19797 12047 19855 12053
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 23017 12047 23075 12053
rect 23385 12087 23443 12093
rect 23385 12053 23397 12087
rect 23431 12084 23443 12087
rect 23566 12084 23572 12096
rect 23431 12056 23572 12084
rect 23431 12053 23443 12056
rect 23385 12047 23443 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 24302 12084 24308 12096
rect 23707 12056 24308 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24486 12044 24492 12096
rect 24544 12084 24550 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 24544 12056 24593 12084
rect 24544 12044 24550 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 24857 12087 24915 12093
rect 24857 12053 24869 12087
rect 24903 12084 24915 12087
rect 25958 12084 25964 12096
rect 24903 12056 25964 12084
rect 24903 12053 24915 12056
rect 24857 12047 24915 12053
rect 25958 12044 25964 12056
rect 26016 12044 26022 12096
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 4706 11840 4712 11892
rect 4764 11840 4770 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5166 11880 5172 11892
rect 5040 11852 5172 11880
rect 5040 11840 5046 11852
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7006 11840 7012 11892
rect 7064 11840 7070 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7742 11880 7748 11892
rect 7147 11852 7748 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10042 11880 10048 11892
rect 9732 11852 10048 11880
rect 9732 11840 9738 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10686 11840 10692 11892
rect 10744 11840 10750 11892
rect 12158 11840 12164 11892
rect 12216 11840 12222 11892
rect 12434 11840 12440 11892
rect 12492 11840 12498 11892
rect 12802 11840 12808 11892
rect 12860 11840 12866 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 2038 11772 2044 11824
rect 2096 11772 2102 11824
rect 4614 11812 4620 11824
rect 3068 11784 4620 11812
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1627 11648 1961 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2958 11636 2964 11688
rect 3016 11636 3022 11688
rect 3068 11685 3096 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7024 11812 7052 11840
rect 13096 11812 13124 11843
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13504 11852 13553 11880
rect 13504 11840 13510 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 14274 11840 14280 11892
rect 14332 11840 14338 11892
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 14516 11852 14749 11880
rect 14516 11840 14522 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 14737 11843 14795 11849
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15620 11852 15853 11880
rect 15620 11840 15626 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 15841 11843 15899 11849
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16206 11880 16212 11892
rect 16071 11852 16212 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11849 16359 11883
rect 16301 11843 16359 11849
rect 7024 11784 12940 11812
rect 13096 11784 13768 11812
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3476 11716 3985 11744
rect 3476 11704 3482 11716
rect 3973 11713 3985 11716
rect 4019 11744 4031 11747
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 4019 11716 4077 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 5068 11747 5126 11753
rect 5068 11713 5080 11747
rect 5114 11744 5126 11747
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 5114 11716 7021 11744
rect 5114 11713 5126 11716
rect 5068 11707 5126 11713
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11645 3111 11679
rect 3053 11639 3111 11645
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 3252 11608 3280 11639
rect 2648 11580 3280 11608
rect 2648 11568 2654 11580
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 3786 11500 3792 11552
rect 3844 11500 3850 11552
rect 4080 11540 4108 11707
rect 4798 11636 4804 11688
rect 4856 11636 4862 11688
rect 6362 11636 6368 11688
rect 6420 11636 6426 11688
rect 7300 11608 7328 11707
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 7944 11753 7972 11784
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7760 11676 7788 11707
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8536 11716 8677 11744
rect 8536 11704 8542 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 10870 11744 10876 11756
rect 9723 11716 10876 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11296 11716 11713 11744
rect 11296 11704 11302 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 12802 11744 12808 11756
rect 12759 11716 12808 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 7432 11648 9996 11676
rect 7432 11636 7438 11648
rect 8294 11608 8300 11620
rect 6196 11580 7328 11608
rect 7484 11580 8300 11608
rect 5442 11540 5448 11552
rect 4080 11512 5448 11540
rect 5442 11500 5448 11512
rect 5500 11540 5506 11552
rect 6196 11549 6224 11580
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 5500 11512 6193 11540
rect 5500 11500 5506 11512
rect 6181 11509 6193 11512
rect 6227 11509 6239 11543
rect 6181 11503 6239 11509
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 7484 11540 7512 11580
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 6328 11512 7512 11540
rect 6328 11500 6334 11512
rect 7558 11500 7564 11552
rect 7616 11500 7622 11552
rect 7834 11500 7840 11552
rect 7892 11500 7898 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 9858 11540 9864 11552
rect 8803 11512 9864 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 9968 11540 9996 11648
rect 10042 11636 10048 11688
rect 10100 11636 10106 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11112 11648 11529 11676
rect 11112 11636 11118 11648
rect 11517 11645 11529 11648
rect 11563 11676 11575 11679
rect 12066 11676 12072 11688
rect 11563 11648 12072 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 10060 11608 10088 11636
rect 12728 11608 12756 11707
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 10060 11580 12756 11608
rect 12912 11608 12940 11784
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 13136 11716 13277 11744
rect 13136 11704 13142 11716
rect 13265 11713 13277 11716
rect 13311 11744 13323 11747
rect 13538 11744 13544 11756
rect 13311 11716 13544 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13740 11753 13768 11784
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 14200 11744 14228 11840
rect 14292 11812 14320 11840
rect 14292 11784 15792 11812
rect 15764 11753 15792 11784
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14200 11716 14289 11744
rect 13725 11707 13783 11713
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16316 11744 16344 11843
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 24397 11883 24455 11889
rect 17092 11852 20208 11880
rect 17092 11840 17098 11852
rect 19518 11812 19524 11824
rect 16592 11784 19524 11812
rect 16255 11716 16344 11744
rect 16485 11747 16543 11753
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16485 11713 16497 11747
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11676 14151 11679
rect 14458 11676 14464 11688
rect 14139 11648 14464 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 15764 11676 15792 11707
rect 16500 11676 16528 11707
rect 15764 11648 16528 11676
rect 16592 11608 16620 11784
rect 18708 11753 18736 11784
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 20180 11753 20208 11852
rect 24397 11849 24409 11883
rect 24443 11880 24455 11883
rect 26053 11883 26111 11889
rect 24443 11852 24900 11880
rect 24443 11849 24455 11852
rect 24397 11843 24455 11849
rect 20524 11815 20582 11821
rect 20524 11781 20536 11815
rect 20570 11812 20582 11815
rect 21266 11812 21272 11824
rect 20570 11784 21272 11812
rect 20570 11781 20582 11784
rect 20524 11775 20582 11781
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 21634 11772 21640 11824
rect 21692 11812 21698 11824
rect 21913 11815 21971 11821
rect 21913 11812 21925 11815
rect 21692 11784 21925 11812
rect 21692 11772 21698 11784
rect 21913 11781 21925 11784
rect 21959 11781 21971 11815
rect 21913 11775 21971 11781
rect 22002 11772 22008 11824
rect 22060 11772 22066 11824
rect 23290 11772 23296 11824
rect 23348 11772 23354 11824
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11744 23259 11747
rect 23308 11744 23336 11772
rect 23247 11716 23336 11744
rect 23477 11747 23535 11753
rect 23247 11713 23259 11716
rect 23201 11707 23259 11713
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 24026 11744 24032 11756
rect 23523 11716 24032 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 12912 11580 16620 11608
rect 18524 11676 18552 11707
rect 24026 11704 24032 11716
rect 24084 11704 24090 11756
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11713 24639 11747
rect 24872 11744 24900 11852
rect 26053 11849 26065 11883
rect 26099 11880 26111 11883
rect 27062 11880 27068 11892
rect 26099 11852 27068 11880
rect 26099 11849 26111 11852
rect 26053 11843 26111 11849
rect 27062 11840 27068 11852
rect 27120 11880 27126 11892
rect 27120 11852 27200 11880
rect 27120 11840 27126 11852
rect 24940 11815 24998 11821
rect 24940 11781 24952 11815
rect 24986 11812 24998 11815
rect 26418 11812 26424 11824
rect 24986 11784 26424 11812
rect 24986 11781 24998 11784
rect 24940 11775 24998 11781
rect 26418 11772 26424 11784
rect 26476 11772 26482 11824
rect 26970 11744 26976 11756
rect 24872 11716 26976 11744
rect 24581 11707 24639 11713
rect 19058 11676 19064 11688
rect 18524 11648 19064 11676
rect 18524 11540 18552 11648
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 20254 11636 20260 11688
rect 20312 11636 20318 11688
rect 22738 11636 22744 11688
rect 22796 11636 22802 11688
rect 23658 11636 23664 11688
rect 23716 11636 23722 11688
rect 23750 11636 23756 11688
rect 23808 11676 23814 11688
rect 24596 11676 24624 11707
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 27172 11753 27200 11852
rect 28166 11840 28172 11892
rect 28224 11840 28230 11892
rect 28353 11883 28411 11889
rect 28353 11849 28365 11883
rect 28399 11880 28411 11883
rect 28442 11880 28448 11892
rect 28399 11852 28448 11880
rect 28399 11849 28411 11852
rect 28353 11843 28411 11849
rect 28442 11840 28448 11852
rect 28500 11840 28506 11892
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27430 11704 27436 11756
rect 27488 11704 27494 11756
rect 27525 11747 27583 11753
rect 27525 11713 27537 11747
rect 27571 11744 27583 11747
rect 27982 11744 27988 11756
rect 27571 11716 27988 11744
rect 27571 11713 27583 11716
rect 27525 11707 27583 11713
rect 27982 11704 27988 11716
rect 28040 11704 28046 11756
rect 28261 11747 28319 11753
rect 28261 11713 28273 11747
rect 28307 11744 28319 11747
rect 28534 11744 28540 11756
rect 28307 11716 28540 11744
rect 28307 11713 28319 11716
rect 28261 11707 28319 11713
rect 28534 11704 28540 11716
rect 28592 11704 28598 11756
rect 23808 11648 24624 11676
rect 24673 11679 24731 11685
rect 23808 11636 23814 11648
rect 24673 11645 24685 11679
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 26237 11679 26295 11685
rect 26237 11645 26249 11679
rect 26283 11676 26295 11679
rect 26283 11648 26648 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 19981 11611 20039 11617
rect 19981 11577 19993 11611
rect 20027 11577 20039 11611
rect 23474 11608 23480 11620
rect 19981 11571 20039 11577
rect 21192 11580 23480 11608
rect 9968 11512 18552 11540
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18690 11540 18696 11552
rect 18647 11512 18696 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 19996 11540 20024 11571
rect 21192 11540 21220 11580
rect 23474 11568 23480 11580
rect 23532 11568 23538 11620
rect 19996 11512 21220 11540
rect 21634 11500 21640 11552
rect 21692 11500 21698 11552
rect 23014 11500 23020 11552
rect 23072 11500 23078 11552
rect 24118 11500 24124 11552
rect 24176 11500 24182 11552
rect 24688 11540 24716 11639
rect 26620 11552 26648 11648
rect 27338 11636 27344 11688
rect 27396 11676 27402 11688
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 27396 11648 27721 11676
rect 27396 11636 27402 11648
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 26973 11611 27031 11617
rect 26973 11577 26985 11611
rect 27019 11608 27031 11611
rect 27019 11580 27384 11608
rect 27019 11577 27031 11580
rect 26973 11571 27031 11577
rect 24854 11540 24860 11552
rect 24688 11512 24860 11540
rect 24854 11500 24860 11512
rect 24912 11500 24918 11552
rect 26602 11500 26608 11552
rect 26660 11500 26666 11552
rect 26786 11500 26792 11552
rect 26844 11500 26850 11552
rect 27246 11500 27252 11552
rect 27304 11500 27310 11552
rect 27356 11540 27384 11580
rect 28074 11540 28080 11552
rect 27356 11512 28080 11540
rect 28074 11500 28080 11512
rect 28132 11500 28138 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 2038 11296 2044 11348
rect 2096 11296 2102 11348
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11305 2743 11339
rect 2685 11299 2743 11305
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 6638 11336 6644 11348
rect 5491 11308 6644 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 2133 11271 2191 11277
rect 2133 11237 2145 11271
rect 2179 11237 2191 11271
rect 2133 11231 2191 11237
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2148 11132 2176 11231
rect 2498 11200 2504 11212
rect 2332 11172 2504 11200
rect 2332 11141 2360 11172
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 2700 11200 2728 11299
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 6788 11308 7512 11336
rect 6788 11296 6794 11308
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 4706 11268 4712 11280
rect 3651 11240 4712 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 5169 11271 5227 11277
rect 5169 11237 5181 11271
rect 5215 11268 5227 11271
rect 5534 11268 5540 11280
rect 5215 11240 5540 11268
rect 5215 11237 5227 11240
rect 5169 11231 5227 11237
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 7484 11268 7512 11308
rect 8128 11308 9413 11336
rect 8128 11268 8156 11308
rect 9401 11305 9413 11308
rect 9447 11336 9459 11339
rect 10134 11336 10140 11348
rect 9447 11308 10140 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 11882 11336 11888 11348
rect 11563 11308 11888 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 11882 11296 11888 11308
rect 11940 11336 11946 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11940 11308 11989 11336
rect 11940 11296 11946 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 19352 11308 20760 11336
rect 7484 11240 8156 11268
rect 8297 11271 8355 11277
rect 8297 11237 8309 11271
rect 8343 11237 8355 11271
rect 8297 11231 8355 11237
rect 8573 11271 8631 11277
rect 8573 11237 8585 11271
rect 8619 11268 8631 11271
rect 9861 11271 9919 11277
rect 8619 11240 9260 11268
rect 8619 11237 8631 11240
rect 8573 11231 8631 11237
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 2700 11172 3157 11200
rect 3145 11169 3157 11172
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 3418 11160 3424 11212
rect 3476 11160 3482 11212
rect 3786 11160 3792 11212
rect 3844 11160 3850 11212
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4203 11172 4537 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 6730 11200 6736 11212
rect 4525 11163 4583 11169
rect 5276 11172 6736 11200
rect 1903 11104 2176 11132
rect 2317 11135 2375 11141
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2317 11101 2329 11135
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2682 11132 2688 11144
rect 2464 11104 2688 11132
rect 2464 11092 2470 11104
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3436 11132 3464 11160
rect 3016 11104 3464 11132
rect 3804 11132 3832 11160
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3804 11104 3985 11132
rect 3016 11092 3022 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4080 11064 4108 11095
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 5276 11132 5304 11172
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 7834 11160 7840 11212
rect 7892 11160 7898 11212
rect 8312 11200 8340 11231
rect 9232 11209 9260 11240
rect 9861 11237 9873 11271
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 10321 11271 10379 11277
rect 10321 11237 10333 11271
rect 10367 11268 10379 11271
rect 14458 11268 14464 11280
rect 10367 11240 11836 11268
rect 10367 11237 10379 11240
rect 10321 11231 10379 11237
rect 9033 11203 9091 11209
rect 8312 11172 8800 11200
rect 4387 11104 5304 11132
rect 5353 11135 5411 11141
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5442 11132 5448 11144
rect 5399 11104 5448 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5442 11092 5448 11104
rect 5500 11132 5506 11144
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 5500 11104 5641 11132
rect 5500 11092 5506 11104
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 7558 11092 7564 11144
rect 7616 11092 7622 11144
rect 4264 11064 4292 11092
rect 7852 11064 7880 11160
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 8772 11141 8800 11172
rect 9033 11169 9045 11203
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11169 9275 11203
rect 9876 11200 9904 11231
rect 9876 11172 10548 11200
rect 9217 11163 9275 11169
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11101 8815 11135
rect 9048 11132 9076 11163
rect 9582 11132 9588 11144
rect 9048 11104 9588 11132
rect 8757 11095 8815 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10520 11141 10548 11172
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11808 11209 11836 11240
rect 11900 11240 14464 11268
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11204 11172 11621 11200
rect 11204 11160 11210 11172
rect 11609 11169 11621 11172
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10836 11104 10885 11132
rect 10836 11092 10842 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 2746 11036 4108 11064
rect 4172 11036 4292 11064
rect 7222 11036 7880 11064
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 2746 10996 2774 11036
rect 2648 10968 2774 10996
rect 3789 10999 3847 11005
rect 2648 10956 2654 10968
rect 3789 10965 3801 10999
rect 3835 10996 3847 10999
rect 4172 10996 4200 11036
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 10888 11064 10916 11095
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 11020 11104 11069 11132
rect 11020 11092 11026 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11900 11064 11928 11240
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 14737 11271 14795 11277
rect 14737 11268 14749 11271
rect 14700 11240 14749 11268
rect 14700 11228 14706 11240
rect 14737 11237 14749 11240
rect 14783 11237 14795 11271
rect 14737 11231 14795 11237
rect 17310 11200 17316 11212
rect 12544 11172 15332 11200
rect 12544 11141 12572 11172
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 12544 11064 12572 11095
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12676 11104 12817 11132
rect 12676 11092 12682 11104
rect 12805 11101 12817 11104
rect 12851 11132 12863 11135
rect 13170 11132 13176 11144
rect 12851 11104 13176 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14148 11104 14381 11132
rect 14148 11092 14154 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 8444 11036 10824 11064
rect 10888 11036 11928 11064
rect 11983 11036 12572 11064
rect 14384 11064 14412 11095
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 15304 11141 15332 11172
rect 15396 11172 17316 11200
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15396 11064 15424 11172
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17494 11160 17500 11212
rect 17552 11160 17558 11212
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 17678 11092 17684 11144
rect 17736 11092 17742 11144
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 19352 11141 19380 11308
rect 20732 11268 20760 11308
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20956 11308 21005 11336
rect 20956 11296 20962 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 22060 11308 22661 11336
rect 22060 11296 22066 11308
rect 22649 11305 22661 11308
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 23017 11339 23075 11345
rect 23017 11305 23029 11339
rect 23063 11336 23075 11339
rect 23658 11336 23664 11348
rect 23063 11308 23664 11336
rect 23063 11305 23075 11308
rect 23017 11299 23075 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24118 11296 24124 11348
rect 24176 11296 24182 11348
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 26881 11339 26939 11345
rect 26881 11336 26893 11339
rect 25648 11308 26893 11336
rect 25648 11296 25654 11308
rect 26881 11305 26893 11308
rect 26927 11305 26939 11339
rect 26881 11299 26939 11305
rect 26988 11308 28304 11336
rect 24394 11268 24400 11280
rect 20732 11240 24400 11268
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 26602 11228 26608 11280
rect 26660 11268 26666 11280
rect 26988 11268 27016 11308
rect 26660 11240 27016 11268
rect 26660 11228 26666 11240
rect 28276 11212 28304 11308
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11169 19671 11203
rect 24854 11200 24860 11212
rect 19613 11163 19671 11169
rect 20824 11172 24860 11200
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17828 11104 18245 11132
rect 17828 11092 17834 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11101 19395 11135
rect 19628 11132 19656 11163
rect 20824 11132 20852 11172
rect 24854 11160 24860 11172
rect 24912 11200 24918 11212
rect 25225 11203 25283 11209
rect 25225 11200 25237 11203
rect 24912 11172 25237 11200
rect 24912 11160 24918 11172
rect 25225 11169 25237 11172
rect 25271 11169 25283 11203
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 25225 11163 25283 11169
rect 26252 11172 27169 11200
rect 19628 11104 20852 11132
rect 19337 11095 19395 11101
rect 14384 11036 15424 11064
rect 15565 11067 15623 11073
rect 8444 11024 8450 11036
rect 3835 10968 4200 10996
rect 3835 10965 3847 10968
rect 3789 10959 3847 10965
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 7098 10996 7104 11008
rect 4304 10968 7104 10996
rect 4304 10956 4310 10968
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7616 10968 7757 10996
rect 7616 10956 7622 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 10796 10996 10824 11036
rect 11983 10996 12011 11036
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 15654 11064 15660 11076
rect 15611 11036 15660 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 18892 11064 18920 11095
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20956 11104 21097 11132
rect 20956 11092 20962 11104
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21634 11092 21640 11144
rect 21692 11132 21698 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21692 11104 21833 11132
rect 21692 11092 21698 11104
rect 21821 11101 21833 11104
rect 21867 11132 21879 11135
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 21867 11104 22569 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23201 11135 23259 11141
rect 23201 11132 23213 11135
rect 23072 11104 23213 11132
rect 23072 11092 23078 11104
rect 23201 11101 23213 11104
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23477 11135 23535 11141
rect 23477 11101 23489 11135
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 17144 11036 18920 11064
rect 19880 11067 19938 11073
rect 17144 11008 17172 11036
rect 19880 11033 19892 11067
rect 19926 11064 19938 11067
rect 22465 11067 22523 11073
rect 22465 11064 22477 11067
rect 19926 11036 22477 11064
rect 19926 11033 19938 11036
rect 19880 11027 19938 11033
rect 22465 11033 22477 11036
rect 22511 11033 22523 11067
rect 23492 11064 23520 11095
rect 23566 11092 23572 11144
rect 23624 11132 23630 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23624 11104 23673 11132
rect 23624 11092 23630 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24176 11104 24409 11132
rect 24176 11092 24182 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24486 11092 24492 11144
rect 24544 11132 24550 11144
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24544 11104 24593 11132
rect 24544 11092 24550 11104
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 25240 11132 25268 11163
rect 26252 11132 26280 11172
rect 27157 11169 27169 11172
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 28258 11160 28264 11212
rect 28316 11160 28322 11212
rect 25240 11104 26280 11132
rect 26878 11092 26884 11144
rect 26936 11132 26942 11144
rect 27065 11135 27123 11141
rect 27065 11132 27077 11135
rect 26936 11104 27077 11132
rect 26936 11092 26942 11104
rect 27065 11101 27077 11104
rect 27111 11101 27123 11135
rect 27065 11095 27123 11101
rect 27424 11135 27482 11141
rect 27424 11101 27436 11135
rect 27470 11132 27482 11135
rect 28166 11132 28172 11144
rect 27470 11104 28172 11132
rect 27470 11101 27482 11104
rect 27424 11095 27482 11101
rect 28166 11092 28172 11104
rect 28224 11092 28230 11144
rect 24780 11064 24808 11092
rect 23492 11036 24808 11064
rect 25492 11067 25550 11073
rect 22465 11027 22523 11033
rect 25492 11033 25504 11067
rect 25538 11064 25550 11067
rect 26142 11064 26148 11076
rect 25538 11036 26148 11064
rect 25538 11033 25550 11036
rect 25492 11027 25550 11033
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 10796 10968 12011 10996
rect 7745 10959 7803 10965
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 17126 10956 17132 11008
rect 17184 10956 17190 11008
rect 18138 10956 18144 11008
rect 18196 10956 18202 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 18325 10999 18383 11005
rect 18325 10996 18337 10999
rect 18288 10968 18337 10996
rect 18288 10956 18294 10968
rect 18325 10965 18337 10968
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 18693 10999 18751 11005
rect 18693 10965 18705 10999
rect 18739 10996 18751 10999
rect 18782 10996 18788 11008
rect 18739 10968 18788 10996
rect 18739 10965 18751 10968
rect 18693 10959 18751 10965
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 21729 10999 21787 11005
rect 21729 10996 21741 10999
rect 21140 10968 21741 10996
rect 21140 10956 21146 10968
rect 21729 10965 21741 10968
rect 21775 10965 21787 10999
rect 21729 10959 21787 10965
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 24210 10996 24216 11008
rect 22336 10968 24216 10996
rect 22336 10956 22342 10968
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 25038 10956 25044 11008
rect 25096 10956 25102 11008
rect 27522 10956 27528 11008
rect 27580 10996 27586 11008
rect 28537 10999 28595 11005
rect 28537 10996 28549 10999
rect 27580 10968 28549 10996
rect 27580 10956 27586 10968
rect 28537 10965 28549 10968
rect 28583 10965 28595 10999
rect 28537 10959 28595 10965
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 2958 10792 2964 10804
rect 2639 10764 2964 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 5350 10792 5356 10804
rect 3384 10764 5356 10792
rect 3384 10752 3390 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 5626 10752 5632 10804
rect 5684 10752 5690 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7742 10792 7748 10804
rect 6972 10764 7748 10792
rect 6972 10752 6978 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 10042 10752 10048 10804
rect 10100 10752 10106 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10192 10764 10425 10792
rect 10192 10752 10198 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 10962 10752 10968 10804
rect 11020 10752 11026 10804
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 12802 10792 12808 10804
rect 11563 10764 12808 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13633 10795 13691 10801
rect 13633 10761 13645 10795
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 13909 10795 13967 10801
rect 13909 10761 13921 10795
rect 13955 10792 13967 10795
rect 14550 10792 14556 10804
rect 13955 10764 14556 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 2406 10724 2412 10736
rect 1596 10696 2412 10724
rect 1596 10668 1624 10696
rect 2406 10684 2412 10696
rect 2464 10684 2470 10736
rect 4798 10724 4804 10736
rect 2700 10696 4804 10724
rect 1578 10616 1584 10668
rect 1636 10616 1642 10668
rect 2700 10665 2728 10696
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 2685 10659 2743 10665
rect 1857 10619 1915 10625
rect 1964 10628 2360 10656
rect 1872 10588 1900 10619
rect 1964 10597 1992 10628
rect 1412 10560 1900 10588
rect 1949 10591 2007 10597
rect 1412 10529 1440 10560
rect 1949 10557 1961 10591
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 1397 10523 1455 10529
rect 1397 10489 1409 10523
rect 1443 10489 1455 10523
rect 1397 10483 1455 10489
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 2148 10520 2176 10551
rect 1719 10492 2176 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 2332 10452 2360 10628
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2952 10659 3010 10665
rect 2952 10625 2964 10659
rect 2998 10656 3010 10659
rect 3510 10656 3516 10668
rect 2998 10628 3516 10656
rect 2998 10625 3010 10628
rect 2952 10619 3010 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4172 10665 4200 10696
rect 4798 10684 4804 10696
rect 4856 10724 4862 10736
rect 6104 10724 6132 10752
rect 4856 10696 6132 10724
rect 4856 10684 4862 10696
rect 6362 10684 6368 10736
rect 6420 10684 6426 10736
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 4424 10659 4482 10665
rect 4424 10625 4436 10659
rect 4470 10656 4482 10659
rect 4890 10656 4896 10668
rect 4470 10628 4896 10656
rect 4470 10625 4482 10628
rect 4424 10619 4482 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5258 10656 5264 10668
rect 5040 10628 5264 10656
rect 5040 10616 5046 10628
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5592 10628 5825 10656
rect 5592 10616 5598 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6380 10656 6408 10684
rect 6135 10628 6408 10656
rect 6632 10659 6690 10665
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6632 10625 6644 10659
rect 6678 10656 6690 10659
rect 7190 10656 7196 10668
rect 6678 10628 7196 10656
rect 6678 10625 6690 10628
rect 6632 10619 6690 10625
rect 4264 10588 4292 10616
rect 6104 10588 6132 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9916 10628 9965 10656
rect 9916 10616 9922 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 10060 10656 10088 10752
rect 13357 10727 13415 10733
rect 13357 10724 13369 10727
rect 11256 10696 11836 10724
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10060 10628 10885 10656
rect 9953 10619 10011 10625
rect 10873 10625 10885 10628
rect 10919 10656 10931 10659
rect 11256 10656 11284 10696
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10919 10628 11345 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11701 10659 11759 10665
rect 11333 10619 11391 10625
rect 11440 10654 11652 10656
rect 11701 10654 11713 10659
rect 11440 10628 11713 10654
rect 3988 10560 4292 10588
rect 5552 10560 6132 10588
rect 6365 10591 6423 10597
rect 3988 10452 4016 10560
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 5552 10529 5580 10560
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 5537 10523 5595 10529
rect 5537 10520 5549 10523
rect 5316 10492 5549 10520
rect 5316 10480 5322 10492
rect 5537 10489 5549 10492
rect 5583 10489 5595 10523
rect 5537 10483 5595 10489
rect 6086 10480 6092 10532
rect 6144 10520 6150 10532
rect 6380 10520 6408 10551
rect 7834 10548 7840 10600
rect 7892 10548 7898 10600
rect 8018 10548 8024 10600
rect 8076 10548 8082 10600
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 10778 10588 10784 10600
rect 9815 10560 10784 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 6144 10492 6408 10520
rect 11149 10523 11207 10529
rect 6144 10480 6150 10492
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 11440 10520 11468 10628
rect 11624 10626 11713 10628
rect 11701 10625 11713 10626
rect 11747 10625 11759 10659
rect 11808 10656 11836 10696
rect 11992 10696 13369 10724
rect 11992 10665 12020 10696
rect 13357 10693 13369 10696
rect 13403 10693 13415 10727
rect 13648 10724 13676 10755
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 14700 10764 15117 10792
rect 14700 10752 14706 10764
rect 15105 10761 15117 10764
rect 15151 10761 15163 10795
rect 15105 10755 15163 10761
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 16022 10792 16028 10804
rect 15243 10764 16028 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 18138 10792 18144 10804
rect 17727 10764 18144 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 19518 10752 19524 10804
rect 19576 10752 19582 10804
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 24213 10795 24271 10801
rect 19760 10764 23428 10792
rect 19760 10752 19766 10764
rect 17126 10724 17132 10736
rect 13648 10696 14136 10724
rect 13357 10687 13415 10693
rect 11977 10659 12035 10665
rect 11808 10628 11928 10656
rect 11701 10619 11759 10625
rect 11514 10548 11520 10600
rect 11572 10588 11578 10600
rect 11790 10588 11796 10600
rect 11572 10560 11796 10588
rect 11572 10548 11578 10560
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 11900 10588 11928 10628
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 12986 10656 12992 10668
rect 11977 10619 12035 10625
rect 12084 10628 12992 10656
rect 12084 10588 12112 10628
rect 12986 10616 12992 10628
rect 13044 10656 13050 10668
rect 14108 10665 14136 10696
rect 14200 10696 15424 10724
rect 14200 10665 14228 10696
rect 15396 10668 15424 10696
rect 16960 10696 17132 10724
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 13044 10628 13277 10656
rect 13044 10616 13050 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14323 10628 14657 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 11900 10560 12112 10588
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10588 12587 10591
rect 12618 10588 12624 10600
rect 12575 10560 12624 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 12544 10520 12572 10551
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 12802 10588 12808 10600
rect 12759 10560 12808 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 13832 10588 13860 10619
rect 14200 10588 14228 10619
rect 15378 10616 15384 10668
rect 15436 10616 15442 10668
rect 15838 10616 15844 10668
rect 15896 10616 15902 10668
rect 16960 10665 16988 10696
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 18690 10684 18696 10736
rect 18748 10684 18754 10736
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17773 10659 17831 10665
rect 17083 10628 17724 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 13780 10560 14228 10588
rect 13780 10548 13786 10560
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 15712 10560 17172 10588
rect 15712 10548 15718 10560
rect 11195 10492 11468 10520
rect 12268 10492 12572 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 2332 10424 4016 10452
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4338 10452 4344 10464
rect 4111 10424 4344 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 5902 10412 5908 10464
rect 5960 10412 5966 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 12268 10452 12296 10492
rect 7156 10424 12296 10452
rect 7156 10412 7162 10424
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 12400 10424 12449 10452
rect 12400 10412 12406 10424
rect 12437 10421 12449 10424
rect 12483 10452 12495 10455
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12483 10424 12909 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 16022 10412 16028 10464
rect 16080 10412 16086 10464
rect 16758 10412 16764 10464
rect 16816 10412 16822 10464
rect 17144 10452 17172 10560
rect 17218 10548 17224 10600
rect 17276 10548 17282 10600
rect 17696 10588 17724 10628
rect 17773 10625 17785 10659
rect 17819 10656 17831 10659
rect 18230 10656 18236 10668
rect 17819 10628 18236 10656
rect 17819 10625 17831 10628
rect 17773 10619 17831 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 19536 10656 19564 10752
rect 20432 10727 20490 10733
rect 20432 10693 20444 10727
rect 20478 10724 20490 10727
rect 21082 10724 21088 10736
rect 20478 10696 21088 10724
rect 20478 10693 20490 10696
rect 20432 10687 20490 10693
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 21634 10684 21640 10736
rect 21692 10684 21698 10736
rect 22278 10684 22284 10736
rect 22336 10684 22342 10736
rect 22388 10696 23060 10724
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19536 10628 19625 10656
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 21652 10656 21680 10684
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 19613 10619 19671 10625
rect 19904 10628 21588 10656
rect 21652 10628 22017 10656
rect 18046 10588 18052 10600
rect 17696 10560 18052 10588
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 18690 10588 18696 10600
rect 18187 10560 18696 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 19904 10520 19932 10628
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 20036 10560 20177 10588
rect 20036 10548 20042 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 21450 10548 21456 10600
rect 21508 10548 21514 10600
rect 21560 10588 21588 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22296 10656 22324 10684
rect 22388 10665 22416 10696
rect 23032 10665 23060 10696
rect 23106 10684 23112 10736
rect 23164 10684 23170 10736
rect 23290 10724 23296 10736
rect 23216 10696 23296 10724
rect 22005 10619 22063 10625
rect 22112 10628 22324 10656
rect 22373 10659 22431 10665
rect 22112 10588 22140 10628
rect 22373 10625 22385 10659
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 23017 10659 23075 10665
rect 23017 10625 23029 10659
rect 23063 10656 23075 10659
rect 23216 10656 23244 10696
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 23400 10668 23428 10764
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24486 10792 24492 10804
rect 24259 10764 24492 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 25038 10752 25044 10804
rect 25096 10752 25102 10804
rect 26142 10752 26148 10804
rect 26200 10792 26206 10804
rect 27249 10795 27307 10801
rect 26200 10764 26924 10792
rect 26200 10752 26206 10764
rect 23934 10684 23940 10736
rect 23992 10724 23998 10736
rect 24581 10727 24639 10733
rect 23992 10696 24164 10724
rect 23992 10684 23998 10696
rect 23382 10656 23388 10668
rect 23063 10628 23244 10656
rect 23308 10628 23388 10656
rect 23063 10625 23075 10628
rect 23017 10619 23075 10625
rect 22848 10588 22876 10619
rect 23308 10597 23336 10628
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 24136 10665 24164 10696
rect 24581 10693 24593 10727
rect 24627 10724 24639 10727
rect 24946 10724 24952 10736
rect 24627 10696 24952 10724
rect 24627 10693 24639 10696
rect 24581 10687 24639 10693
rect 24946 10684 24952 10696
rect 25004 10684 25010 10736
rect 25056 10724 25084 10752
rect 25133 10727 25191 10733
rect 25133 10724 25145 10727
rect 25056 10696 25145 10724
rect 25133 10693 25145 10696
rect 25179 10693 25191 10727
rect 25133 10687 25191 10693
rect 25584 10727 25642 10733
rect 25584 10693 25596 10727
rect 25630 10724 25642 10727
rect 26786 10724 26792 10736
rect 25630 10696 26792 10724
rect 25630 10693 25642 10696
rect 25584 10687 25642 10693
rect 26786 10684 26792 10696
rect 26844 10684 26850 10736
rect 26896 10724 26924 10764
rect 27249 10761 27261 10795
rect 27295 10792 27307 10795
rect 27338 10792 27344 10804
rect 27295 10764 27344 10792
rect 27295 10761 27307 10764
rect 27249 10755 27307 10761
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 28169 10727 28227 10733
rect 28169 10724 28181 10727
rect 26896 10696 28181 10724
rect 28169 10693 28181 10696
rect 28215 10693 28227 10727
rect 28169 10687 28227 10693
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 26418 10656 26424 10668
rect 25280 10628 26424 10656
rect 25280 10616 25286 10628
rect 26418 10616 26424 10628
rect 26476 10616 26482 10668
rect 26878 10616 26884 10668
rect 26936 10656 26942 10668
rect 27154 10656 27160 10668
rect 26936 10628 27160 10656
rect 26936 10616 26942 10628
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 27433 10659 27491 10665
rect 27433 10656 27445 10659
rect 27304 10628 27445 10656
rect 27304 10616 27310 10628
rect 27433 10625 27445 10628
rect 27479 10625 27491 10659
rect 27433 10619 27491 10625
rect 28258 10616 28264 10668
rect 28316 10616 28322 10668
rect 21560 10560 22140 10588
rect 22204 10560 22876 10588
rect 23293 10591 23351 10597
rect 19208 10492 19932 10520
rect 21468 10520 21496 10548
rect 22204 10529 22232 10560
rect 23293 10557 23305 10591
rect 23339 10557 23351 10591
rect 23477 10591 23535 10597
rect 23477 10588 23489 10591
rect 23293 10551 23351 10557
rect 23400 10560 23489 10588
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 21468 10492 21833 10520
rect 19208 10480 19214 10492
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 22189 10523 22247 10529
rect 22189 10489 22201 10523
rect 22235 10489 22247 10523
rect 22189 10483 22247 10489
rect 22649 10523 22707 10529
rect 22649 10489 22661 10523
rect 22695 10520 22707 10523
rect 23400 10520 23428 10560
rect 23477 10557 23489 10560
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10588 23995 10591
rect 24486 10588 24492 10600
rect 23983 10560 24492 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 25317 10591 25375 10597
rect 25317 10588 25329 10591
rect 24912 10560 25329 10588
rect 24912 10548 24918 10560
rect 25317 10557 25329 10560
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 27522 10548 27528 10600
rect 27580 10548 27586 10600
rect 24762 10520 24768 10532
rect 22695 10492 23428 10520
rect 23492 10492 24768 10520
rect 22695 10489 22707 10492
rect 22649 10483 22707 10489
rect 19702 10452 19708 10464
rect 17144 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 19794 10412 19800 10464
rect 19852 10412 19858 10464
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 21545 10455 21603 10461
rect 21545 10452 21557 10455
rect 21508 10424 21557 10452
rect 21508 10412 21514 10424
rect 21545 10421 21557 10424
rect 21591 10421 21603 10455
rect 21545 10415 21603 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 23492 10452 23520 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 27430 10520 27436 10532
rect 26620 10492 27436 10520
rect 22152 10424 23520 10452
rect 22152 10412 22158 10424
rect 23566 10412 23572 10464
rect 23624 10452 23630 10464
rect 26620 10452 26648 10492
rect 27430 10480 27436 10492
rect 27488 10480 27494 10532
rect 23624 10424 26648 10452
rect 23624 10412 23630 10424
rect 26694 10412 26700 10464
rect 26752 10412 26758 10464
rect 26973 10455 27031 10461
rect 26973 10421 26985 10455
rect 27019 10452 27031 10455
rect 27706 10452 27712 10464
rect 27019 10424 27712 10452
rect 27019 10421 27031 10424
rect 26973 10415 27031 10421
rect 27706 10412 27712 10424
rect 27764 10412 27770 10464
rect 28353 10455 28411 10461
rect 28353 10421 28365 10455
rect 28399 10452 28411 10455
rect 28399 10424 28948 10452
rect 28399 10421 28411 10424
rect 28353 10415 28411 10421
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2866 10248 2872 10260
rect 2363 10220 2872 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3326 10248 3332 10260
rect 3068 10220 3332 10248
rect 1581 10183 1639 10189
rect 1581 10149 1593 10183
rect 1627 10180 1639 10183
rect 3068 10180 3096 10220
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 4338 10248 4344 10260
rect 3436 10220 4344 10248
rect 1627 10152 3096 10180
rect 3145 10183 3203 10189
rect 1627 10149 1639 10152
rect 1581 10143 1639 10149
rect 3145 10149 3157 10183
rect 3191 10149 3203 10183
rect 3145 10143 3203 10149
rect 2590 10072 2596 10124
rect 2648 10072 2654 10124
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 2608 10044 2636 10072
rect 2547 10016 2636 10044
rect 3053 10047 3111 10053
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3160 10044 3188 10143
rect 3436 10053 3464 10220
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 4890 10208 4896 10260
rect 4948 10208 4954 10260
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 5718 10248 5724 10260
rect 5491 10220 5724 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5902 10208 5908 10260
rect 5960 10208 5966 10260
rect 7834 10208 7840 10260
rect 7892 10208 7898 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 8076 10220 8309 10248
rect 8076 10208 8082 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 15286 10248 15292 10260
rect 11848 10220 15292 10248
rect 11848 10208 11854 10220
rect 15286 10208 15292 10220
rect 15344 10248 15350 10260
rect 15344 10220 15976 10248
rect 15344 10208 15350 10220
rect 5920 10180 5948 10208
rect 4172 10152 5948 10180
rect 6641 10183 6699 10189
rect 4172 10053 4200 10152
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 7650 10180 7656 10192
rect 6687 10152 7656 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 7852 10180 7880 10208
rect 8386 10180 8392 10192
rect 7852 10152 8392 10180
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 13906 10180 13912 10192
rect 9324 10152 13912 10180
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10112 5227 10115
rect 5534 10112 5540 10124
rect 5215 10084 5540 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5644 10084 8432 10112
rect 5644 10056 5672 10084
rect 3099 10016 3188 10044
rect 3329 10047 3387 10053
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3421 10047 3479 10053
rect 3421 10044 3433 10047
rect 3375 10016 3433 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3421 10013 3433 10016
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5258 10044 5264 10056
rect 5123 10016 5264 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5350 10004 5356 10056
rect 5408 10004 5414 10056
rect 5442 10004 5448 10056
rect 5500 10004 5506 10056
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 6871 10016 6929 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 2593 9979 2651 9985
rect 2593 9945 2605 9979
rect 2639 9976 2651 9979
rect 2958 9976 2964 9988
rect 2639 9948 2964 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3513 9979 3571 9985
rect 3513 9945 3525 9979
rect 3559 9976 3571 9979
rect 4430 9976 4436 9988
rect 3559 9948 4436 9976
rect 3559 9945 3571 9948
rect 3513 9939 3571 9945
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 5460 9976 5488 10004
rect 6365 9979 6423 9985
rect 6365 9976 6377 9979
rect 5460 9948 6377 9976
rect 6365 9945 6377 9948
rect 6411 9945 6423 9979
rect 6365 9939 6423 9945
rect 6932 9920 6960 10007
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7064 10016 7205 10044
rect 7064 10004 7070 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7558 10044 7564 10056
rect 7515 10016 7564 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7285 9979 7343 9985
rect 7285 9945 7297 9979
rect 7331 9976 7343 9979
rect 7668 9976 7696 10007
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 7800 10016 8217 10044
rect 7800 10004 7806 10016
rect 8205 10013 8217 10016
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 7331 9948 7696 9976
rect 8404 9976 8432 10084
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 9324 10044 9352 10152
rect 13906 10140 13912 10152
rect 13964 10140 13970 10192
rect 11517 10115 11575 10121
rect 9508 10084 10456 10112
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 8536 10016 9413 10044
rect 8536 10004 8542 10016
rect 9401 10013 9413 10016
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9508 9976 9536 10084
rect 10428 10056 10456 10084
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11882 10112 11888 10124
rect 11563 10084 11888 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12342 10072 12348 10124
rect 12400 10072 12406 10124
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10468 10016 11284 10044
rect 10468 10004 10474 10016
rect 8404 9948 9536 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 11149 9979 11207 9985
rect 11149 9976 11161 9979
rect 9824 9948 11161 9976
rect 9824 9936 9830 9948
rect 11149 9945 11161 9948
rect 11195 9945 11207 9979
rect 11256 9976 11284 10016
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 13722 10004 13728 10056
rect 13780 10053 13786 10056
rect 13780 10044 13791 10053
rect 15304 10044 15332 10208
rect 15378 10140 15384 10192
rect 15436 10180 15442 10192
rect 15948 10180 15976 10220
rect 16022 10208 16028 10260
rect 16080 10208 16086 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 17276 10220 17601 10248
rect 17276 10208 17282 10220
rect 17589 10217 17601 10220
rect 17635 10217 17647 10251
rect 17589 10211 17647 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 21177 10251 21235 10257
rect 18012 10220 21036 10248
rect 18012 10208 18018 10220
rect 19061 10183 19119 10189
rect 15436 10152 15516 10180
rect 15948 10152 18736 10180
rect 15436 10140 15442 10152
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 13780 10016 13825 10044
rect 15304 10016 15393 10044
rect 13780 10007 13791 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15488 10044 15516 10152
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10112 15623 10115
rect 16209 10115 16267 10121
rect 16209 10112 16221 10115
rect 15611 10084 16221 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 16209 10081 16221 10084
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 16758 10072 16764 10124
rect 16816 10072 16822 10124
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17957 10115 18015 10121
rect 17276 10084 17540 10112
rect 17276 10072 17282 10084
rect 16114 10044 16120 10056
rect 15488 10016 16120 10044
rect 15381 10007 15439 10013
rect 13780 10004 13786 10007
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 16776 10044 16804 10072
rect 17512 10053 17540 10084
rect 17957 10081 17969 10115
rect 18003 10112 18015 10115
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18003 10084 18613 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18708 10112 18736 10152
rect 19061 10149 19073 10183
rect 19107 10180 19119 10183
rect 19426 10180 19432 10192
rect 19107 10152 19432 10180
rect 19107 10149 19119 10152
rect 19061 10143 19119 10149
rect 19426 10140 19432 10152
rect 19484 10180 19490 10192
rect 19613 10183 19671 10189
rect 19613 10180 19625 10183
rect 19484 10152 19625 10180
rect 19484 10140 19490 10152
rect 19613 10149 19625 10152
rect 19659 10149 19671 10183
rect 19613 10143 19671 10149
rect 19150 10112 19156 10124
rect 18708 10084 19156 10112
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 16776 10016 17417 10044
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17543 10016 17877 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 18708 10044 18736 10084
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19245 10115 19303 10121
rect 19245 10081 19257 10115
rect 19291 10112 19303 10115
rect 19702 10112 19708 10124
rect 19291 10084 19708 10112
rect 19291 10081 19303 10084
rect 19245 10075 19303 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 18463 10016 18736 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 16298 9976 16304 9988
rect 11256 9948 16304 9976
rect 11149 9939 11207 9945
rect 16298 9936 16304 9948
rect 16356 9976 16362 9988
rect 18230 9976 18236 9988
rect 16356 9948 18236 9976
rect 16356 9936 16362 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 18340 9976 18368 10007
rect 18782 10004 18788 10056
rect 18840 10004 18846 10056
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 19024 10038 19104 10044
rect 19306 10038 19441 10044
rect 19024 10016 19441 10038
rect 19024 10004 19030 10016
rect 19076 10010 19334 10016
rect 19429 10013 19441 10016
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20165 10047 20223 10053
rect 20165 10044 20177 10047
rect 19944 10016 20177 10044
rect 19944 10004 19950 10016
rect 20165 10013 20177 10016
rect 20211 10044 20223 10047
rect 20898 10044 20904 10056
rect 20211 10016 20904 10044
rect 20211 10013 20223 10016
rect 20165 10007 20223 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 18800 9976 18828 10004
rect 18340 9948 18828 9976
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 18932 9948 19196 9976
rect 18932 9936 18938 9948
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 5718 9908 5724 9920
rect 4019 9880 5724 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 7006 9868 7012 9920
rect 7064 9868 7070 9920
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 10137 9911 10195 9917
rect 10137 9877 10149 9911
rect 10183 9908 10195 9911
rect 11790 9908 11796 9920
rect 10183 9880 11796 9908
rect 10183 9877 10195 9880
rect 10137 9871 10195 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 11940 9880 12173 9908
rect 11940 9868 11946 9880
rect 12161 9877 12173 9880
rect 12207 9908 12219 9911
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12207 9880 13001 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 14090 9908 14096 9920
rect 13587 9880 14096 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 17034 9908 17040 9920
rect 14608 9880 17040 9908
rect 14608 9868 14614 9880
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 17221 9911 17279 9917
rect 17221 9877 17233 9911
rect 17267 9908 17279 9911
rect 17678 9908 17684 9920
rect 17267 9880 17684 9908
rect 17267 9877 17279 9880
rect 17221 9871 17279 9877
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18966 9908 18972 9920
rect 18187 9880 18972 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19168 9908 19196 9948
rect 19306 9948 20668 9976
rect 19306 9908 19334 9948
rect 19168 9880 19334 9908
rect 20640 9908 20668 9948
rect 20714 9936 20720 9988
rect 20772 9936 20778 9988
rect 21008 9976 21036 10220
rect 21177 10217 21189 10251
rect 21223 10248 21235 10251
rect 22094 10248 22100 10260
rect 21223 10220 22100 10248
rect 21223 10217 21235 10220
rect 21177 10211 21235 10217
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 22281 10251 22339 10257
rect 22281 10217 22293 10251
rect 22327 10248 22339 10251
rect 22327 10220 23060 10248
rect 22327 10217 22339 10220
rect 22281 10211 22339 10217
rect 21358 10140 21364 10192
rect 21416 10140 21422 10192
rect 21634 10180 21640 10192
rect 21468 10152 21640 10180
rect 21082 10004 21088 10056
rect 21140 10004 21146 10056
rect 21468 10044 21496 10152
rect 21634 10140 21640 10152
rect 21692 10180 21698 10192
rect 21913 10183 21971 10189
rect 21692 10152 21864 10180
rect 21692 10140 21698 10152
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 21836 10112 21864 10152
rect 21913 10149 21925 10183
rect 21959 10180 21971 10183
rect 22925 10183 22983 10189
rect 21959 10152 22692 10180
rect 21959 10149 21971 10152
rect 21913 10143 21971 10149
rect 22664 10121 22692 10152
rect 22925 10149 22937 10183
rect 22971 10149 22983 10183
rect 23032 10180 23060 10220
rect 23198 10208 23204 10260
rect 23256 10248 23262 10260
rect 23293 10251 23351 10257
rect 23293 10248 23305 10251
rect 23256 10220 23305 10248
rect 23256 10208 23262 10220
rect 23293 10217 23305 10220
rect 23339 10217 23351 10251
rect 23293 10211 23351 10217
rect 23661 10251 23719 10257
rect 23661 10217 23673 10251
rect 23707 10248 23719 10251
rect 24118 10248 24124 10260
rect 23707 10220 24124 10248
rect 23707 10217 23719 10220
rect 23661 10211 23719 10217
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 24486 10208 24492 10260
rect 24544 10248 24550 10260
rect 24765 10251 24823 10257
rect 24765 10248 24777 10251
rect 24544 10220 24777 10248
rect 24544 10208 24550 10220
rect 24765 10217 24777 10220
rect 24811 10217 24823 10251
rect 27062 10248 27068 10260
rect 24765 10211 24823 10217
rect 26252 10220 27068 10248
rect 26252 10180 26280 10220
rect 27062 10208 27068 10220
rect 27120 10208 27126 10260
rect 28920 10180 28948 10424
rect 23032 10152 26280 10180
rect 26344 10152 28948 10180
rect 22925 10143 22983 10149
rect 22649 10115 22707 10121
rect 21836 10084 22600 10112
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 21468 10016 21557 10044
rect 21545 10013 21557 10016
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 21637 10047 21695 10053
rect 21637 10013 21649 10047
rect 21683 10013 21695 10047
rect 21744 10044 21772 10072
rect 22097 10047 22155 10053
rect 22097 10044 22109 10047
rect 21744 10016 22109 10044
rect 21637 10007 21695 10013
rect 22097 10013 22109 10016
rect 22143 10013 22155 10047
rect 22097 10007 22155 10013
rect 21652 9976 21680 10007
rect 22186 10004 22192 10056
rect 22244 10004 22250 10056
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10013 22523 10047
rect 22572 10044 22600 10084
rect 22649 10081 22661 10115
rect 22695 10081 22707 10115
rect 22940 10112 22968 10143
rect 23014 10112 23020 10124
rect 22940 10084 23020 10112
rect 22649 10075 22707 10081
rect 23014 10072 23020 10084
rect 23072 10072 23078 10124
rect 23106 10072 23112 10124
rect 23164 10112 23170 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 23164 10084 24593 10112
rect 23164 10072 23170 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 25038 10072 25044 10124
rect 25096 10112 25102 10124
rect 25225 10115 25283 10121
rect 25225 10112 25237 10115
rect 25096 10084 25237 10112
rect 25096 10072 25102 10084
rect 25225 10081 25237 10084
rect 25271 10081 25283 10115
rect 25225 10075 25283 10081
rect 26142 10072 26148 10124
rect 26200 10072 26206 10124
rect 26234 10072 26240 10124
rect 26292 10072 26298 10124
rect 26344 10121 26372 10152
rect 26329 10115 26387 10121
rect 26329 10081 26341 10115
rect 26375 10081 26387 10115
rect 26329 10075 26387 10081
rect 26694 10072 26700 10124
rect 26752 10112 26758 10124
rect 27065 10115 27123 10121
rect 27065 10112 27077 10115
rect 26752 10084 27077 10112
rect 26752 10072 26758 10084
rect 27065 10081 27077 10084
rect 27111 10081 27123 10115
rect 27065 10075 27123 10081
rect 27801 10115 27859 10121
rect 27801 10081 27813 10115
rect 27847 10112 27859 10115
rect 28258 10112 28264 10124
rect 27847 10084 28264 10112
rect 27847 10081 27859 10084
rect 27801 10075 27859 10081
rect 28258 10072 28264 10084
rect 28316 10072 28322 10124
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 22572 10016 23213 10044
rect 22465 10007 22523 10013
rect 23201 10013 23213 10016
rect 23247 10044 23259 10047
rect 23290 10044 23296 10056
rect 23247 10016 23296 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 22480 9976 22508 10007
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 23842 10004 23848 10056
rect 23900 10004 23906 10056
rect 23934 10004 23940 10056
rect 23992 10044 23998 10056
rect 24121 10047 24179 10053
rect 24121 10044 24133 10047
rect 23992 10016 24133 10044
rect 23992 10004 23998 10016
rect 24121 10013 24133 10016
rect 24167 10013 24179 10047
rect 24121 10007 24179 10013
rect 24210 10004 24216 10056
rect 24268 10044 24274 10056
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 24268 10016 24409 10044
rect 24268 10004 24274 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 26252 10044 26280 10072
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 26252 10016 26525 10044
rect 24397 10007 24455 10013
rect 26513 10013 26525 10016
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 27982 10004 27988 10056
rect 28040 10004 28046 10056
rect 23566 9976 23572 9988
rect 21008 9948 21680 9976
rect 21744 9948 23572 9976
rect 21744 9908 21772 9948
rect 23566 9936 23572 9948
rect 23624 9936 23630 9988
rect 25317 9979 25375 9985
rect 25317 9945 25329 9979
rect 25363 9945 25375 9979
rect 28534 9976 28540 9988
rect 25317 9939 25375 9945
rect 26896 9948 28540 9976
rect 20640 9880 21772 9908
rect 21821 9911 21879 9917
rect 21821 9877 21833 9911
rect 21867 9908 21879 9911
rect 23474 9908 23480 9920
rect 21867 9880 23480 9908
rect 21867 9877 21879 9880
rect 21821 9871 21879 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 23937 9911 23995 9917
rect 23937 9877 23949 9911
rect 23983 9908 23995 9911
rect 24946 9908 24952 9920
rect 23983 9880 24952 9908
rect 23983 9877 23995 9880
rect 23937 9871 23995 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 25130 9868 25136 9920
rect 25188 9908 25194 9920
rect 25325 9908 25353 9939
rect 25188 9880 25353 9908
rect 25188 9868 25194 9880
rect 25406 9868 25412 9920
rect 25464 9908 25470 9920
rect 26896 9908 26924 9948
rect 28534 9936 28540 9948
rect 28592 9936 28598 9988
rect 25464 9880 26924 9908
rect 26973 9911 27031 9917
rect 25464 9868 25470 9880
rect 26973 9877 26985 9911
rect 27019 9908 27031 9911
rect 27614 9908 27620 9920
rect 27019 9880 27620 9908
rect 27019 9877 27031 9880
rect 26973 9871 27031 9877
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 27709 9911 27767 9917
rect 27709 9877 27721 9911
rect 27755 9908 27767 9911
rect 27798 9908 27804 9920
rect 27755 9880 27804 9908
rect 27755 9877 27767 9880
rect 27709 9871 27767 9877
rect 27798 9868 27804 9880
rect 27856 9868 27862 9920
rect 28442 9868 28448 9920
rect 28500 9868 28506 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2924 9676 3924 9704
rect 2924 9664 2930 9676
rect 3050 9596 3056 9648
rect 3108 9596 3114 9648
rect 3896 9645 3924 9676
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 7193 9707 7251 9713
rect 5592 9676 6592 9704
rect 5592 9664 5598 9676
rect 3881 9639 3939 9645
rect 3881 9605 3893 9639
rect 3927 9605 3939 9639
rect 3881 9599 3939 9605
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 5626 9636 5632 9648
rect 5307 9608 5632 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6086 9596 6092 9648
rect 6144 9596 6150 9648
rect 6564 9645 6592 9676
rect 7193 9673 7205 9707
rect 7239 9673 7251 9707
rect 7193 9667 7251 9673
rect 8849 9707 8907 9713
rect 8849 9673 8861 9707
rect 8895 9704 8907 9707
rect 9582 9704 9588 9716
rect 8895 9676 9588 9704
rect 8895 9673 8907 9676
rect 8849 9667 8907 9673
rect 6549 9639 6607 9645
rect 6549 9605 6561 9639
rect 6595 9605 6607 9639
rect 7208 9636 7236 9667
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11756 9676 11805 9704
rect 11756 9664 11762 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 12345 9707 12403 9713
rect 12345 9673 12357 9707
rect 12391 9704 12403 9707
rect 12526 9704 12532 9716
rect 12391 9676 12532 9704
rect 12391 9673 12403 9676
rect 12345 9667 12403 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13906 9704 13912 9716
rect 13740 9676 13912 9704
rect 7653 9639 7711 9645
rect 7653 9636 7665 9639
rect 7208 9608 7665 9636
rect 6549 9599 6607 9605
rect 7653 9605 7665 9608
rect 7699 9605 7711 9639
rect 7653 9599 7711 9605
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8444 9608 8585 9636
rect 8444 9596 8450 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8573 9599 8631 9605
rect 8680 9608 9168 9636
rect 8680 9580 8708 9608
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 1872 9500 1900 9531
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4488 9540 4721 9568
rect 4488 9528 4494 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4798 9528 4804 9580
rect 4856 9528 4862 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 9030 9528 9036 9580
rect 9088 9528 9094 9580
rect 9140 9577 9168 9608
rect 11716 9608 12848 9636
rect 11716 9577 11744 9608
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 9539 9540 10977 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 11848 9540 12173 9568
rect 11848 9528 11854 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12575 9540 12664 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 1412 9472 1900 9500
rect 1412 9441 1440 9472
rect 2130 9460 2136 9512
rect 2188 9460 2194 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 1397 9435 1455 9441
rect 1397 9401 1409 9435
rect 1443 9401 1455 9435
rect 1397 9395 1455 9401
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 2332 9432 2360 9463
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 2832 9472 2973 9500
rect 2832 9460 2838 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 2961 9463 3019 9469
rect 3620 9472 3801 9500
rect 1820 9404 2360 9432
rect 3513 9435 3571 9441
rect 1820 9392 1826 9404
rect 3513 9401 3525 9435
rect 3559 9432 3571 9435
rect 3620 9432 3648 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4816 9500 4844 9528
rect 4571 9472 4844 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5408 9472 6469 9500
rect 5408 9460 5414 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 7558 9460 7564 9512
rect 7616 9460 7622 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 3559 9404 3648 9432
rect 3559 9401 3571 9404
rect 3513 9395 3571 9401
rect 3620 9376 3648 9404
rect 4341 9435 4399 9441
rect 4341 9401 4353 9435
rect 4387 9432 4399 9435
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4387 9404 4905 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4893 9401 4905 9404
rect 4939 9432 4951 9435
rect 5258 9432 5264 9444
rect 4939 9404 5264 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6972 9404 7021 9432
rect 6972 9392 6978 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 9692 9432 9720 9463
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 10100 9472 10241 9500
rect 10100 9460 10106 9472
rect 10229 9469 10241 9472
rect 10275 9469 10287 9503
rect 10229 9463 10287 9469
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 10870 9500 10876 9512
rect 10459 9472 10876 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 12636 9441 12664 9540
rect 12710 9528 12716 9580
rect 12768 9528 12774 9580
rect 12820 9577 12848 9608
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 13538 9568 13544 9580
rect 12851 9540 13544 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 13740 9577 13768 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 14090 9664 14096 9716
rect 14148 9664 14154 9716
rect 14642 9664 14648 9716
rect 14700 9664 14706 9716
rect 19260 9676 20576 9704
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 14108 9568 14136 9664
rect 14660 9636 14688 9664
rect 18874 9636 18880 9648
rect 14660 9608 14964 9636
rect 14936 9577 14964 9608
rect 17144 9608 18880 9636
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 14108 9540 14657 9568
rect 13725 9531 13783 9537
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15657 9571 15715 9577
rect 15657 9537 15669 9571
rect 15703 9568 15715 9571
rect 16022 9568 16028 9580
rect 15703 9540 16028 9568
rect 15703 9537 15715 9540
rect 15657 9531 15715 9537
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 17144 9577 17172 9608
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 19260 9636 19288 9676
rect 18984 9608 19288 9636
rect 20548 9636 20576 9676
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21174 9704 21180 9716
rect 20772 9676 21180 9704
rect 20772 9664 20778 9676
rect 21174 9664 21180 9676
rect 21232 9704 21238 9716
rect 21634 9704 21640 9716
rect 21232 9676 21640 9704
rect 21232 9664 21238 9676
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21821 9707 21879 9713
rect 21821 9673 21833 9707
rect 21867 9704 21879 9707
rect 23750 9704 23756 9716
rect 21867 9676 23756 9704
rect 21867 9673 21879 9676
rect 21821 9667 21879 9673
rect 23750 9664 23756 9676
rect 23808 9664 23814 9716
rect 23842 9664 23848 9716
rect 23900 9704 23906 9716
rect 23900 9676 24808 9704
rect 23900 9664 23906 9676
rect 20548 9608 20944 9636
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 12728 9500 12756 9528
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12728 9472 13001 9500
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 13955 9472 14504 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14476 9441 14504 9472
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 15838 9460 15844 9512
rect 15896 9460 15902 9512
rect 17052 9500 17080 9531
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17460 9540 17877 9568
rect 17460 9528 17466 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18196 9540 18613 9568
rect 18196 9528 18202 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 17052 9472 17264 9500
rect 11977 9435 12035 9441
rect 11977 9432 11989 9435
rect 9692 9404 11989 9432
rect 7009 9395 7067 9401
rect 11977 9401 11989 9404
rect 12023 9401 12035 9435
rect 11977 9395 12035 9401
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 14461 9435 14519 9441
rect 14461 9401 14473 9435
rect 14507 9401 14519 9435
rect 14461 9395 14519 9401
rect 17236 9376 17264 9472
rect 17310 9460 17316 9512
rect 17368 9460 17374 9512
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 17678 9392 17684 9444
rect 17736 9432 17742 9444
rect 18984 9432 19012 9608
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19208 9540 20269 9568
rect 19208 9528 19214 9540
rect 20088 9512 20116 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20346 9528 20352 9580
rect 20404 9528 20410 9580
rect 20622 9528 20628 9580
rect 20680 9528 20686 9580
rect 20916 9577 20944 9608
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21266 9568 21272 9580
rect 21223 9540 21272 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21266 9528 21272 9540
rect 21324 9568 21330 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21324 9540 21465 9568
rect 21324 9528 21330 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 22738 9568 22744 9580
rect 22060 9540 22744 9568
rect 22060 9528 22066 9540
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 22830 9528 22836 9580
rect 22888 9528 22894 9580
rect 23017 9571 23075 9577
rect 23017 9537 23029 9571
rect 23063 9568 23075 9571
rect 23198 9568 23204 9580
rect 23063 9540 23204 9568
rect 23063 9537 23075 9540
rect 23017 9531 23075 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 23290 9528 23296 9580
rect 23348 9568 23354 9580
rect 23661 9571 23719 9577
rect 23661 9568 23673 9571
rect 23348 9540 23673 9568
rect 23348 9528 23354 9540
rect 23661 9537 23673 9540
rect 23707 9568 23719 9571
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 23707 9540 24685 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 24673 9537 24685 9540
rect 24719 9537 24731 9571
rect 24780 9568 24808 9676
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 25004 9676 25912 9704
rect 25004 9664 25010 9676
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25409 9639 25467 9645
rect 25409 9636 25421 9639
rect 24912 9608 25421 9636
rect 24912 9596 24918 9608
rect 25409 9605 25421 9608
rect 25455 9605 25467 9639
rect 25409 9599 25467 9605
rect 25884 9577 25912 9676
rect 26694 9664 26700 9716
rect 26752 9664 26758 9716
rect 27706 9664 27712 9716
rect 27764 9664 27770 9716
rect 27982 9664 27988 9716
rect 28040 9704 28046 9716
rect 28169 9707 28227 9713
rect 28169 9704 28181 9707
rect 28040 9676 28181 9704
rect 28040 9664 28046 9676
rect 28169 9673 28181 9676
rect 28215 9673 28227 9707
rect 28169 9667 28227 9673
rect 28442 9664 28448 9716
rect 28500 9664 28506 9716
rect 25958 9596 25964 9648
rect 26016 9636 26022 9648
rect 26712 9636 26740 9664
rect 26016 9608 26556 9636
rect 26712 9608 27016 9636
rect 26016 9596 26022 9608
rect 25869 9571 25927 9577
rect 24780 9540 25452 9568
rect 24673 9531 24731 9537
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9500 19395 9503
rect 19426 9500 19432 9512
rect 19383 9472 19432 9500
rect 19383 9469 19395 9472
rect 19337 9463 19395 9469
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19518 9460 19524 9512
rect 19576 9460 19582 9512
rect 20070 9460 20076 9512
rect 20128 9460 20134 9512
rect 21726 9460 21732 9512
rect 21784 9460 21790 9512
rect 22094 9460 22100 9512
rect 22152 9460 22158 9512
rect 22278 9460 22284 9512
rect 22336 9460 22342 9512
rect 24489 9503 24547 9509
rect 24489 9469 24501 9503
rect 24535 9500 24547 9503
rect 24946 9500 24952 9512
rect 24535 9472 24952 9500
rect 24535 9469 24547 9472
rect 24489 9463 24547 9469
rect 24946 9460 24952 9472
rect 25004 9460 25010 9512
rect 17736 9404 19012 9432
rect 19245 9435 19303 9441
rect 17736 9392 17742 9404
rect 19245 9401 19257 9435
rect 19291 9432 19303 9435
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 19291 9404 19993 9432
rect 19291 9401 19303 9404
rect 19245 9395 19303 9401
rect 19981 9401 19993 9404
rect 20027 9432 20039 9435
rect 20027 9404 20208 9432
rect 20027 9401 20039 9404
rect 19981 9395 20039 9401
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 2222 9364 2228 9376
rect 1719 9336 2228 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 8478 9364 8484 9376
rect 3936 9336 8484 9364
rect 3936 9324 3942 9336
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10594 9364 10600 9376
rect 10183 9336 10600 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 14090 9364 14096 9376
rect 13679 9336 14096 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15528 9336 16037 9364
rect 15528 9324 15534 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17218 9324 17224 9376
rect 17276 9324 17282 9376
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 17828 9336 18245 9364
rect 17828 9324 17834 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 19702 9324 19708 9376
rect 19760 9364 19766 9376
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 19760 9336 20085 9364
rect 19760 9324 19766 9336
rect 20073 9333 20085 9336
rect 20119 9333 20131 9367
rect 20180 9364 20208 9404
rect 20346 9364 20352 9376
rect 20180 9336 20352 9364
rect 20073 9327 20131 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20438 9324 20444 9376
rect 20496 9324 20502 9376
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 21266 9324 21272 9376
rect 21324 9324 21330 9376
rect 21637 9367 21695 9373
rect 21637 9333 21649 9367
rect 21683 9364 21695 9367
rect 21744 9364 21772 9460
rect 23106 9392 23112 9444
rect 23164 9432 23170 9444
rect 23201 9435 23259 9441
rect 23201 9432 23213 9435
rect 23164 9404 23213 9432
rect 23164 9392 23170 9404
rect 23201 9401 23213 9404
rect 23247 9401 23259 9435
rect 25424 9432 25452 9540
rect 25869 9537 25881 9571
rect 25915 9537 25927 9571
rect 25869 9531 25927 9537
rect 26234 9528 26240 9580
rect 26292 9568 26298 9580
rect 26528 9577 26556 9608
rect 26513 9571 26571 9577
rect 26292 9540 26464 9568
rect 26292 9528 26298 9540
rect 26053 9435 26111 9441
rect 26053 9432 26065 9435
rect 25424 9404 26065 9432
rect 23201 9395 23259 9401
rect 26053 9401 26065 9404
rect 26099 9401 26111 9435
rect 26053 9395 26111 9401
rect 21683 9336 21772 9364
rect 21683 9333 21695 9336
rect 21637 9327 21695 9333
rect 22738 9324 22744 9376
rect 22796 9324 22802 9376
rect 25038 9324 25044 9376
rect 25096 9364 25102 9376
rect 25685 9367 25743 9373
rect 25685 9364 25697 9367
rect 25096 9336 25697 9364
rect 25096 9324 25102 9336
rect 25685 9333 25697 9336
rect 25731 9333 25743 9367
rect 25685 9327 25743 9333
rect 26326 9324 26332 9376
rect 26384 9324 26390 9376
rect 26436 9364 26464 9540
rect 26513 9537 26525 9571
rect 26559 9537 26571 9571
rect 26513 9531 26571 9537
rect 26786 9528 26792 9580
rect 26844 9528 26850 9580
rect 26988 9577 27016 9608
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9537 27031 9571
rect 26973 9531 27031 9537
rect 27062 9528 27068 9580
rect 27120 9568 27126 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27120 9540 27445 9568
rect 27120 9528 27126 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27724 9568 27752 9664
rect 27890 9596 27896 9648
rect 27948 9636 27954 9648
rect 28077 9639 28135 9645
rect 28077 9636 28089 9639
rect 27948 9608 28089 9636
rect 27948 9596 27954 9608
rect 28077 9605 28089 9608
rect 28123 9636 28135 9639
rect 28460 9636 28488 9664
rect 28123 9608 28488 9636
rect 28123 9605 28135 9608
rect 28077 9599 28135 9605
rect 28353 9571 28411 9577
rect 28353 9568 28365 9571
rect 27724 9540 28365 9568
rect 27433 9531 27491 9537
rect 28353 9537 28365 9540
rect 28399 9537 28411 9571
rect 28353 9531 28411 9537
rect 27338 9460 27344 9512
rect 27396 9500 27402 9512
rect 27617 9503 27675 9509
rect 27617 9500 27629 9503
rect 27396 9472 27629 9500
rect 27396 9460 27402 9472
rect 27617 9469 27629 9472
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 26605 9435 26663 9441
rect 26605 9401 26617 9435
rect 26651 9432 26663 9435
rect 27982 9432 27988 9444
rect 26651 9404 27988 9432
rect 26651 9401 26663 9404
rect 26605 9395 26663 9401
rect 27982 9392 27988 9404
rect 28040 9392 28046 9444
rect 26694 9364 26700 9376
rect 26436 9336 26700 9364
rect 26694 9324 26700 9336
rect 26752 9364 26758 9376
rect 26878 9364 26884 9376
rect 26752 9336 26884 9364
rect 26752 9324 26758 9336
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 27062 9324 27068 9376
rect 27120 9324 27126 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 2130 9120 2136 9172
rect 2188 9120 2194 9172
rect 2774 9120 2780 9172
rect 2832 9120 2838 9172
rect 3510 9120 3516 9172
rect 3568 9120 3574 9172
rect 5350 9120 5356 9172
rect 5408 9120 5414 9172
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7374 9160 7380 9172
rect 6319 9132 7380 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 8352 9132 8401 9160
rect 8352 9120 8358 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9030 9160 9036 9172
rect 8619 9132 9036 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9214 9120 9220 9172
rect 9272 9120 9278 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9160 9827 9163
rect 10042 9160 10048 9172
rect 9815 9132 10048 9160
rect 9815 9129 9827 9132
rect 9769 9123 9827 9129
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10594 9120 10600 9172
rect 10652 9120 10658 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13817 9163 13875 9169
rect 13817 9160 13829 9163
rect 13228 9132 13829 9160
rect 13228 9120 13234 9132
rect 13817 9129 13829 9132
rect 13863 9129 13875 9163
rect 13817 9123 13875 9129
rect 14090 9120 14096 9172
rect 14148 9120 14154 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 15160 9132 15301 9160
rect 15160 9120 15166 9132
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 15838 9160 15844 9172
rect 15703 9132 15844 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 17037 9163 17095 9169
rect 17037 9129 17049 9163
rect 17083 9160 17095 9163
rect 17310 9160 17316 9172
rect 17083 9132 17316 9160
rect 17083 9129 17095 9132
rect 17037 9123 17095 9129
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17405 9163 17463 9169
rect 17405 9129 17417 9163
rect 17451 9160 17463 9163
rect 18046 9160 18052 9172
rect 17451 9132 18052 9160
rect 17451 9129 17463 9132
rect 17405 9123 17463 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 18233 9163 18291 9169
rect 18233 9129 18245 9163
rect 18279 9160 18291 9163
rect 18782 9160 18788 9172
rect 18279 9132 18788 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19518 9160 19524 9172
rect 18923 9132 19524 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19518 9120 19524 9132
rect 19576 9120 19582 9172
rect 20162 9120 20168 9172
rect 20220 9120 20226 9172
rect 21634 9160 21640 9172
rect 20640 9132 21640 9160
rect 2148 9092 2176 9120
rect 6362 9092 6368 9104
rect 2148 9064 4568 9092
rect 3878 9024 3884 9036
rect 2148 8996 2452 9024
rect 2148 8965 2176 8996
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2056 8888 2084 8919
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2280 8928 2329 8956
rect 2280 8916 2286 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2424 8956 2452 8996
rect 2746 8996 3884 9024
rect 2746 8956 2774 8996
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 4246 9024 4252 9036
rect 4019 8996 4252 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 2424 8928 2774 8956
rect 2869 8959 2927 8965
rect 2317 8919 2375 8925
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2884 8888 2912 8919
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 2056 8860 2912 8888
rect 2792 8832 2820 8860
rect 1854 8780 1860 8832
rect 1912 8780 1918 8832
rect 2774 8780 2780 8832
rect 2832 8780 2838 8832
rect 4540 8820 4568 9064
rect 4724 9064 6368 9092
rect 4724 9033 4752 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 7190 9052 7196 9104
rect 7248 9052 7254 9104
rect 8478 9092 8484 9104
rect 7392 9064 8484 9092
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 5316 8996 5549 9024
rect 5316 8984 5322 8996
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6914 9024 6920 9036
rect 6227 8996 6920 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7392 9033 7420 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7616 8996 7665 9024
rect 7616 8984 7622 8996
rect 7653 8993 7665 8996
rect 7699 9024 7711 9027
rect 9232 9024 9260 9120
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 7699 8996 8340 9024
rect 9232 8996 9321 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6503 8928 6653 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6641 8925 6653 8928
rect 6687 8956 6699 8959
rect 6822 8956 6828 8968
rect 6687 8928 6828 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 8312 8965 8340 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 10612 9024 10640 9120
rect 12710 9092 12716 9104
rect 10980 9064 12716 9092
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10612 8996 10885 9024
rect 9309 8987 9367 8993
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8720 8928 8769 8956
rect 8720 8916 8726 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10410 8956 10416 8968
rect 9907 8928 10416 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 4617 8891 4675 8897
rect 4617 8857 4629 8891
rect 4663 8888 4675 8891
rect 5368 8888 5396 8916
rect 4663 8860 5396 8888
rect 5629 8891 5687 8897
rect 4663 8857 4675 8860
rect 4617 8851 4675 8857
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5718 8888 5724 8900
rect 5675 8860 5724 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 7466 8848 7472 8900
rect 7524 8848 7530 8900
rect 9140 8888 9168 8919
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10980 8956 11008 9064
rect 12710 9052 12716 9064
rect 12768 9052 12774 9104
rect 11609 9027 11667 9033
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 11882 9024 11888 9036
rect 11655 8996 11888 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 14108 9033 14136 9120
rect 20640 9104 20668 9132
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22189 9163 22247 9169
rect 22189 9160 22201 9163
rect 22152 9132 22201 9160
rect 22152 9120 22158 9132
rect 22189 9129 22201 9132
rect 22235 9129 22247 9163
rect 22189 9123 22247 9129
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 22796 9132 23673 9160
rect 22796 9120 22802 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 24026 9120 24032 9172
rect 24084 9120 24090 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 25225 9163 25283 9169
rect 25225 9160 25237 9163
rect 25188 9132 25237 9160
rect 25188 9120 25194 9132
rect 25225 9129 25237 9132
rect 25271 9129 25283 9163
rect 26602 9160 26608 9172
rect 25225 9123 25283 9129
rect 25332 9132 26608 9160
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14461 9095 14519 9101
rect 14461 9092 14473 9095
rect 14240 9064 14473 9092
rect 14240 9052 14246 9064
rect 14461 9061 14473 9064
rect 14507 9061 14519 9095
rect 14461 9055 14519 9061
rect 16684 9064 19840 9092
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 9024 14335 9027
rect 14921 9027 14979 9033
rect 14921 9024 14933 9027
rect 14323 8996 14933 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 14921 8993 14933 8996
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 15212 8996 16160 9024
rect 10520 8928 11008 8956
rect 10520 8888 10548 8928
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11756 8928 11805 8956
rect 11756 8916 11762 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 13722 8916 13728 8968
rect 13780 8916 13786 8968
rect 15212 8965 15240 8996
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8956 14887 8959
rect 15197 8959 15255 8965
rect 15197 8956 15209 8959
rect 14875 8928 15209 8956
rect 14875 8925 14887 8928
rect 14829 8919 14887 8925
rect 15197 8925 15209 8928
rect 15243 8925 15255 8959
rect 15197 8919 15255 8925
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 15930 8956 15936 8968
rect 15887 8928 15936 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16132 8965 16160 8996
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16298 8956 16304 8968
rect 16163 8928 16304 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 16482 8956 16488 8968
rect 16439 8928 16488 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16684 8965 16712 9064
rect 16850 8984 16856 9036
rect 16908 8984 16914 9036
rect 19610 9024 19616 9036
rect 17880 8996 19616 9024
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16632 8928 16681 8956
rect 16632 8916 16638 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16758 8916 16764 8968
rect 16816 8916 16822 8968
rect 16868 8956 16896 8984
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 16868 8928 17233 8956
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17310 8916 17316 8968
rect 17368 8916 17374 8968
rect 17880 8965 17908 8996
rect 19610 8984 19616 8996
rect 19668 8984 19674 9036
rect 19702 8984 19708 9036
rect 19760 8984 19766 9036
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 18187 8928 18797 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8925 19119 8959
rect 19061 8919 19119 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 19720 8956 19748 8984
rect 19475 8928 19748 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 8312 8860 10548 8888
rect 8312 8820 8340 8860
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 16022 8848 16028 8900
rect 16080 8888 16086 8900
rect 17788 8888 17816 8919
rect 18156 8888 18184 8919
rect 19076 8888 19104 8919
rect 16080 8860 17816 8888
rect 17880 8860 18184 8888
rect 18616 8860 19104 8888
rect 16080 8848 16086 8860
rect 17880 8832 17908 8860
rect 4540 8792 8340 8820
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8570 8820 8576 8832
rect 8444 8792 8576 8820
rect 8444 8780 8450 8792
rect 8570 8780 8576 8792
rect 8628 8820 8634 8832
rect 9030 8820 9036 8832
rect 8628 8792 9036 8820
rect 8628 8780 8634 8792
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 10560 8792 11529 8820
rect 10560 8780 10566 8792
rect 11517 8789 11529 8792
rect 11563 8820 11575 8823
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 11563 8792 12265 8820
rect 11563 8789 11575 8792
rect 11517 8783 11575 8789
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 12253 8783 12311 8789
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16850 8820 16856 8832
rect 16531 8792 16856 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 16945 8823 17003 8829
rect 16945 8789 16957 8823
rect 16991 8820 17003 8823
rect 17494 8820 17500 8832
rect 16991 8792 17500 8820
rect 16991 8789 17003 8792
rect 16945 8783 17003 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17586 8780 17592 8832
rect 17644 8780 17650 8832
rect 17862 8780 17868 8832
rect 17920 8780 17926 8832
rect 18046 8780 18052 8832
rect 18104 8780 18110 8832
rect 18616 8829 18644 8860
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8789 18659 8823
rect 18601 8783 18659 8789
rect 19610 8780 19616 8832
rect 19668 8780 19674 8832
rect 19702 8780 19708 8832
rect 19760 8780 19766 8832
rect 19812 8820 19840 9064
rect 20622 9052 20628 9104
rect 20680 9052 20686 9104
rect 20993 9095 21051 9101
rect 20993 9061 21005 9095
rect 21039 9092 21051 9095
rect 21453 9095 21511 9101
rect 21453 9092 21465 9095
rect 21039 9064 21465 9092
rect 21039 9061 21051 9064
rect 20993 9055 21051 9061
rect 21453 9061 21465 9064
rect 21499 9092 21511 9095
rect 21499 9064 23336 9092
rect 21499 9061 21511 9064
rect 21453 9055 21511 9061
rect 20162 8984 20168 9036
rect 20220 9024 20226 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 20220 8996 20361 9024
rect 20220 8984 20226 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20772 8996 21281 9024
rect 20772 8984 20778 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 23106 8984 23112 9036
rect 23164 8984 23170 9036
rect 23308 9033 23336 9064
rect 23474 9052 23480 9104
rect 23532 9092 23538 9104
rect 25332 9092 25360 9132
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 27062 9120 27068 9172
rect 27120 9120 27126 9172
rect 27614 9120 27620 9172
rect 27672 9120 27678 9172
rect 23532 9064 25360 9092
rect 23532 9052 23538 9064
rect 23293 9027 23351 9033
rect 23293 8993 23305 9027
rect 23339 8993 23351 9027
rect 24397 9027 24455 9033
rect 24397 9024 24409 9027
rect 23293 8987 23351 8993
rect 23400 8996 24409 9024
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 20070 8916 20076 8968
rect 20128 8916 20134 8968
rect 20530 8916 20536 8968
rect 20588 8916 20594 8968
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21542 8956 21548 8968
rect 21131 8928 21548 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21821 8959 21879 8965
rect 21821 8956 21833 8959
rect 21692 8928 21833 8956
rect 21692 8916 21698 8928
rect 21821 8925 21833 8928
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 19904 8888 19932 8916
rect 20714 8888 20720 8900
rect 19904 8860 20720 8888
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 22020 8888 22048 8919
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22520 8928 22569 8956
rect 22520 8916 22526 8928
rect 22557 8925 22569 8928
rect 22603 8925 22615 8959
rect 23124 8956 23152 8984
rect 23400 8956 23428 8996
rect 24397 8993 24409 8996
rect 24443 8993 24455 9027
rect 24397 8987 24455 8993
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 25409 9027 25467 9033
rect 25409 9024 25421 9027
rect 24912 8996 25421 9024
rect 24912 8984 24918 8996
rect 25409 8993 25421 8996
rect 25455 8993 25467 9027
rect 25409 8987 25467 8993
rect 26973 9027 27031 9033
rect 26973 8993 26985 9027
rect 27019 9024 27031 9027
rect 27080 9024 27108 9120
rect 27019 8996 27108 9024
rect 27632 9024 27660 9120
rect 27709 9027 27767 9033
rect 27709 9024 27721 9027
rect 27632 8996 27721 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 27709 8993 27721 8996
rect 27755 8993 27767 9027
rect 27709 8987 27767 8993
rect 23124 8928 23428 8956
rect 22557 8919 22615 8925
rect 23474 8916 23480 8968
rect 23532 8916 23538 8968
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 24228 8888 24256 8919
rect 24578 8916 24584 8968
rect 24636 8916 24642 8968
rect 24762 8916 24768 8968
rect 24820 8956 24826 8968
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 24820 8928 25145 8956
rect 24820 8916 24826 8928
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 27614 8956 27620 8968
rect 27203 8928 27620 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 27614 8916 27620 8928
rect 27672 8916 27678 8968
rect 27798 8916 27804 8968
rect 27856 8916 27862 8968
rect 27893 8959 27951 8965
rect 27893 8925 27905 8959
rect 27939 8925 27951 8959
rect 27893 8919 27951 8925
rect 21048 8860 22048 8888
rect 22572 8860 24256 8888
rect 21048 8848 21054 8860
rect 22572 8832 22600 8860
rect 24394 8848 24400 8900
rect 24452 8888 24458 8900
rect 24854 8888 24860 8900
rect 24452 8860 24860 8888
rect 24452 8848 24458 8860
rect 24854 8848 24860 8860
rect 24912 8888 24918 8900
rect 25676 8891 25734 8897
rect 24912 8860 25176 8888
rect 24912 8848 24918 8860
rect 22002 8820 22008 8832
rect 19812 8792 22008 8820
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22554 8780 22560 8832
rect 22612 8780 22618 8832
rect 23014 8780 23020 8832
rect 23072 8820 23078 8832
rect 23201 8823 23259 8829
rect 23201 8820 23213 8823
rect 23072 8792 23213 8820
rect 23072 8780 23078 8792
rect 23201 8789 23213 8792
rect 23247 8789 23259 8823
rect 23201 8783 23259 8789
rect 25038 8780 25044 8832
rect 25096 8780 25102 8832
rect 25148 8820 25176 8860
rect 25676 8857 25688 8891
rect 25722 8888 25734 8891
rect 27816 8888 27844 8916
rect 25722 8860 27844 8888
rect 25722 8857 25734 8860
rect 25676 8851 25734 8857
rect 26789 8823 26847 8829
rect 26789 8820 26801 8823
rect 25148 8792 26801 8820
rect 26789 8789 26801 8792
rect 26835 8789 26847 8823
rect 26789 8783 26847 8789
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 27908 8820 27936 8919
rect 26936 8792 27936 8820
rect 26936 8780 26942 8792
rect 28350 8780 28356 8832
rect 28408 8780 28414 8832
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 1762 8616 1768 8628
rect 1719 8588 1768 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 1854 8576 1860 8628
rect 1912 8576 1918 8628
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8585 2191 8619
rect 2133 8579 2191 8585
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2455 8588 2774 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 1596 8489 1624 8576
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1872 8480 1900 8576
rect 2148 8548 2176 8579
rect 2746 8548 2774 8588
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4709 8619 4767 8625
rect 4709 8616 4721 8619
rect 4212 8588 4721 8616
rect 4212 8576 4218 8588
rect 4709 8585 4721 8588
rect 4755 8585 4767 8619
rect 4709 8579 4767 8585
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 2148 8520 2636 8548
rect 2746 8520 4108 8548
rect 2608 8489 2636 8520
rect 4080 8489 4108 8520
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4525 8551 4583 8557
rect 4525 8548 4537 8551
rect 4304 8520 4537 8548
rect 4304 8508 4310 8520
rect 4525 8517 4537 8520
rect 4571 8517 4583 8551
rect 5644 8548 5672 8579
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7524 8588 8033 8616
rect 7524 8576 7530 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 10870 8576 10876 8628
rect 10928 8576 10934 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 11112 8588 11161 8616
rect 11112 8576 11118 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 11698 8616 11704 8628
rect 11655 8588 11704 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11793 8619 11851 8625
rect 11793 8585 11805 8619
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 4525 8511 4583 8517
rect 5092 8520 5672 8548
rect 5727 8520 6040 8548
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1872 8452 2053 8480
rect 1581 8443 1639 8449
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2685 8443 2743 8449
rect 2884 8452 3157 8480
rect 2332 8412 2360 8443
rect 2700 8412 2728 8443
rect 2774 8412 2780 8424
rect 2332 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2884 8344 2912 8452
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 5092 8489 5120 8520
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4396 8452 4629 8480
rect 4396 8440 4402 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5727 8480 5755 8520
rect 6012 8489 6040 8520
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 7064 8520 7389 8548
rect 7064 8508 7070 8520
rect 7377 8517 7389 8520
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 7708 8520 8248 8548
rect 7708 8508 7714 8520
rect 8220 8489 8248 8520
rect 8956 8520 9444 8548
rect 8956 8492 8984 8520
rect 5399 8452 5755 8480
rect 5813 8483 5871 8489
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6135 8452 6653 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8938 8480 8944 8492
rect 8343 8452 8944 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 2958 8372 2964 8424
rect 3016 8372 3022 8424
rect 3878 8372 3884 8424
rect 3936 8372 3942 8424
rect 4632 8412 4660 8443
rect 5828 8412 5856 8443
rect 4632 8384 5856 8412
rect 1903 8316 2912 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 5810 8344 5816 8356
rect 3660 8316 5816 8344
rect 3660 8304 3666 8316
rect 5810 8304 5816 8316
rect 5868 8344 5874 8356
rect 6012 8344 6040 8443
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 5868 8316 6040 8344
rect 5868 8304 5874 8316
rect 6362 8304 6368 8356
rect 6420 8304 6426 8356
rect 6472 8344 6500 8375
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7558 8372 7564 8424
rect 7616 8372 7622 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8527 8384 9137 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 8570 8344 8576 8356
rect 6472 8316 8576 8344
rect 8570 8304 8576 8316
rect 8628 8344 8634 8356
rect 8665 8347 8723 8353
rect 8665 8344 8677 8347
rect 8628 8316 8677 8344
rect 8628 8304 8634 8316
rect 8665 8313 8677 8316
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 9306 8304 9312 8356
rect 9364 8304 9370 8356
rect 9416 8344 9444 8520
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 9732 8520 9781 8548
rect 9732 8508 9738 8520
rect 9769 8517 9781 8520
rect 9815 8517 9827 8551
rect 9769 8511 9827 8517
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 11808 8548 11836 8579
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 16482 8616 16488 8628
rect 14332 8588 16488 8616
rect 14332 8576 14338 8588
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 17957 8619 18015 8625
rect 17957 8585 17969 8619
rect 18003 8616 18015 8619
rect 18690 8616 18696 8628
rect 18003 8588 18696 8616
rect 18003 8585 18015 8588
rect 17957 8579 18015 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 20441 8619 20499 8625
rect 19760 8588 20300 8616
rect 19760 8576 19766 8588
rect 10376 8520 10824 8548
rect 10376 8508 10382 8520
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 10796 8489 10824 8520
rect 11348 8520 11836 8548
rect 12084 8520 18184 8548
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 10962 8480 10968 8492
rect 10827 8452 10968 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11348 8489 11376 8520
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11563 8452 11989 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10502 8412 10508 8424
rect 9723 8384 10508 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10686 8372 10692 8424
rect 10744 8372 10750 8424
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11532 8412 11560 8443
rect 11204 8384 11560 8412
rect 12084 8412 12112 8520
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12986 8480 12992 8492
rect 12216 8452 12992 8480
rect 12216 8440 12222 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14148 8452 14933 8480
rect 14148 8440 14154 8452
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15396 8489 15424 8520
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 12084 8384 12265 8412
rect 11204 8372 11210 8384
rect 12253 8381 12265 8384
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 13081 8415 13139 8421
rect 13081 8412 13093 8415
rect 12483 8384 13093 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13081 8381 13093 8384
rect 13127 8381 13139 8415
rect 13081 8375 13139 8381
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 16209 8415 16267 8421
rect 16209 8412 16221 8415
rect 15611 8384 16221 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 16209 8381 16221 8384
rect 16255 8381 16267 8415
rect 16776 8412 16804 8443
rect 17034 8440 17040 8492
rect 17092 8440 17098 8492
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17770 8480 17776 8492
rect 17359 8452 17776 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17920 8452 18061 8480
rect 17920 8440 17926 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18156 8480 18184 8520
rect 18230 8508 18236 8560
rect 18288 8548 18294 8560
rect 19153 8551 19211 8557
rect 19153 8548 19165 8551
rect 18288 8520 19165 8548
rect 18288 8508 18294 8520
rect 19153 8517 19165 8520
rect 19199 8548 19211 8551
rect 19334 8548 19340 8560
rect 19199 8520 19340 8548
rect 19199 8517 19211 8520
rect 19153 8511 19211 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19426 8508 19432 8560
rect 19484 8548 19490 8560
rect 19978 8548 19984 8560
rect 19484 8520 19984 8548
rect 19484 8508 19490 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 20070 8508 20076 8560
rect 20128 8508 20134 8560
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18156 8452 18429 8480
rect 18049 8443 18107 8449
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 20088 8480 20116 8508
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 20088 8452 20177 8480
rect 18417 8443 18475 8449
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20272 8480 20300 8588
rect 20441 8585 20453 8619
rect 20487 8616 20499 8619
rect 20530 8616 20536 8628
rect 20487 8588 20536 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20990 8576 20996 8628
rect 21048 8576 21054 8628
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21315 8588 22094 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 20714 8508 20720 8560
rect 20772 8508 20778 8560
rect 22066 8548 22094 8588
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 22244 8588 22477 8616
rect 22244 8576 22250 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 22554 8576 22560 8628
rect 22612 8576 22618 8628
rect 22649 8619 22707 8625
rect 22649 8585 22661 8619
rect 22695 8616 22707 8619
rect 23474 8616 23480 8628
rect 22695 8588 23480 8616
rect 22695 8585 22707 8588
rect 22649 8579 22707 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 23845 8619 23903 8625
rect 23845 8585 23857 8619
rect 23891 8616 23903 8619
rect 24578 8616 24584 8628
rect 23891 8588 24584 8616
rect 23891 8585 23903 8588
rect 23845 8579 23903 8585
rect 24578 8576 24584 8588
rect 24636 8576 24642 8628
rect 26326 8576 26332 8628
rect 26384 8576 26390 8628
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28445 8619 28503 8625
rect 28445 8616 28457 8619
rect 28408 8588 28457 8616
rect 28408 8576 28414 8588
rect 28445 8585 28457 8588
rect 28491 8585 28503 8619
rect 28445 8579 28503 8585
rect 22572 8548 22600 8576
rect 23934 8548 23940 8560
rect 21008 8520 21864 8548
rect 22066 8520 22600 8548
rect 22664 8520 23940 8548
rect 20625 8483 20683 8489
rect 20625 8480 20637 8483
rect 20272 8452 20637 8480
rect 20165 8443 20223 8449
rect 20625 8449 20637 8452
rect 20671 8449 20683 8483
rect 20732 8480 20760 8508
rect 21008 8492 21036 8520
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20732 8452 20913 8480
rect 20625 8443 20683 8449
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 20990 8440 20996 8492
rect 21048 8440 21054 8492
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 17402 8412 17408 8424
rect 16776 8384 17408 8412
rect 16209 8375 16267 8381
rect 12268 8344 12296 8375
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17543 8384 18153 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8412 18659 8415
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 18647 8384 20269 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 21192 8412 21220 8443
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 21836 8421 21864 8520
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 22462 8440 22468 8492
rect 22520 8480 22526 8492
rect 22557 8483 22615 8489
rect 22557 8480 22569 8483
rect 22520 8452 22569 8480
rect 22520 8440 22526 8452
rect 22557 8449 22569 8452
rect 22603 8480 22615 8483
rect 22664 8480 22692 8520
rect 22603 8452 22692 8480
rect 22603 8449 22615 8452
rect 22557 8443 22615 8449
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 23768 8489 23796 8520
rect 23934 8508 23940 8520
rect 23992 8508 23998 8560
rect 24762 8508 24768 8560
rect 24820 8508 24826 8560
rect 24854 8508 24860 8560
rect 24912 8508 24918 8560
rect 25038 8508 25044 8560
rect 25096 8548 25102 8560
rect 25096 8520 26096 8548
rect 25096 8508 25102 8520
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22796 8452 23029 8480
rect 22796 8440 22802 8452
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24780 8480 24808 8508
rect 24268 8452 24808 8480
rect 24268 8440 24274 8452
rect 20257 8375 20315 8381
rect 20732 8384 21220 8412
rect 21821 8415 21879 8421
rect 9416 8316 12296 8344
rect 15197 8347 15255 8353
rect 15197 8313 15209 8347
rect 15243 8344 15255 8347
rect 15654 8344 15660 8356
rect 15243 8316 15660 8344
rect 15243 8313 15255 8316
rect 15197 8307 15255 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 20732 8353 20760 8384
rect 21821 8381 21833 8415
rect 21867 8412 21879 8415
rect 22922 8412 22928 8424
rect 21867 8384 22928 8412
rect 21867 8381 21879 8384
rect 21821 8375 21879 8381
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 23198 8372 23204 8424
rect 23256 8372 23262 8424
rect 24394 8372 24400 8424
rect 24452 8372 24458 8424
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 24872 8412 24900 8508
rect 26068 8489 26096 8520
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 26237 8483 26295 8489
rect 26237 8449 26249 8483
rect 26283 8480 26295 8483
rect 26344 8480 26372 8576
rect 26283 8452 26372 8480
rect 26283 8449 26295 8452
rect 26237 8443 26295 8449
rect 26970 8440 26976 8492
rect 27028 8440 27034 8492
rect 27065 8483 27123 8489
rect 27065 8449 27077 8483
rect 27111 8480 27123 8483
rect 28368 8480 28396 8576
rect 27111 8452 28396 8480
rect 27111 8449 27123 8452
rect 27065 8443 27123 8449
rect 25317 8415 25375 8421
rect 25317 8412 25329 8415
rect 24872 8384 25329 8412
rect 25317 8381 25329 8384
rect 25363 8381 25375 8415
rect 25317 8375 25375 8381
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 26878 8412 26884 8424
rect 25884 8384 26884 8412
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 20717 8347 20775 8353
rect 16899 8316 20668 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 3050 8276 3056 8288
rect 2823 8248 3056 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5132 8248 5457 8276
rect 5132 8236 5138 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 6380 8276 6408 8304
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6380 8248 6837 8276
rect 5445 8239 5503 8245
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 10226 8276 10232 8288
rect 7340 8248 10232 8276
rect 7340 8236 7346 8248
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 12710 8236 12716 8288
rect 12768 8236 12774 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 14737 8279 14795 8285
rect 14737 8276 14749 8279
rect 14700 8248 14749 8276
rect 14700 8236 14706 8248
rect 14737 8245 14749 8248
rect 14783 8245 14795 8279
rect 14737 8239 14795 8245
rect 15838 8236 15844 8288
rect 15896 8236 15902 8288
rect 17129 8279 17187 8285
rect 17129 8245 17141 8279
rect 17175 8276 17187 8279
rect 17862 8276 17868 8288
rect 17175 8248 17868 8276
rect 17175 8245 17187 8248
rect 17129 8239 17187 8245
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 19058 8236 19064 8288
rect 19116 8236 19122 8288
rect 20640 8276 20668 8316
rect 20717 8313 20729 8347
rect 20763 8313 20775 8347
rect 23382 8344 23388 8356
rect 20717 8307 20775 8313
rect 21376 8316 23388 8344
rect 21376 8276 21404 8316
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 23566 8304 23572 8356
rect 23624 8304 23630 8356
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8344 24087 8347
rect 25792 8344 25820 8372
rect 24075 8316 25820 8344
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 20640 8248 21404 8276
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 22462 8276 22468 8288
rect 21508 8248 22468 8276
rect 21508 8236 21514 8248
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 22646 8236 22652 8288
rect 22704 8276 22710 8288
rect 25884 8276 25912 8384
rect 26878 8372 26884 8384
rect 26936 8372 26942 8424
rect 26988 8412 27016 8440
rect 27249 8415 27307 8421
rect 27249 8412 27261 8415
rect 26988 8384 27261 8412
rect 27249 8381 27261 8384
rect 27295 8381 27307 8415
rect 27249 8375 27307 8381
rect 27801 8415 27859 8421
rect 27801 8381 27813 8415
rect 27847 8412 27859 8415
rect 27890 8412 27896 8424
rect 27847 8384 27896 8412
rect 27847 8381 27859 8384
rect 27801 8375 27859 8381
rect 27890 8372 27896 8384
rect 27948 8372 27954 8424
rect 27982 8372 27988 8424
rect 28040 8372 28046 8424
rect 22704 8248 25912 8276
rect 22704 8236 22710 8248
rect 25958 8236 25964 8288
rect 26016 8236 26022 8288
rect 26142 8236 26148 8288
rect 26200 8276 26206 8288
rect 26421 8279 26479 8285
rect 26421 8276 26433 8279
rect 26200 8248 26433 8276
rect 26200 8236 26206 8248
rect 26421 8245 26433 8248
rect 26467 8245 26479 8279
rect 26421 8239 26479 8245
rect 27522 8236 27528 8288
rect 27580 8236 27586 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3602 8072 3608 8084
rect 2832 8044 3608 8072
rect 2832 8032 2838 8044
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4304 8044 4997 8072
rect 4304 8032 4310 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 10042 8072 10048 8084
rect 4985 8035 5043 8041
rect 5828 8044 10048 8072
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 5828 8004 5856 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 12710 8032 12716 8084
rect 12768 8032 12774 8084
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8072 14243 8075
rect 14550 8072 14556 8084
rect 14231 8044 14556 8072
rect 14231 8041 14243 8044
rect 14185 8035 14243 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 18782 8072 18788 8084
rect 16816 8044 18788 8072
rect 16816 8032 16822 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 19058 8032 19064 8084
rect 19116 8072 19122 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19116 8044 19625 8072
rect 19116 8032 19122 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 20070 8032 20076 8084
rect 20128 8032 20134 8084
rect 20622 8072 20628 8084
rect 20272 8044 20628 8072
rect 7006 8004 7012 8016
rect 4948 7976 5856 8004
rect 5920 7976 7012 8004
rect 4948 7964 4954 7976
rect 4801 7939 4859 7945
rect 3896 7908 4752 7936
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 2746 7840 3372 7868
rect 1664 7803 1722 7809
rect 1664 7769 1676 7803
rect 1710 7800 1722 7803
rect 2746 7800 2774 7840
rect 1710 7772 2774 7800
rect 1710 7769 1722 7772
rect 1664 7763 1722 7769
rect 3234 7760 3240 7812
rect 3292 7760 3298 7812
rect 3344 7800 3372 7840
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 3896 7877 3924 7908
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3844 7840 3893 7868
rect 3844 7828 3850 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 4724 7868 4752 7908
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5074 7936 5080 7948
rect 4847 7908 5080 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5920 7945 5948 7976
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 9582 8004 9588 8016
rect 7432 7976 9588 8004
rect 7432 7964 7438 7976
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 8128 7945 8156 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6052 7908 6837 7936
rect 6052 7896 6058 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7936 8355 7939
rect 9306 7936 9312 7948
rect 8343 7908 9312 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11020 7908 11621 7936
rect 11020 7896 11026 7908
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11940 7908 12081 7936
rect 11940 7896 11946 7908
rect 12069 7905 12081 7908
rect 12115 7936 12127 7939
rect 12728 7936 12756 8032
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12115 7908 12388 7936
rect 12728 7908 12817 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 4724 7840 5549 7868
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 4525 7803 4583 7809
rect 4525 7800 4537 7803
rect 3344 7772 4537 7800
rect 4525 7769 4537 7772
rect 4571 7769 4583 7803
rect 5552 7800 5580 7831
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6420 7840 6561 7868
rect 6420 7828 6426 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6730 7868 6736 7880
rect 6687 7840 6736 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7098 7800 7104 7812
rect 5552 7772 7104 7800
rect 4525 7763 4583 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 7484 7800 7512 7831
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8628 7840 8769 7868
rect 8628 7828 8634 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 9171 7840 9720 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9582 7800 9588 7812
rect 7484 7772 9588 7800
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 9692 7800 9720 7840
rect 9766 7830 9772 7882
rect 9824 7877 9830 7882
rect 9824 7868 9834 7877
rect 9824 7840 9867 7868
rect 9824 7831 9834 7840
rect 9824 7830 9830 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11204 7840 11437 7868
rect 11204 7828 11210 7840
rect 11425 7837 11437 7840
rect 11471 7868 11483 7871
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11471 7840 11529 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12360 7868 12388 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13035 7908 13645 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 15856 7936 15884 8032
rect 17681 8007 17739 8013
rect 16040 7976 17448 8004
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 13780 7908 15516 7936
rect 15856 7908 15945 7936
rect 13780 7896 13786 7908
rect 12360 7840 13492 7868
rect 10036 7803 10094 7809
rect 9692 7772 9996 7800
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7732 3571 7735
rect 4338 7732 4344 7744
rect 3559 7704 4344 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 4338 7692 4344 7704
rect 4396 7732 4402 7744
rect 5166 7732 5172 7744
rect 4396 7704 5172 7732
rect 4396 7692 4402 7704
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 5626 7692 5632 7744
rect 5684 7692 5690 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 7282 7732 7288 7744
rect 5960 7704 7288 7732
rect 5960 7692 5966 7704
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7524 7704 8033 7732
rect 7524 7692 7530 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9088 7704 9689 7732
rect 9088 7692 9094 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9968 7732 9996 7772
rect 10036 7769 10048 7803
rect 10082 7800 10094 7803
rect 12434 7800 12440 7812
rect 10082 7772 12440 7800
rect 10082 7769 10094 7772
rect 10036 7763 10094 7769
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 13464 7800 13492 7840
rect 13538 7828 13544 7880
rect 13596 7828 13602 7880
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14274 7868 14280 7880
rect 14056 7840 14280 7868
rect 14056 7828 14062 7840
rect 14274 7828 14280 7840
rect 14332 7868 14338 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 14332 7840 14381 7868
rect 14332 7828 14338 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14608 7840 14657 7868
rect 14608 7828 14614 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7837 15255 7871
rect 15197 7831 15255 7837
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15488 7868 15516 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 16040 7868 16068 7976
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 16163 7908 16773 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 15488 7840 16068 7868
rect 15381 7831 15439 7837
rect 15212 7800 15240 7831
rect 13464 7772 15240 7800
rect 15396 7800 15424 7831
rect 16206 7828 16212 7880
rect 16264 7868 16270 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 16264 7840 16681 7868
rect 16264 7828 16270 7840
rect 16669 7837 16681 7840
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17420 7877 17448 7976
rect 17681 7973 17693 8007
rect 17727 7973 17739 8007
rect 17681 7967 17739 7973
rect 17696 7936 17724 7967
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 20088 8004 20116 8032
rect 17920 7976 20116 8004
rect 17920 7964 17926 7976
rect 18417 7939 18475 7945
rect 17696 7908 18184 7936
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18156 7877 18184 7908
rect 18417 7905 18429 7939
rect 18463 7936 18475 7939
rect 19058 7936 19064 7948
rect 18463 7908 19064 7936
rect 18463 7905 18475 7908
rect 18417 7899 18475 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 20070 7936 20076 7948
rect 19291 7908 20076 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17828 7840 17877 7868
rect 17828 7828 17834 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 17880 7800 17908 7831
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 19702 7868 19708 7880
rect 19475 7840 19708 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 18230 7800 18236 7812
rect 15396 7772 16988 7800
rect 17880 7772 18236 7800
rect 11146 7732 11152 7744
rect 9968 7704 11152 7732
rect 9677 7695 9735 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11238 7692 11244 7744
rect 11296 7692 11302 7744
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 13449 7735 13507 7741
rect 13449 7732 13461 7735
rect 13228 7704 13461 7732
rect 13228 7692 13234 7704
rect 13449 7701 13461 7704
rect 13495 7701 13507 7735
rect 13449 7695 13507 7701
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15194 7732 15200 7744
rect 15151 7704 15200 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16960 7741 16988 7772
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 20272 7800 20300 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 20714 8032 20720 8084
rect 20772 8032 20778 8084
rect 21545 8075 21603 8081
rect 21545 8041 21557 8075
rect 21591 8072 21603 8075
rect 22002 8072 22008 8084
rect 21591 8044 22008 8072
rect 21591 8041 21603 8044
rect 21545 8035 21603 8041
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 23106 8072 23112 8084
rect 22888 8044 23112 8072
rect 22888 8032 22894 8044
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 23198 8032 23204 8084
rect 23256 8072 23262 8084
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 23256 8044 23489 8072
rect 23256 8032 23262 8044
rect 23477 8041 23489 8044
rect 23523 8041 23535 8075
rect 23477 8035 23535 8041
rect 24397 8075 24455 8081
rect 24397 8041 24409 8075
rect 24443 8072 24455 8075
rect 24578 8072 24584 8084
rect 24443 8044 24584 8072
rect 24443 8041 24455 8044
rect 24397 8035 24455 8041
rect 24578 8032 24584 8044
rect 24636 8032 24642 8084
rect 24762 8032 24768 8084
rect 24820 8032 24826 8084
rect 25314 8032 25320 8084
rect 25372 8072 25378 8084
rect 26142 8072 26148 8084
rect 25372 8044 26148 8072
rect 25372 8032 25378 8044
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 28132 8044 28273 8072
rect 28132 8032 28138 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 20732 8004 20760 8032
rect 20364 7976 21404 8004
rect 20364 7877 20392 7976
rect 20456 7908 21220 7936
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 18524 7772 20300 7800
rect 18524 7744 18552 7772
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 16172 7704 16589 7732
rect 16172 7692 16178 7704
rect 16577 7701 16589 7704
rect 16623 7701 16635 7735
rect 16577 7695 16635 7701
rect 16945 7735 17003 7741
rect 16945 7701 16957 7735
rect 16991 7701 17003 7735
rect 16945 7695 17003 7701
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17276 7704 17509 7732
rect 17276 7692 17282 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18414 7732 18420 7744
rect 18003 7704 18420 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18506 7692 18512 7744
rect 18564 7692 18570 7744
rect 19061 7735 19119 7741
rect 19061 7701 19073 7735
rect 19107 7732 19119 7735
rect 19518 7732 19524 7744
rect 19107 7704 19524 7732
rect 19107 7701 19119 7704
rect 19061 7695 19119 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 20165 7735 20223 7741
rect 20165 7701 20177 7735
rect 20211 7732 20223 7735
rect 20456 7732 20484 7908
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21192 7877 21220 7908
rect 21266 7896 21272 7948
rect 21324 7896 21330 7948
rect 21376 7936 21404 7976
rect 21450 7964 21456 8016
rect 21508 8004 21514 8016
rect 27157 8007 27215 8013
rect 21508 7976 24801 8004
rect 21508 7964 21514 7976
rect 22281 7939 22339 7945
rect 21376 7908 21956 7936
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7837 21235 7871
rect 21284 7868 21312 7896
rect 21928 7877 21956 7908
rect 22281 7905 22293 7939
rect 22327 7936 22339 7939
rect 23198 7936 23204 7948
rect 22327 7908 23204 7936
rect 22327 7905 22339 7908
rect 22281 7899 22339 7905
rect 23198 7896 23204 7908
rect 23256 7896 23262 7948
rect 24026 7936 24032 7948
rect 23308 7908 24032 7936
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 21284 7840 21465 7868
rect 21177 7831 21235 7837
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22186 7868 22192 7880
rect 22143 7840 22192 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 20533 7803 20591 7809
rect 20533 7769 20545 7803
rect 20579 7769 20591 7803
rect 21468 7800 21496 7831
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 23308 7864 23336 7908
rect 24026 7896 24032 7908
rect 24084 7936 24090 7948
rect 24210 7936 24216 7948
rect 24084 7908 24216 7936
rect 24084 7896 24090 7908
rect 24210 7896 24216 7908
rect 24268 7896 24274 7948
rect 23385 7871 23443 7877
rect 23385 7864 23397 7871
rect 23308 7837 23397 7864
rect 23431 7837 23443 7871
rect 23308 7836 23443 7837
rect 23385 7831 23443 7836
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 22848 7800 22876 7831
rect 21468 7772 22876 7800
rect 20533 7763 20591 7769
rect 20211 7704 20484 7732
rect 20548 7732 20576 7763
rect 20898 7732 20904 7744
rect 20548 7704 20904 7732
rect 20211 7701 20223 7704
rect 20165 7695 20223 7701
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 20990 7692 20996 7744
rect 21048 7692 21054 7744
rect 21174 7692 21180 7744
rect 21232 7732 21238 7744
rect 21729 7735 21787 7741
rect 21729 7732 21741 7735
rect 21232 7704 21741 7732
rect 21232 7692 21238 7704
rect 21729 7701 21741 7704
rect 21775 7701 21787 7735
rect 21729 7695 21787 7701
rect 22738 7692 22744 7744
rect 22796 7692 22802 7744
rect 22922 7692 22928 7744
rect 22980 7692 22986 7744
rect 23201 7735 23259 7741
rect 23201 7701 23213 7735
rect 23247 7732 23259 7735
rect 23676 7732 23704 7831
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24121 7871 24179 7877
rect 24121 7868 24133 7871
rect 23900 7840 24133 7868
rect 23900 7828 23906 7840
rect 24121 7837 24133 7840
rect 24167 7868 24179 7871
rect 24486 7868 24492 7880
rect 24167 7840 24492 7868
rect 24167 7837 24179 7840
rect 24121 7831 24179 7837
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 24596 7800 24624 7831
rect 23952 7772 24624 7800
rect 23952 7741 23980 7772
rect 23247 7704 23704 7732
rect 23937 7735 23995 7741
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 23937 7701 23949 7735
rect 23983 7701 23995 7735
rect 23937 7695 23995 7701
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24688 7732 24716 7831
rect 24773 7800 24801 7976
rect 27157 7973 27169 8007
rect 27203 8004 27215 8007
rect 27430 8004 27436 8016
rect 27203 7976 27436 8004
rect 27203 7973 27215 7976
rect 27157 7967 27215 7973
rect 27430 7964 27436 7976
rect 27488 8004 27494 8016
rect 27617 8007 27675 8013
rect 27617 8004 27629 8007
rect 27488 7976 27629 8004
rect 27488 7964 27494 7976
rect 27617 7973 27629 7976
rect 27663 7973 27675 8007
rect 27617 7967 27675 7973
rect 28166 7964 28172 8016
rect 28224 7964 28230 8016
rect 24946 7896 24952 7948
rect 25004 7896 25010 7948
rect 26510 7896 26516 7948
rect 26568 7896 26574 7948
rect 25216 7871 25274 7877
rect 25216 7837 25228 7871
rect 25262 7868 25274 7871
rect 25958 7868 25964 7880
rect 25262 7840 25964 7868
rect 25262 7837 25274 7840
rect 25216 7831 25274 7837
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 26694 7828 26700 7880
rect 26752 7828 26758 7880
rect 26786 7828 26792 7880
rect 26844 7868 26850 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 26844 7840 27261 7868
rect 26844 7828 26850 7840
rect 27249 7837 27261 7840
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 28077 7871 28135 7877
rect 28077 7837 28089 7871
rect 28123 7868 28135 7871
rect 28184 7868 28212 7964
rect 28123 7840 28212 7868
rect 28537 7871 28595 7877
rect 28123 7837 28135 7840
rect 28077 7831 28135 7837
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 28626 7868 28632 7880
rect 28583 7840 28632 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 27448 7800 27476 7831
rect 28626 7828 28632 7840
rect 28684 7828 28690 7880
rect 24773 7772 27476 7800
rect 24176 7704 24716 7732
rect 24176 7692 24182 7704
rect 26142 7692 26148 7744
rect 26200 7732 26206 7744
rect 26329 7735 26387 7741
rect 26329 7732 26341 7735
rect 26200 7704 26341 7732
rect 26200 7692 26206 7704
rect 26329 7701 26341 7704
rect 26375 7701 26387 7735
rect 26329 7695 26387 7701
rect 28350 7692 28356 7744
rect 28408 7692 28414 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 3510 7528 3516 7540
rect 1636 7500 3516 7528
rect 1636 7488 1642 7500
rect 2148 7469 2176 7500
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4672 7500 5089 7528
rect 4672 7488 4678 7500
rect 5077 7497 5089 7500
rect 5123 7528 5135 7531
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5123 7500 5825 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6144 7500 6377 7528
rect 6144 7488 6150 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 10594 7528 10600 7540
rect 6365 7491 6423 7497
rect 6748 7500 10600 7528
rect 2133 7463 2191 7469
rect 2133 7429 2145 7463
rect 2179 7460 2191 7463
rect 3786 7460 3792 7472
rect 2179 7432 2213 7460
rect 2516 7432 3792 7460
rect 2179 7429 2191 7432
rect 2133 7423 2191 7429
rect 2516 7401 2544 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 1627 7364 2513 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3605 7395 3663 7401
rect 2915 7364 3464 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 2792 7324 2820 7355
rect 2332 7296 2820 7324
rect 3053 7327 3111 7333
rect 2332 7265 2360 7296
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 2317 7259 2375 7265
rect 2317 7225 2329 7259
rect 2363 7225 2375 7259
rect 2317 7219 2375 7225
rect 2593 7259 2651 7265
rect 2593 7225 2605 7259
rect 2639 7256 2651 7259
rect 3068 7256 3096 7287
rect 2639 7228 3096 7256
rect 2639 7225 2651 7228
rect 2593 7219 2651 7225
rect 3436 7188 3464 7364
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 3651 7364 4108 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 3786 7284 3792 7336
rect 3844 7284 3850 7336
rect 4080 7324 4108 7364
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4212 7364 4629 7392
rect 4212 7352 4218 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5902 7392 5908 7404
rect 5215 7364 5908 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 4338 7324 4344 7336
rect 4080 7296 4344 7324
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 5000 7324 5028 7352
rect 4479 7296 5028 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5316 7296 5365 7324
rect 5316 7284 5322 7296
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 6012 7324 6040 7355
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6748 7401 6776 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 11238 7488 11244 7540
rect 11296 7488 11302 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 14642 7488 14648 7540
rect 14700 7488 14706 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15252 7500 15301 7528
rect 15252 7488 15258 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 7000 7463 7058 7469
rect 7000 7429 7012 7463
rect 7046 7460 7058 7463
rect 7466 7460 7472 7472
rect 7046 7432 7472 7460
rect 7046 7429 7058 7432
rect 7000 7423 7058 7429
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 9766 7460 9772 7472
rect 8220 7432 9772 7460
rect 8220 7401 8248 7432
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 9858 7420 9864 7472
rect 9916 7420 9922 7472
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 10781 7463 10839 7469
rect 10781 7460 10793 7463
rect 10744 7432 10793 7460
rect 10744 7420 10750 7432
rect 10781 7429 10793 7432
rect 10827 7429 10839 7463
rect 10781 7423 10839 7429
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6420 7364 6561 7392
rect 6420 7352 6426 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 8205 7395 8263 7401
rect 6733 7355 6791 7361
rect 6840 7364 7788 7392
rect 6840 7324 6868 7364
rect 6012 7296 6868 7324
rect 7760 7324 7788 7364
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8472 7395 8530 7401
rect 8472 7361 8484 7395
rect 8518 7392 8530 7395
rect 9030 7392 9036 7404
rect 8518 7364 9036 7392
rect 8518 7361 8530 7364
rect 8472 7355 8530 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9582 7352 9588 7404
rect 9640 7352 9646 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11256 7392 11284 7488
rect 13170 7460 13176 7472
rect 13096 7432 13176 7460
rect 11195 7364 11284 7392
rect 11517 7395 11575 7401
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 13096 7392 13124 7432
rect 13170 7420 13176 7432
rect 13228 7460 13234 7472
rect 13725 7463 13783 7469
rect 13725 7460 13737 7463
rect 13228 7432 13737 7460
rect 13228 7420 13234 7432
rect 13725 7429 13737 7432
rect 13771 7429 13783 7463
rect 13725 7423 13783 7429
rect 11563 7364 13124 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13504 7364 14013 7392
rect 13504 7352 13510 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14332 7364 14565 7392
rect 14332 7352 14338 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14660 7392 14688 7488
rect 15304 7460 15332 7491
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 16206 7528 16212 7540
rect 15804 7500 16212 7528
rect 15804 7488 15810 7500
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 17678 7528 17684 7540
rect 16899 7500 17684 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 18656 7500 19533 7528
rect 18656 7488 18662 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 19521 7491 19579 7497
rect 19702 7488 19708 7540
rect 19760 7488 19766 7540
rect 20254 7488 20260 7540
rect 20312 7528 20318 7540
rect 20312 7500 21128 7528
rect 20312 7488 20318 7500
rect 17310 7460 17316 7472
rect 15304 7432 15700 7460
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14660 7364 14841 7392
rect 14553 7355 14611 7361
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 15672 7401 15700 7432
rect 16960 7432 17316 7460
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 16960 7401 16988 7432
rect 17310 7420 17316 7432
rect 17368 7460 17374 7472
rect 19150 7460 19156 7472
rect 17368 7432 17724 7460
rect 17368 7420 17374 7432
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17083 7364 17417 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 8312 7324 8340 7352
rect 7760 7296 8340 7324
rect 5353 7287 5411 7293
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 3878 7256 3884 7268
rect 3559 7228 3884 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3878 7216 3884 7228
rect 3936 7256 3942 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3936 7228 3985 7256
rect 3936 7216 3942 7228
rect 3973 7225 3985 7228
rect 4019 7225 4031 7259
rect 4890 7256 4896 7268
rect 3973 7219 4031 7225
rect 4080 7228 4896 7256
rect 4080 7188 4108 7228
rect 4890 7216 4896 7228
rect 4948 7256 4954 7268
rect 6730 7256 6736 7268
rect 4948 7228 6736 7256
rect 4948 7216 4954 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 9600 7265 9628 7352
rect 17696 7336 17724 7432
rect 17788 7432 19156 7460
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 9585 7259 9643 7265
rect 9585 7225 9597 7259
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 3436 7160 4108 7188
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 6914 7188 6920 7200
rect 6135 7160 6920 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 8110 7188 8116 7200
rect 7156 7160 8116 7188
rect 7156 7148 7162 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9784 7188 9812 7287
rect 10965 7259 11023 7265
rect 10965 7225 10977 7259
rect 11011 7256 11023 7259
rect 11716 7256 11744 7287
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12124 7296 12357 7324
rect 12124 7284 12130 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 11011 7228 11744 7256
rect 11011 7225 11023 7228
rect 10965 7219 11023 7225
rect 11146 7188 11152 7200
rect 9784 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7188 11210 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11204 7160 11897 7188
rect 11204 7148 11210 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 12360 7188 12388 7287
rect 12526 7284 12532 7336
rect 12584 7284 12590 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7324 13047 7327
rect 13078 7324 13084 7336
rect 13035 7296 13084 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7293 13323 7327
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 13265 7287 13323 7293
rect 13924 7296 14657 7324
rect 13280 7256 13308 7287
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 13280 7228 13829 7256
rect 13817 7225 13829 7228
rect 13863 7225 13875 7259
rect 13817 7219 13875 7225
rect 13924 7188 13952 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7293 15899 7327
rect 15841 7287 15899 7293
rect 15381 7259 15439 7265
rect 15381 7225 15393 7259
rect 15427 7256 15439 7259
rect 15856 7256 15884 7287
rect 17126 7284 17132 7336
rect 17184 7284 17190 7336
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 17678 7284 17684 7336
rect 17736 7284 17742 7336
rect 17144 7256 17172 7284
rect 15427 7228 15884 7256
rect 15948 7228 17172 7256
rect 15427 7225 15439 7228
rect 15381 7219 15439 7225
rect 12360 7160 13952 7188
rect 14369 7191 14427 7197
rect 11885 7151 11943 7157
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 15948 7188 15976 7228
rect 14415 7160 15976 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 16114 7148 16120 7200
rect 16172 7148 16178 7200
rect 17236 7188 17264 7284
rect 17310 7216 17316 7268
rect 17368 7256 17374 7268
rect 17788 7256 17816 7432
rect 19150 7420 19156 7432
rect 19208 7420 19214 7472
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 21100 7469 21128 7500
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21416 7500 21487 7528
rect 21416 7488 21422 7500
rect 20349 7463 20407 7469
rect 20349 7460 20361 7463
rect 19392 7432 20361 7460
rect 19392 7420 19398 7432
rect 20349 7429 20361 7432
rect 20395 7429 20407 7463
rect 20349 7423 20407 7429
rect 21085 7463 21143 7469
rect 21085 7429 21097 7463
rect 21131 7429 21143 7463
rect 21085 7423 21143 7429
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 18414 7352 18420 7404
rect 18472 7392 18478 7404
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18472 7364 18889 7392
rect 18472 7352 18478 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19475 7364 19748 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7324 18015 7327
rect 18506 7324 18512 7336
rect 18003 7296 18512 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 17368 7228 17816 7256
rect 17865 7259 17923 7265
rect 17368 7216 17374 7228
rect 17865 7225 17877 7259
rect 17911 7256 17923 7259
rect 18325 7259 18383 7265
rect 18325 7256 18337 7259
rect 17911 7228 18337 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 18325 7225 18337 7228
rect 18371 7256 18383 7259
rect 18708 7256 18736 7287
rect 19720 7268 19748 7364
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 20070 7352 20076 7404
rect 20128 7352 20134 7404
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 21192 7392 21220 7488
rect 20303 7364 21220 7392
rect 21284 7392 21312 7488
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 21284 7364 21373 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 20088 7324 20116 7352
rect 21459 7324 21487 7500
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22244 7500 22477 7528
rect 22244 7488 22250 7500
rect 22465 7497 22477 7500
rect 22511 7497 22523 7531
rect 22646 7528 22652 7540
rect 22465 7491 22523 7497
rect 22572 7500 22652 7528
rect 21634 7420 21640 7472
rect 21692 7460 21698 7472
rect 22572 7460 22600 7500
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 22796 7500 23213 7528
rect 22796 7488 22802 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23201 7491 23259 7497
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 23842 7528 23848 7540
rect 23532 7500 23848 7528
rect 23532 7488 23538 7500
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 24486 7488 24492 7540
rect 24544 7528 24550 7540
rect 25501 7531 25559 7537
rect 24544 7500 25452 7528
rect 24544 7488 24550 7500
rect 25424 7460 25452 7500
rect 25501 7497 25513 7531
rect 25547 7528 25559 7531
rect 25547 7500 25728 7528
rect 25547 7497 25559 7500
rect 25501 7491 25559 7497
rect 25700 7460 25728 7500
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 25832 7500 28212 7528
rect 25832 7488 25838 7500
rect 21692 7432 22600 7460
rect 22664 7432 24992 7460
rect 25424 7432 25636 7460
rect 25700 7432 27200 7460
rect 21692 7420 21698 7432
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 20088 7296 21833 7324
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22005 7327 22063 7333
rect 22005 7293 22017 7327
rect 22051 7293 22063 7327
rect 22005 7287 22063 7293
rect 18371 7228 18736 7256
rect 19337 7259 19395 7265
rect 18371 7225 18383 7228
rect 18325 7219 18383 7225
rect 19337 7225 19349 7259
rect 19383 7256 19395 7259
rect 19518 7256 19524 7268
rect 19383 7228 19524 7256
rect 19383 7225 19395 7228
rect 19337 7219 19395 7225
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 19702 7216 19708 7268
rect 19760 7216 19766 7268
rect 20073 7259 20131 7265
rect 20073 7225 20085 7259
rect 20119 7256 20131 7259
rect 22020 7256 22048 7287
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 20119 7228 22048 7256
rect 20119 7225 20131 7228
rect 20073 7219 20131 7225
rect 21082 7188 21088 7200
rect 17236 7160 21088 7188
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 21542 7148 21548 7200
rect 21600 7188 21606 7200
rect 22664 7188 22692 7432
rect 23474 7352 23480 7404
rect 23532 7352 23538 7404
rect 24964 7392 24992 7432
rect 25608 7392 25636 7432
rect 25682 7392 25688 7404
rect 24964 7364 25544 7392
rect 25608 7364 25688 7392
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 23382 7324 23388 7336
rect 22787 7296 23388 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 23382 7284 23388 7296
rect 23440 7284 23446 7336
rect 23569 7327 23627 7333
rect 23569 7293 23581 7327
rect 23615 7293 23627 7327
rect 23569 7287 23627 7293
rect 23753 7327 23811 7333
rect 23753 7293 23765 7327
rect 23799 7293 23811 7327
rect 23753 7287 23811 7293
rect 21600 7160 22692 7188
rect 21600 7148 21606 7160
rect 23290 7148 23296 7200
rect 23348 7148 23354 7200
rect 23584 7188 23612 7287
rect 23768 7256 23796 7287
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 25406 7324 25412 7336
rect 24268 7296 25412 7324
rect 24268 7284 24274 7296
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25516 7324 25544 7364
rect 25682 7352 25688 7364
rect 25740 7352 25746 7404
rect 25774 7352 25780 7404
rect 25832 7392 25838 7404
rect 25961 7395 26019 7401
rect 25961 7392 25973 7395
rect 25832 7364 25973 7392
rect 25832 7352 25838 7364
rect 25961 7361 25973 7364
rect 26007 7361 26019 7395
rect 25961 7355 26019 7361
rect 26142 7352 26148 7404
rect 26200 7352 26206 7404
rect 27172 7401 27200 7432
rect 27157 7395 27215 7401
rect 27157 7361 27169 7395
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27430 7352 27436 7404
rect 27488 7352 27494 7404
rect 28184 7401 28212 7500
rect 28169 7395 28227 7401
rect 28169 7361 28181 7395
rect 28215 7361 28227 7395
rect 28169 7355 28227 7361
rect 27617 7327 27675 7333
rect 27617 7324 27629 7327
rect 25516 7296 27629 7324
rect 27617 7293 27629 7296
rect 27663 7293 27675 7327
rect 27617 7287 27675 7293
rect 26973 7259 27031 7265
rect 26973 7256 26985 7259
rect 23768 7228 26985 7256
rect 26973 7225 26985 7228
rect 27019 7225 27031 7259
rect 26973 7219 27031 7225
rect 25314 7188 25320 7200
rect 23584 7160 25320 7188
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 25777 7191 25835 7197
rect 25777 7157 25789 7191
rect 25823 7188 25835 7191
rect 25866 7188 25872 7200
rect 25823 7160 25872 7188
rect 25823 7157 25835 7160
rect 25777 7151 25835 7157
rect 25866 7148 25872 7160
rect 25924 7148 25930 7200
rect 26050 7148 26056 7200
rect 26108 7188 26114 7200
rect 26697 7191 26755 7197
rect 26697 7188 26709 7191
rect 26108 7160 26709 7188
rect 26108 7148 26114 7160
rect 26697 7157 26709 7160
rect 26743 7157 26755 7191
rect 26697 7151 26755 7157
rect 27890 7148 27896 7200
rect 27948 7148 27954 7200
rect 28258 7148 28264 7200
rect 28316 7148 28322 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3844 6956 3893 6984
rect 3844 6944 3850 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 4154 6944 4160 6996
rect 4212 6944 4218 6996
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5258 6984 5264 6996
rect 5215 6956 5264 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5368 6956 6408 6984
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 5368 6916 5396 6956
rect 4396 6888 5396 6916
rect 6380 6916 6408 6956
rect 6822 6944 6828 6996
rect 6880 6944 6886 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7064 6956 7389 6984
rect 7064 6944 7070 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 8294 6944 8300 6996
rect 8352 6944 8358 6996
rect 9858 6944 9864 6996
rect 9916 6944 9922 6996
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 12250 6984 12256 6996
rect 11563 6956 12256 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12434 6944 12440 6996
rect 12492 6944 12498 6996
rect 13078 6944 13084 6996
rect 13136 6944 13142 6996
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14608 6956 14749 6984
rect 14608 6944 14614 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 14737 6947 14795 6953
rect 15562 6944 15568 6996
rect 15620 6944 15626 6996
rect 15930 6944 15936 6996
rect 15988 6944 15994 6996
rect 16022 6944 16028 6996
rect 16080 6944 16086 6996
rect 17313 6987 17371 6993
rect 17313 6953 17325 6987
rect 17359 6984 17371 6987
rect 18138 6984 18144 6996
rect 17359 6956 18144 6984
rect 17359 6953 17371 6956
rect 17313 6947 17371 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 19886 6984 19892 6996
rect 18923 6956 19892 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 21542 6984 21548 6996
rect 20732 6956 21548 6984
rect 8312 6916 8340 6944
rect 6380 6888 8340 6916
rect 10428 6888 11928 6916
rect 4396 6876 4402 6888
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3878 6848 3884 6860
rect 3292 6820 3884 6848
rect 3292 6808 3298 6820
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 5442 6808 5448 6860
rect 5500 6808 5506 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 6972 6820 7205 6848
rect 6972 6808 6978 6820
rect 7193 6817 7205 6820
rect 7239 6817 7251 6851
rect 10428 6848 10456 6888
rect 7193 6811 7251 6817
rect 8036 6820 10456 6848
rect 10520 6820 10916 6848
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2774 6780 2780 6792
rect 2455 6752 2780 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3568 6752 3801 6780
rect 3568 6740 3574 6752
rect 3789 6749 3801 6752
rect 3835 6780 3847 6783
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3835 6752 4077 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4065 6743 4123 6749
rect 4172 6752 4353 6780
rect 4172 6656 4200 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 8036 6780 8064 6820
rect 7055 6752 8064 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8168 6752 8309 6780
rect 8168 6740 8174 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 8812 6752 9413 6780
rect 8812 6740 8818 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 5712 6715 5770 6721
rect 5712 6681 5724 6715
rect 5758 6712 5770 6715
rect 6362 6712 6368 6724
rect 5758 6684 6368 6712
rect 5758 6681 5770 6684
rect 5712 6675 5770 6681
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 6730 6672 6736 6724
rect 6788 6712 6794 6724
rect 9030 6712 9036 6724
rect 6788 6684 9036 6712
rect 6788 6672 6794 6684
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 9508 6712 9536 6743
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 10520 6789 10548 6820
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9640 6752 9781 6780
rect 9640 6740 9646 6752
rect 9769 6749 9781 6752
rect 9815 6780 9827 6783
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 9815 6752 10241 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10778 6740 10784 6792
rect 10836 6740 10842 6792
rect 10888 6780 10916 6820
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11112 6820 11805 6848
rect 11112 6808 11118 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11900 6848 11928 6888
rect 12342 6876 12348 6928
rect 12400 6916 12406 6928
rect 13446 6916 13452 6928
rect 12400 6888 13452 6916
rect 12400 6876 12406 6888
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 15948 6916 15976 6944
rect 14415 6888 15976 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 11974 6848 11980 6860
rect 11900 6820 11980 6848
rect 11793 6811 11851 6817
rect 11974 6808 11980 6820
rect 12032 6848 12038 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12032 6820 12541 6848
rect 12032 6808 12038 6820
rect 12529 6817 12541 6820
rect 12575 6848 12587 6851
rect 16040 6848 16068 6944
rect 16761 6919 16819 6925
rect 16761 6885 16773 6919
rect 16807 6916 16819 6919
rect 17954 6916 17960 6928
rect 16807 6888 17960 6916
rect 16807 6885 16819 6888
rect 16761 6879 16819 6885
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 20732 6916 20760 6956
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 22186 6944 22192 6996
rect 22244 6984 22250 6996
rect 22741 6987 22799 6993
rect 22741 6984 22753 6987
rect 22244 6956 22753 6984
rect 22244 6944 22250 6956
rect 22741 6953 22753 6956
rect 22787 6953 22799 6987
rect 22741 6947 22799 6953
rect 23842 6944 23848 6996
rect 23900 6984 23906 6996
rect 26234 6984 26240 6996
rect 23900 6956 26240 6984
rect 23900 6944 23906 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 26602 6944 26608 6996
rect 26660 6984 26666 6996
rect 26697 6987 26755 6993
rect 26697 6984 26709 6987
rect 26660 6956 26709 6984
rect 26660 6944 26666 6956
rect 26697 6953 26709 6956
rect 26743 6953 26755 6987
rect 26697 6947 26755 6953
rect 18104 6888 20760 6916
rect 20824 6888 22232 6916
rect 18104 6876 18110 6888
rect 16574 6848 16580 6860
rect 12575 6820 13768 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 10888 6752 11652 6780
rect 11624 6712 11652 6752
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13630 6780 13636 6792
rect 13403 6752 13636 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 11974 6712 11980 6724
rect 9140 6684 9352 6712
rect 9508 6684 10088 6712
rect 11624 6684 11980 6712
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2866 6644 2872 6656
rect 2547 6616 2872 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3510 6604 3516 6656
rect 3568 6604 3574 6656
rect 4154 6604 4160 6656
rect 4212 6604 4218 6656
rect 4982 6604 4988 6656
rect 5040 6604 5046 6656
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 9140 6644 9168 6684
rect 8159 6616 9168 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 9214 6604 9220 6656
rect 9272 6604 9278 6656
rect 9324 6644 9352 6684
rect 9490 6644 9496 6656
rect 9324 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 10060 6653 10088 6684
rect 11974 6672 11980 6684
rect 12032 6672 12038 6724
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12728 6712 12756 6743
rect 12124 6684 12756 6712
rect 12124 6672 12130 6684
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 13372 6644 13400 6743
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13740 6721 13768 6820
rect 14292 6820 15240 6848
rect 14292 6792 14320 6820
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 14056 6752 14105 6780
rect 14056 6740 14062 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 15212 6789 15240 6820
rect 15304 6820 16068 6848
rect 16500 6820 16580 6848
rect 15304 6789 15332 6820
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 13725 6715 13783 6721
rect 13725 6681 13737 6715
rect 13771 6712 13783 6715
rect 14476 6712 14504 6740
rect 13771 6684 14504 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 10643 6616 13400 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 14148 6616 14197 6644
rect 14148 6604 14154 6616
rect 14185 6613 14197 6616
rect 14231 6613 14243 6647
rect 14568 6644 14596 6743
rect 14660 6712 14688 6743
rect 15102 6712 15108 6724
rect 14660 6684 15108 6712
rect 15102 6672 15108 6684
rect 15160 6712 15166 6724
rect 15304 6712 15332 6743
rect 15160 6684 15332 6712
rect 15160 6672 15166 6684
rect 15764 6656 15792 6743
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16500 6789 16528 6820
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 17586 6848 17592 6860
rect 17236 6820 17592 6848
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15896 6752 15945 6780
rect 15896 6740 15902 6752
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 16224 6712 16252 6743
rect 15948 6684 16252 6712
rect 15948 6656 15976 6684
rect 16574 6672 16580 6724
rect 16632 6672 16638 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 16960 6712 16988 6743
rect 17034 6740 17040 6792
rect 17092 6789 17098 6792
rect 17092 6783 17119 6789
rect 17107 6780 17119 6783
rect 17236 6780 17264 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 18598 6808 18604 6860
rect 18656 6848 18662 6860
rect 20824 6848 20852 6888
rect 18656 6820 20852 6848
rect 18656 6808 18662 6820
rect 20898 6808 20904 6860
rect 20956 6808 20962 6860
rect 21450 6808 21456 6860
rect 21508 6848 21514 6860
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 21508 6820 21833 6848
rect 21508 6808 21514 6820
rect 21821 6817 21833 6820
rect 21867 6817 21879 6851
rect 22204 6848 22232 6888
rect 22278 6876 22284 6928
rect 22336 6876 22342 6928
rect 23382 6876 23388 6928
rect 23440 6916 23446 6928
rect 24489 6919 24547 6925
rect 24489 6916 24501 6919
rect 23440 6888 24501 6916
rect 23440 6876 23446 6888
rect 24489 6885 24501 6888
rect 24535 6885 24547 6919
rect 27522 6916 27528 6928
rect 24489 6879 24547 6885
rect 24964 6888 27528 6916
rect 22370 6848 22376 6860
rect 22204 6820 22376 6848
rect 21821 6811 21879 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6848 22615 6851
rect 22922 6848 22928 6860
rect 22603 6820 22928 6848
rect 22603 6817 22615 6820
rect 22557 6811 22615 6817
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 23566 6808 23572 6860
rect 23624 6808 23630 6860
rect 24762 6848 24768 6860
rect 24596 6820 24768 6848
rect 17107 6752 17264 6780
rect 17107 6749 17119 6752
rect 17092 6743 17119 6749
rect 17092 6740 17098 6743
rect 17310 6740 17316 6792
rect 17368 6740 17374 6792
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17773 6783 17831 6789
rect 17543 6752 17632 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17328 6712 17356 6740
rect 16816 6684 17356 6712
rect 16816 6672 16822 6684
rect 14642 6644 14648 6656
rect 14568 6616 14648 6644
rect 14185 6607 14243 6613
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15286 6644 15292 6656
rect 15059 6616 15292 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15378 6604 15384 6656
rect 15436 6604 15442 6656
rect 15746 6604 15752 6656
rect 15804 6604 15810 6656
rect 15930 6604 15936 6656
rect 15988 6604 15994 6656
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 16206 6644 16212 6656
rect 16071 6616 16212 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16298 6604 16304 6656
rect 16356 6604 16362 6656
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17402 6644 17408 6656
rect 17175 6616 17408 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17604 6653 17632 6752
rect 17773 6749 17785 6783
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 17788 6712 17816 6743
rect 17862 6740 17868 6792
rect 17920 6780 17926 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17920 6752 18061 6780
rect 17920 6740 17926 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6780 18383 6783
rect 18506 6780 18512 6792
rect 18371 6752 18512 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6780 18843 6783
rect 19061 6783 19119 6789
rect 19061 6780 19073 6783
rect 18831 6752 19073 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 19061 6749 19073 6752
rect 19107 6780 19119 6783
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19107 6752 19257 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19245 6749 19257 6752
rect 19291 6780 19303 6783
rect 19334 6780 19340 6792
rect 19291 6752 19340 6780
rect 19291 6749 19303 6752
rect 19245 6743 19303 6749
rect 18800 6712 18828 6743
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19978 6740 19984 6792
rect 20036 6740 20042 6792
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 21600 6752 21649 6780
rect 21600 6740 21606 6752
rect 21637 6749 21649 6752
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 17788 6684 18828 6712
rect 17788 6656 17816 6684
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 20073 6715 20131 6721
rect 20073 6712 20085 6715
rect 19208 6684 20085 6712
rect 19208 6672 19214 6684
rect 20073 6681 20085 6684
rect 20119 6681 20131 6715
rect 20073 6675 20131 6681
rect 20533 6715 20591 6721
rect 20533 6681 20545 6715
rect 20579 6681 20591 6715
rect 20533 6675 20591 6681
rect 20625 6715 20683 6721
rect 20625 6681 20637 6715
rect 20671 6712 20683 6715
rect 21358 6712 21364 6724
rect 20671 6684 21364 6712
rect 20671 6681 20683 6684
rect 20625 6675 20683 6681
rect 17589 6647 17647 6653
rect 17589 6613 17601 6647
rect 17635 6613 17647 6647
rect 17589 6607 17647 6613
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 18230 6604 18236 6656
rect 18288 6604 18294 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 18601 6647 18659 6653
rect 18601 6613 18613 6647
rect 18647 6644 18659 6647
rect 19058 6644 19064 6656
rect 18647 6616 19064 6644
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 19300 6616 19901 6644
rect 19300 6604 19306 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 20548 6644 20576 6675
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 23124 6712 23152 6743
rect 24210 6740 24216 6792
rect 24268 6740 24274 6792
rect 24421 6783 24479 6789
rect 24421 6749 24433 6783
rect 24467 6780 24479 6783
rect 24596 6780 24624 6820
rect 24762 6808 24768 6820
rect 24820 6808 24826 6860
rect 24467 6752 24624 6780
rect 24673 6783 24731 6789
rect 24467 6749 24479 6752
rect 24421 6743 24479 6749
rect 24673 6749 24685 6783
rect 24719 6780 24731 6783
rect 24854 6780 24860 6792
rect 24719 6752 24860 6780
rect 24719 6749 24731 6752
rect 24673 6743 24731 6749
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 23382 6712 23388 6724
rect 21928 6684 23388 6712
rect 21928 6644 21956 6684
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 23661 6715 23719 6721
rect 23661 6681 23673 6715
rect 23707 6712 23719 6715
rect 24964 6712 24992 6888
rect 27522 6876 27528 6888
rect 27580 6916 27586 6928
rect 28169 6919 28227 6925
rect 28169 6916 28181 6919
rect 27580 6888 28181 6916
rect 27580 6876 27586 6888
rect 28169 6885 28181 6888
rect 28215 6885 28227 6919
rect 28169 6879 28227 6885
rect 25130 6808 25136 6860
rect 25188 6848 25194 6860
rect 26145 6851 26203 6857
rect 26145 6848 26157 6851
rect 25188 6820 26157 6848
rect 25188 6808 25194 6820
rect 26145 6817 26157 6820
rect 26191 6817 26203 6851
rect 26145 6811 26203 6817
rect 26602 6808 26608 6860
rect 26660 6848 26666 6860
rect 27065 6851 27123 6857
rect 27065 6848 27077 6851
rect 26660 6820 27077 6848
rect 26660 6808 26666 6820
rect 27065 6817 27077 6820
rect 27111 6817 27123 6851
rect 27065 6811 27123 6817
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 25133 6715 25191 6721
rect 25133 6712 25145 6715
rect 23707 6684 24900 6712
rect 24964 6684 25145 6712
rect 23707 6681 23719 6684
rect 23661 6675 23719 6681
rect 20548 6616 21956 6644
rect 19889 6607 19947 6613
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 22060 6616 23213 6644
rect 22060 6604 22066 6616
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 24670 6604 24676 6656
rect 24728 6644 24734 6656
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 24728 6616 24777 6644
rect 24728 6604 24734 6616
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24872 6644 24900 6684
rect 25133 6681 25145 6684
rect 25179 6681 25191 6715
rect 25133 6675 25191 6681
rect 25222 6672 25228 6724
rect 25280 6672 25286 6724
rect 25406 6672 25412 6724
rect 25464 6712 25470 6724
rect 25777 6715 25835 6721
rect 25777 6712 25789 6715
rect 25464 6684 25789 6712
rect 25464 6672 25470 6684
rect 25777 6681 25789 6684
rect 25823 6681 25835 6715
rect 25884 6712 25912 6743
rect 27246 6740 27252 6792
rect 27304 6740 27310 6792
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6780 27859 6783
rect 27890 6780 27896 6792
rect 27847 6752 27896 6780
rect 27847 6749 27859 6752
rect 27801 6743 27859 6749
rect 27890 6740 27896 6752
rect 27948 6740 27954 6792
rect 27982 6740 27988 6792
rect 28040 6740 28046 6792
rect 25884 6684 26372 6712
rect 25777 6675 25835 6681
rect 26344 6656 26372 6684
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 24872 6616 25973 6644
rect 24765 6607 24823 6613
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 26326 6604 26332 6656
rect 26384 6604 26390 6656
rect 27709 6647 27767 6653
rect 27709 6613 27721 6647
rect 27755 6644 27767 6647
rect 27798 6644 27804 6656
rect 27755 6616 27804 6644
rect 27755 6613 27767 6616
rect 27709 6607 27767 6613
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6409 5687 6443
rect 5629 6403 5687 6409
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 5644 6372 5672 6403
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6420 6412 7021 6440
rect 6420 6400 6426 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 8754 6400 8760 6452
rect 8812 6400 8818 6452
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6409 11759 6443
rect 11701 6403 11759 6409
rect 1452 6344 5488 6372
rect 5644 6344 7420 6372
rect 1452 6332 1458 6344
rect 2792 6313 2820 6344
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 3044 6307 3102 6313
rect 2823 6276 2857 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3044 6273 3056 6307
rect 3090 6304 3102 6307
rect 3786 6304 3792 6316
rect 3090 6276 3792 6304
rect 3090 6273 3102 6276
rect 3044 6267 3102 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 4264 6313 4292 6344
rect 5460 6316 5488 6344
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4516 6307 4574 6313
rect 4516 6273 4528 6307
rect 4562 6304 4574 6307
rect 4982 6304 4988 6316
rect 4562 6276 4988 6304
rect 4562 6273 4574 6276
rect 4516 6267 4574 6273
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 6380 6313 6408 6344
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 1995 6208 2774 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2746 6112 2774 6208
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5736 6236 5764 6267
rect 5316 6208 5764 6236
rect 5316 6196 5322 6208
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 6196 6168 6224 6267
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7392 6313 7420 6344
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7156 6276 7297 6304
rect 7156 6264 7162 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 7852 6236 7880 6267
rect 8202 6236 8208 6248
rect 7852 6208 8208 6236
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8496 6236 8524 6267
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9232 6313 9260 6400
rect 11716 6372 11744 6403
rect 12066 6400 12072 6452
rect 12124 6400 12130 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12342 6440 12348 6452
rect 12299 6412 12348 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12584 6412 12725 6440
rect 12584 6400 12590 6412
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 12713 6403 12771 6409
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 13688 6412 13829 6440
rect 13688 6400 13694 6412
rect 13817 6409 13829 6412
rect 13863 6440 13875 6443
rect 14182 6440 14188 6452
rect 13863 6412 14188 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 15194 6400 15200 6452
rect 15252 6400 15258 6452
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 18598 6440 18604 6452
rect 15427 6412 18604 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 11716 6344 12940 6372
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11848 6276 11897 6304
rect 11848 6264 11854 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12066 6304 12072 6316
rect 12023 6276 12072 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 12912 6313 12940 6344
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14182 6304 14188 6316
rect 14047 6276 14188 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14599 6276 14933 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 14921 6273 14933 6276
rect 14967 6304 14979 6307
rect 15212 6304 15240 6400
rect 15304 6372 15332 6400
rect 15304 6344 15516 6372
rect 14967 6276 15240 6304
rect 15289 6307 15347 6313
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 8662 6236 8668 6248
rect 8496 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 9490 6236 9496 6248
rect 8720 6208 9496 6236
rect 8720 6196 8726 6208
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9640 6208 9781 6236
rect 9640 6196 9646 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 9950 6196 9956 6248
rect 10008 6196 10014 6248
rect 10502 6196 10508 6248
rect 10560 6196 10566 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 13078 6236 13084 6248
rect 10735 6208 13084 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13170 6196 13176 6248
rect 13228 6196 13234 6248
rect 13354 6196 13360 6248
rect 13412 6196 13418 6248
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 15304 6236 15332 6267
rect 14660 6208 15332 6236
rect 15488 6236 15516 6344
rect 15580 6313 15608 6412
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 19392 6412 20729 6440
rect 19392 6400 19398 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 21453 6443 21511 6449
rect 21453 6409 21465 6443
rect 21499 6440 21511 6443
rect 22278 6440 22284 6452
rect 21499 6412 22284 6440
rect 21499 6409 21511 6412
rect 21453 6403 21511 6409
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 22664 6412 24992 6440
rect 16758 6372 16764 6384
rect 16592 6344 16764 6372
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 15565 6267 15623 6273
rect 15672 6276 16497 6304
rect 15672 6236 15700 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 15488 6208 15700 6236
rect 15749 6239 15807 6245
rect 7101 6171 7159 6177
rect 7101 6168 7113 6171
rect 3936 6140 4292 6168
rect 3936 6128 3942 6140
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2372 6072 2513 6100
rect 2372 6060 2378 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2746 6072 2780 6112
rect 2501 6063 2559 6069
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 4154 6060 4160 6112
rect 4212 6060 4218 6112
rect 4264 6100 4292 6140
rect 5184 6140 5948 6168
rect 6196 6140 7113 6168
rect 5184 6100 5212 6140
rect 4264 6072 5212 6100
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 5920 6100 5948 6140
rect 7101 6137 7113 6140
rect 7147 6137 7159 6171
rect 10413 6171 10471 6177
rect 7101 6131 7159 6137
rect 7208 6140 9720 6168
rect 7208 6100 7236 6140
rect 5920 6072 7236 6100
rect 7466 6060 7472 6112
rect 7524 6060 7530 6112
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 9692 6100 9720 6140
rect 10413 6137 10425 6171
rect 10459 6168 10471 6171
rect 10778 6168 10784 6180
rect 10459 6140 10784 6168
rect 10459 6137 10471 6140
rect 10413 6131 10471 6137
rect 10778 6128 10784 6140
rect 10836 6168 10842 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10836 6140 10885 6168
rect 10836 6128 10842 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 11054 6128 11060 6180
rect 11112 6168 11118 6180
rect 12434 6168 12440 6180
rect 11112 6140 12440 6168
rect 11112 6128 11118 6140
rect 12434 6128 12440 6140
rect 12492 6168 12498 6180
rect 12802 6168 12808 6180
rect 12492 6140 12808 6168
rect 12492 6128 12498 6140
rect 12802 6128 12808 6140
rect 12860 6168 12866 6180
rect 13556 6168 13584 6196
rect 14660 6168 14688 6208
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 16592 6236 16620 6344
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 20254 6372 20260 6384
rect 16960 6344 20260 6372
rect 16960 6313 16988 6344
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 22664 6316 22692 6412
rect 24964 6384 24992 6412
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 26602 6440 26608 6452
rect 25280 6412 26608 6440
rect 25280 6400 25286 6412
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 26789 6443 26847 6449
rect 26789 6409 26801 6443
rect 26835 6409 26847 6443
rect 26789 6403 26847 6409
rect 22916 6375 22974 6381
rect 22916 6341 22928 6375
rect 22962 6372 22974 6375
rect 23014 6372 23020 6384
rect 22962 6344 23020 6372
rect 22962 6341 22974 6344
rect 22916 6335 22974 6341
rect 23014 6332 23020 6344
rect 23072 6332 23078 6384
rect 24394 6372 24400 6384
rect 23952 6344 24400 6372
rect 23952 6316 23980 6344
rect 24394 6332 24400 6344
rect 24452 6332 24458 6384
rect 24486 6332 24492 6384
rect 24544 6372 24550 6384
rect 24765 6375 24823 6381
rect 24765 6372 24777 6375
rect 24544 6344 24777 6372
rect 24544 6332 24550 6344
rect 24765 6341 24777 6344
rect 24811 6341 24823 6375
rect 24765 6335 24823 6341
rect 24946 6332 24952 6384
rect 25004 6372 25010 6384
rect 25774 6372 25780 6384
rect 25004 6344 25780 6372
rect 25004 6332 25010 6344
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 16945 6307 17003 6313
rect 16715 6276 16896 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 15749 6199 15807 6205
rect 15856 6208 16620 6236
rect 12860 6140 13584 6168
rect 13740 6140 14688 6168
rect 15013 6171 15071 6177
rect 12860 6128 12866 6140
rect 13740 6100 13768 6140
rect 15013 6137 15025 6171
rect 15059 6168 15071 6171
rect 15764 6168 15792 6199
rect 15059 6140 15792 6168
rect 15059 6137 15071 6140
rect 15013 6131 15071 6137
rect 9692 6072 13768 6100
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15856 6100 15884 6208
rect 16022 6128 16028 6180
rect 16080 6168 16086 6180
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 16080 6140 16313 6168
rect 16080 6128 16086 6140
rect 16301 6137 16313 6140
rect 16347 6137 16359 6171
rect 16301 6131 16359 6137
rect 14700 6072 15884 6100
rect 14700 6060 14706 6072
rect 16206 6060 16212 6112
rect 16264 6060 16270 6112
rect 16758 6060 16764 6112
rect 16816 6060 16822 6112
rect 16868 6100 16896 6276
rect 16945 6273 16957 6307
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17212 6307 17270 6313
rect 17212 6273 17224 6307
rect 17258 6304 17270 6307
rect 18785 6307 18843 6313
rect 17258 6276 18736 6304
rect 17258 6273 17270 6276
rect 17212 6267 17270 6273
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 18598 6196 18604 6248
rect 18656 6196 18662 6248
rect 18708 6236 18736 6276
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 19150 6304 19156 6316
rect 18831 6276 19156 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6304 19395 6307
rect 19426 6304 19432 6316
rect 19383 6276 19432 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19604 6307 19662 6313
rect 19604 6273 19616 6307
rect 19650 6304 19662 6307
rect 19650 6276 20944 6304
rect 19650 6273 19662 6276
rect 19604 6267 19662 6273
rect 19260 6236 19288 6264
rect 18708 6208 19288 6236
rect 20806 6196 20812 6248
rect 20864 6196 20870 6248
rect 20916 6236 20944 6276
rect 20990 6264 20996 6316
rect 21048 6264 21054 6316
rect 21913 6307 21971 6313
rect 21913 6273 21925 6307
rect 21959 6304 21971 6307
rect 21959 6276 22600 6304
rect 21959 6273 21971 6276
rect 21913 6267 21971 6273
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 20916 6208 22477 6236
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22572 6236 22600 6276
rect 22646 6264 22652 6316
rect 22704 6264 22710 6316
rect 23934 6304 23940 6316
rect 22756 6276 23940 6304
rect 22756 6236 22784 6276
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 24026 6264 24032 6316
rect 24084 6304 24090 6316
rect 25424 6313 25452 6344
rect 25774 6332 25780 6344
rect 25832 6332 25838 6384
rect 26050 6332 26056 6384
rect 26108 6332 26114 6384
rect 26234 6332 26240 6384
rect 26292 6372 26298 6384
rect 26804 6372 26832 6403
rect 27890 6400 27896 6452
rect 27948 6440 27954 6452
rect 28353 6443 28411 6449
rect 28353 6440 28365 6443
rect 27948 6412 28365 6440
rect 27948 6400 27954 6412
rect 28353 6409 28365 6412
rect 28399 6409 28411 6443
rect 28353 6403 28411 6409
rect 26292 6344 27016 6372
rect 26292 6332 26298 6344
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 24084 6276 24133 6304
rect 24084 6264 24090 6276
rect 24121 6273 24133 6276
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 25676 6307 25734 6313
rect 25676 6273 25688 6307
rect 25722 6304 25734 6307
rect 26068 6304 26096 6332
rect 26988 6313 27016 6344
rect 25722 6276 26096 6304
rect 26973 6307 27031 6313
rect 25722 6273 25734 6276
rect 25676 6267 25734 6273
rect 26973 6273 26985 6307
rect 27019 6273 27031 6307
rect 26973 6267 27031 6273
rect 22572 6208 22784 6236
rect 24673 6239 24731 6245
rect 22465 6199 22523 6205
rect 24673 6205 24685 6239
rect 24719 6236 24731 6239
rect 25130 6236 25136 6248
rect 24719 6208 25136 6236
rect 24719 6205 24731 6208
rect 24673 6199 24731 6205
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 27709 6239 27767 6245
rect 27709 6205 27721 6239
rect 27755 6236 27767 6239
rect 27798 6236 27804 6248
rect 27755 6208 27804 6236
rect 27755 6205 27767 6208
rect 27709 6199 27767 6205
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 27893 6239 27951 6245
rect 27893 6205 27905 6239
rect 27939 6205 27951 6239
rect 27893 6199 27951 6205
rect 18432 6168 18460 6196
rect 18432 6140 19380 6168
rect 17678 6100 17684 6112
rect 16868 6072 17684 6100
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18322 6100 18328 6112
rect 18012 6072 18328 6100
rect 18012 6060 18018 6072
rect 18322 6060 18328 6072
rect 18380 6100 18386 6112
rect 19150 6100 19156 6112
rect 18380 6072 19156 6100
rect 18380 6060 18386 6072
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 19352 6100 19380 6140
rect 20640 6140 22094 6168
rect 20640 6100 20668 6140
rect 19352 6072 20668 6100
rect 22066 6100 22094 6140
rect 23584 6140 24992 6168
rect 23584 6100 23612 6140
rect 22066 6072 23612 6100
rect 24026 6060 24032 6112
rect 24084 6060 24090 6112
rect 24210 6060 24216 6112
rect 24268 6060 24274 6112
rect 24964 6100 24992 6140
rect 25038 6128 25044 6180
rect 25096 6168 25102 6180
rect 25225 6171 25283 6177
rect 25225 6168 25237 6171
rect 25096 6140 25237 6168
rect 25096 6128 25102 6140
rect 25225 6137 25237 6140
rect 25271 6168 25283 6171
rect 25406 6168 25412 6180
rect 25271 6140 25412 6168
rect 25271 6137 25283 6140
rect 25225 6131 25283 6137
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 27908 6168 27936 6199
rect 26344 6140 27936 6168
rect 26344 6100 26372 6140
rect 24964 6072 26372 6100
rect 27614 6060 27620 6112
rect 27672 6060 27678 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 3844 5868 4445 5896
rect 3844 5856 3850 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 5810 5856 5816 5908
rect 5868 5856 5874 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 7616 5868 7665 5896
rect 7616 5856 7622 5868
rect 7653 5865 7665 5868
rect 7699 5896 7711 5899
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 7699 5868 8401 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8389 5865 8401 5868
rect 8435 5865 8447 5899
rect 8389 5859 8447 5865
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 9582 5856 9588 5908
rect 9640 5856 9646 5908
rect 9950 5856 9956 5908
rect 10008 5896 10014 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10008 5868 10885 5896
rect 10008 5856 10014 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 11149 5899 11207 5905
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 11698 5896 11704 5908
rect 11195 5868 11704 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 13078 5856 13084 5908
rect 13136 5856 13142 5908
rect 13170 5856 13176 5908
rect 13228 5856 13234 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13354 5896 13360 5908
rect 13311 5868 13360 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 15746 5856 15752 5908
rect 15804 5856 15810 5908
rect 16022 5856 16028 5908
rect 16080 5856 16086 5908
rect 16206 5856 16212 5908
rect 16264 5856 16270 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17862 5896 17868 5908
rect 17276 5868 17868 5896
rect 17276 5856 17282 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19300 5868 19625 5896
rect 19300 5856 19306 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 20898 5856 20904 5908
rect 20956 5856 20962 5908
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 21416 5868 22094 5896
rect 21416 5856 21422 5868
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1412 5732 2053 5760
rect 1412 5704 1440 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 3436 5760 3464 5856
rect 5828 5769 5856 5856
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3436 5732 3801 5760
rect 2041 5723 2099 5729
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5729 5871 5763
rect 7484 5760 7512 5856
rect 5813 5723 5871 5729
rect 6472 5732 7512 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1854 5692 1860 5704
rect 1627 5664 1860 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 2314 5701 2320 5704
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 2308 5692 2320 5701
rect 2275 5664 2320 5692
rect 1949 5655 2007 5661
rect 2308 5655 2320 5664
rect 1964 5624 1992 5655
rect 2314 5652 2320 5655
rect 2372 5652 2378 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4212 5664 4629 5692
rect 4212 5652 4218 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4755 5664 4905 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 6472 5692 6500 5732
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7800 5732 8217 5760
rect 7800 5720 7806 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8588 5760 8616 5856
rect 11072 5828 11100 5856
rect 9968 5800 11100 5828
rect 9125 5763 9183 5769
rect 9125 5760 9137 5763
rect 8588 5732 9137 5760
rect 8205 5723 8263 5729
rect 9125 5729 9137 5732
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 5675 5664 6500 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6730 5652 6736 5704
rect 6788 5652 6794 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 7208 5664 7297 5692
rect 1412 5596 1992 5624
rect 1412 5565 1440 5596
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5525 1455 5559
rect 1397 5519 1455 5525
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 3050 5556 3056 5568
rect 1811 5528 3056 5556
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 6270 5556 6276 5568
rect 5583 5528 6276 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7208 5565 7236 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7466 5652 7472 5704
rect 7524 5652 7530 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7616 5664 8033 5692
rect 7616 5652 7622 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9968 5701 9996 5800
rect 11238 5788 11244 5840
rect 11296 5788 11302 5840
rect 10042 5720 10048 5772
rect 10100 5720 10106 5772
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 11256 5760 11284 5788
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 10652 5732 11437 5760
rect 10652 5720 10658 5732
rect 11425 5729 11437 5732
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8352 5664 8953 5692
rect 8352 5652 8358 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10704 5664 11069 5692
rect 10704 5624 10732 5664
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11379 5664 11836 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11808 5636 11836 5664
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12820 5692 12848 5856
rect 13188 5760 13216 5856
rect 14093 5831 14151 5837
rect 14093 5797 14105 5831
rect 14139 5797 14151 5831
rect 15764 5828 15792 5856
rect 14093 5791 14151 5797
rect 14292 5800 15792 5828
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13188 5732 13553 5760
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12032 5664 12434 5692
rect 12820 5664 13001 5692
rect 12032 5652 12038 5664
rect 9784 5596 10732 5624
rect 9784 5565 9812 5596
rect 11514 5584 11520 5636
rect 11572 5624 11578 5636
rect 11670 5627 11728 5633
rect 11670 5624 11682 5627
rect 11572 5596 11682 5624
rect 11572 5584 11578 5596
rect 11670 5593 11682 5596
rect 11716 5593 11728 5627
rect 11670 5587 11728 5593
rect 11790 5584 11796 5636
rect 11848 5584 11854 5636
rect 12406 5624 12434 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 14108 5692 14136 5791
rect 14292 5701 14320 5800
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14424 5732 14841 5760
rect 14424 5720 14430 5732
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5760 15071 5763
rect 15286 5760 15292 5772
rect 15059 5732 15292 5760
rect 15059 5729 15071 5732
rect 15013 5723 15071 5729
rect 13495 5664 14136 5692
rect 14277 5695 14335 5701
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5661 14795 5695
rect 14844 5692 14872 5723
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 16040 5760 16068 5856
rect 15795 5732 16068 5760
rect 16224 5760 16252 5856
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 16669 5831 16727 5837
rect 16669 5828 16681 5831
rect 16632 5800 16681 5828
rect 16632 5788 16638 5800
rect 16669 5797 16681 5800
rect 16715 5797 16727 5831
rect 16669 5791 16727 5797
rect 17144 5800 18552 5828
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 16224 5732 16313 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 16301 5729 16313 5732
rect 16347 5729 16359 5763
rect 17144 5760 17172 5800
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 16301 5723 16359 5729
rect 16408 5732 17172 5760
rect 17236 5732 18429 5760
rect 15565 5695 15623 5701
rect 14844 5664 15516 5692
rect 14737 5655 14795 5661
rect 14366 5624 14372 5636
rect 12406 5596 14372 5624
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 14752 5624 14780 5655
rect 15194 5624 15200 5636
rect 14752 5596 15200 5624
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 15488 5624 15516 5664
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 16408 5692 16436 5732
rect 15611 5664 16436 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17236 5692 17264 5732
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18524 5760 18552 5800
rect 18598 5788 18604 5840
rect 18656 5788 18662 5840
rect 19981 5831 20039 5837
rect 19981 5828 19993 5831
rect 19444 5800 19993 5828
rect 19444 5769 19472 5800
rect 19981 5797 19993 5800
rect 20027 5797 20039 5831
rect 19981 5791 20039 5797
rect 19429 5763 19487 5769
rect 18524 5732 19288 5760
rect 18417 5723 18475 5729
rect 16816 5664 17264 5692
rect 17313 5695 17371 5701
rect 16816 5652 16822 5664
rect 17313 5661 17325 5695
rect 17359 5692 17371 5695
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17359 5664 17509 5692
rect 17359 5661 17371 5664
rect 17313 5655 17371 5661
rect 17497 5661 17509 5664
rect 17543 5692 17555 5695
rect 17770 5692 17776 5704
rect 17543 5664 17776 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 17880 5664 18245 5692
rect 17880 5624 17908 5664
rect 18233 5661 18245 5664
rect 18279 5692 18291 5695
rect 18322 5692 18328 5704
rect 18279 5664 18328 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 19260 5701 19288 5732
rect 19429 5729 19441 5763
rect 19475 5729 19487 5763
rect 19794 5760 19800 5772
rect 19429 5723 19487 5729
rect 19536 5732 19800 5760
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19536 5692 19564 5732
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 19886 5720 19892 5772
rect 19944 5760 19950 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 19944 5732 20269 5760
rect 19944 5720 19950 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20916 5760 20944 5856
rect 22066 5828 22094 5868
rect 23566 5856 23572 5908
rect 23624 5856 23630 5908
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 25130 5856 25136 5908
rect 25188 5896 25194 5908
rect 25498 5896 25504 5908
rect 25188 5868 25504 5896
rect 25188 5856 25194 5868
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 26237 5899 26295 5905
rect 26237 5865 26249 5899
rect 26283 5896 26295 5899
rect 26786 5896 26792 5908
rect 26283 5868 26792 5896
rect 26283 5865 26295 5868
rect 26237 5859 26295 5865
rect 26786 5856 26792 5868
rect 26844 5856 26850 5908
rect 27614 5856 27620 5908
rect 27672 5856 27678 5908
rect 27801 5899 27859 5905
rect 27801 5865 27813 5899
rect 27847 5896 27859 5899
rect 28534 5896 28540 5908
rect 27847 5868 28540 5896
rect 27847 5865 27859 5868
rect 27801 5859 27859 5865
rect 23753 5831 23811 5837
rect 23753 5828 23765 5831
rect 22066 5800 23765 5828
rect 23753 5797 23765 5800
rect 23799 5797 23811 5831
rect 23753 5791 23811 5797
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20916 5732 21005 5760
rect 20257 5723 20315 5729
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21177 5763 21235 5769
rect 21177 5729 21189 5763
rect 21223 5760 21235 5763
rect 21223 5732 22784 5760
rect 21223 5729 21235 5732
rect 21177 5723 21235 5729
rect 19291 5664 19564 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 19668 5664 20177 5692
rect 19668 5652 19674 5664
rect 20165 5661 20177 5664
rect 20211 5661 20223 5695
rect 20165 5655 20223 5661
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 15488 5596 17908 5624
rect 18049 5627 18107 5633
rect 18049 5593 18061 5627
rect 18095 5624 18107 5627
rect 19978 5624 19984 5636
rect 18095 5596 19984 5624
rect 18095 5593 18107 5596
rect 18049 5587 18107 5593
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 7156 5528 7205 5556
rect 7156 5516 7162 5528
rect 7193 5525 7205 5528
rect 7239 5525 7251 5559
rect 7193 5519 7251 5525
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5525 9827 5559
rect 9769 5519 9827 5525
rect 10594 5516 10600 5568
rect 10652 5556 10658 5568
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 10652 5528 10701 5556
rect 10652 5516 10658 5528
rect 10689 5525 10701 5528
rect 10735 5525 10747 5559
rect 10689 5519 10747 5525
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 15470 5516 15476 5568
rect 15528 5516 15534 5568
rect 17126 5516 17132 5568
rect 17184 5516 17190 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 18064 5556 18092 5587
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 17736 5528 18092 5556
rect 17736 5516 17742 5528
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 19150 5556 19156 5568
rect 18288 5528 19156 5556
rect 18288 5516 18294 5528
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19794 5556 19800 5568
rect 19392 5528 19800 5556
rect 19392 5516 19398 5528
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 22756 5556 22784 5732
rect 22830 5720 22836 5772
rect 22888 5760 22894 5772
rect 23017 5763 23075 5769
rect 23017 5760 23029 5763
rect 22888 5732 23029 5760
rect 22888 5720 22894 5732
rect 23017 5729 23029 5732
rect 23063 5729 23075 5763
rect 23017 5723 23075 5729
rect 23201 5763 23259 5769
rect 23201 5729 23213 5763
rect 23247 5760 23259 5763
rect 24228 5760 24256 5856
rect 24302 5788 24308 5840
rect 24360 5828 24366 5840
rect 25869 5831 25927 5837
rect 25869 5828 25881 5831
rect 24360 5800 25881 5828
rect 24360 5788 24366 5800
rect 25869 5797 25881 5800
rect 25915 5797 25927 5831
rect 25869 5791 25927 5797
rect 23247 5732 24256 5760
rect 23247 5729 23259 5732
rect 23201 5723 23259 5729
rect 25774 5720 25780 5772
rect 25832 5760 25838 5772
rect 26418 5760 26424 5772
rect 25832 5732 26424 5760
rect 25832 5720 25838 5732
rect 26418 5720 26424 5732
rect 26476 5720 26482 5772
rect 22922 5652 22928 5704
rect 22980 5652 22986 5704
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5661 23995 5695
rect 23937 5655 23995 5661
rect 22833 5627 22891 5633
rect 22833 5593 22845 5627
rect 22879 5624 22891 5627
rect 22940 5624 22968 5652
rect 22879 5596 22968 5624
rect 23952 5624 23980 5655
rect 24026 5652 24032 5704
rect 24084 5652 24090 5704
rect 24118 5652 24124 5704
rect 24176 5692 24182 5704
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 24176 5664 24409 5692
rect 24176 5652 24182 5664
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 24397 5655 24455 5661
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 24728 5664 24992 5692
rect 24728 5652 24734 5664
rect 24854 5624 24860 5636
rect 23952 5596 24860 5624
rect 22879 5593 22891 5596
rect 22833 5587 22891 5593
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 24964 5624 24992 5664
rect 25130 5652 25136 5704
rect 25188 5652 25194 5704
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25590 5692 25596 5704
rect 25363 5664 25596 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 25682 5652 25688 5704
rect 25740 5692 25746 5704
rect 26053 5695 26111 5701
rect 26053 5692 26065 5695
rect 25740 5664 26065 5692
rect 25740 5652 25746 5664
rect 26053 5661 26065 5664
rect 26099 5661 26111 5695
rect 26053 5655 26111 5661
rect 26142 5652 26148 5704
rect 26200 5652 26206 5704
rect 26688 5695 26746 5701
rect 26688 5661 26700 5695
rect 26734 5692 26746 5695
rect 27632 5692 27660 5856
rect 27908 5769 27936 5868
rect 28534 5856 28540 5868
rect 28592 5856 28598 5908
rect 27893 5763 27951 5769
rect 27893 5729 27905 5763
rect 27939 5729 27951 5763
rect 27893 5723 27951 5729
rect 26734 5664 27660 5692
rect 26734 5661 26746 5664
rect 26688 5655 26746 5661
rect 24964 5596 25176 5624
rect 24121 5559 24179 5565
rect 24121 5556 24133 5559
rect 22756 5528 24133 5556
rect 24121 5525 24133 5528
rect 24167 5525 24179 5559
rect 24121 5519 24179 5525
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 25148 5556 25176 5596
rect 27522 5584 27528 5636
rect 27580 5624 27586 5636
rect 28537 5627 28595 5633
rect 28537 5624 28549 5627
rect 27580 5596 28549 5624
rect 27580 5584 27586 5596
rect 28537 5593 28549 5596
rect 28583 5593 28595 5627
rect 28537 5587 28595 5593
rect 28166 5556 28172 5568
rect 25148 5528 28172 5556
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 5074 5352 5080 5364
rect 4755 5324 5080 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6730 5352 6736 5364
rect 6043 5324 6736 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 5736 5284 5764 5315
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 7098 5312 7104 5364
rect 7156 5312 7162 5364
rect 7466 5312 7472 5364
rect 7524 5312 7530 5364
rect 8938 5312 8944 5364
rect 8996 5312 9002 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5321 9183 5355
rect 9125 5315 9183 5321
rect 8294 5284 8300 5296
rect 5736 5256 6224 5284
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 1664 5219 1722 5225
rect 1664 5185 1676 5219
rect 1710 5216 1722 5219
rect 2130 5216 2136 5228
rect 1710 5188 2136 5216
rect 1710 5185 1722 5188
rect 1664 5179 1722 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3568 5188 3801 5216
rect 3568 5176 3574 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4939 5188 5028 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3200 5120 3985 5148
rect 3200 5108 3206 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 5000 5089 5028 5188
rect 5092 5188 5181 5216
rect 5092 5160 5120 5188
rect 5169 5185 5181 5188
rect 5215 5216 5227 5219
rect 5258 5216 5264 5228
rect 5215 5188 5264 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5902 5176 5908 5228
rect 5960 5225 5966 5228
rect 6196 5225 6224 5256
rect 7576 5256 8300 5284
rect 5960 5179 5971 5225
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5185 6239 5219
rect 6181 5179 6239 5185
rect 5960 5176 5966 5179
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6328 5188 6469 5216
rect 6328 5176 6334 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 7401 5219 7459 5225
rect 7401 5185 7413 5219
rect 7447 5216 7459 5219
rect 7576 5216 7604 5256
rect 8294 5244 8300 5256
rect 8352 5284 8358 5296
rect 8956 5284 8984 5312
rect 9140 5284 9168 5315
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9769 5355 9827 5361
rect 9548 5324 9720 5352
rect 9548 5312 9554 5324
rect 9692 5284 9720 5324
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10226 5352 10232 5364
rect 9815 5324 10232 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10594 5312 10600 5364
rect 10652 5312 10658 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11514 5352 11520 5364
rect 11379 5324 11520 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 15470 5312 15476 5364
rect 15528 5312 15534 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16482 5352 16488 5364
rect 16347 5324 16488 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16574 5312 16580 5364
rect 16632 5312 16638 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5321 16727 5355
rect 17310 5352 17316 5364
rect 16669 5315 16727 5321
rect 16776 5324 17316 5352
rect 12066 5284 12072 5296
rect 8352 5256 8524 5284
rect 8956 5256 9076 5284
rect 9140 5256 9628 5284
rect 8352 5244 8358 5256
rect 7447 5188 7604 5216
rect 7447 5185 7459 5188
rect 7401 5179 7459 5185
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8496 5225 8524 5256
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7708 5188 7849 5216
rect 7708 5176 7714 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8389 5219 8447 5225
rect 8159 5188 8248 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 5074 5108 5080 5160
rect 5132 5108 5138 5160
rect 6638 5108 6644 5160
rect 6696 5108 6702 5160
rect 7742 5108 7748 5160
rect 7800 5108 7806 5160
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5049 5043 5083
rect 6546 5080 6552 5092
rect 4985 5043 5043 5049
rect 5092 5052 6552 5080
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 3559 4984 4445 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 4433 4981 4445 4984
rect 4479 5012 4491 5015
rect 5092 5012 5120 5052
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 7653 5083 7711 5089
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 7760 5080 7788 5108
rect 8220 5089 8248 5188
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8527 5188 8953 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9048 5216 9076 5256
rect 9600 5225 9628 5256
rect 9692 5256 12072 5284
rect 9692 5225 9720 5256
rect 12066 5244 12072 5256
rect 12124 5244 12130 5296
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 13817 5287 13875 5293
rect 13136 5256 13676 5284
rect 13136 5244 13142 5256
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9048 5188 9321 5216
rect 8941 5179 8999 5185
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5185 9735 5219
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 9677 5179 9735 5185
rect 9876 5188 10793 5216
rect 8404 5148 8432 5179
rect 8404 5120 8708 5148
rect 7699 5052 7788 5080
rect 8205 5083 8263 5089
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8205 5049 8217 5083
rect 8251 5049 8263 5083
rect 8205 5043 8263 5049
rect 8680 5024 8708 5120
rect 4479 4984 5120 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5258 4972 5264 5024
rect 5316 4972 5322 5024
rect 7929 5015 7987 5021
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8294 5012 8300 5024
rect 7975 4984 8300 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 8444 4984 8585 5012
rect 8444 4972 8450 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 8573 4975 8631 4981
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 8754 4972 8760 5024
rect 8812 4972 8818 5024
rect 8956 5012 8984 5179
rect 9324 5148 9352 5179
rect 9876 5148 9904 5188
rect 10781 5185 10793 5188
rect 10827 5216 10839 5219
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 10827 5188 11713 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11701 5185 11713 5188
rect 11747 5216 11759 5219
rect 11790 5216 11796 5228
rect 11747 5188 11796 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 13648 5225 13676 5256
rect 13817 5253 13829 5287
rect 13863 5284 13875 5287
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13863 5256 14197 5284
rect 13863 5253 13875 5256
rect 13817 5247 13875 5253
rect 14185 5253 14197 5256
rect 14231 5253 14243 5287
rect 14185 5247 14243 5253
rect 14550 5244 14556 5296
rect 14608 5284 14614 5296
rect 14608 5256 15056 5284
rect 14608 5244 14614 5256
rect 15028 5225 15056 5256
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13633 5219 13691 5225
rect 13219 5188 13492 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 9324 5120 9904 5148
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5148 10011 5151
rect 10042 5148 10048 5160
rect 9999 5120 10048 5148
rect 9999 5117 10011 5120
rect 9953 5111 10011 5117
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 9401 5083 9459 5089
rect 9401 5049 9413 5083
rect 9447 5080 9459 5083
rect 10152 5080 10180 5111
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 12621 5151 12679 5157
rect 12621 5148 12633 5151
rect 12584 5120 12633 5148
rect 12584 5108 12590 5120
rect 12621 5117 12633 5120
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 9447 5052 10180 5080
rect 9447 5049 9459 5052
rect 9401 5043 9459 5049
rect 10686 5040 10692 5092
rect 10744 5040 10750 5092
rect 13464 5089 13492 5188
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15488 5216 15516 5312
rect 16209 5287 16267 5293
rect 16209 5253 16221 5287
rect 16255 5284 16267 5287
rect 16592 5284 16620 5312
rect 16255 5256 16620 5284
rect 16255 5253 16267 5256
rect 16209 5247 16267 5253
rect 15565 5219 15623 5225
rect 15565 5216 15577 5219
rect 15488 5188 15577 5216
rect 15013 5179 15071 5185
rect 15565 5185 15577 5188
rect 15611 5185 15623 5219
rect 16485 5219 16543 5225
rect 15565 5179 15623 5185
rect 15672 5188 15884 5216
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 13740 5148 13768 5179
rect 13596 5120 13768 5148
rect 14093 5151 14151 5157
rect 13596 5108 13602 5120
rect 14093 5117 14105 5151
rect 14139 5117 14151 5151
rect 14093 5111 14151 5117
rect 13449 5083 13507 5089
rect 13449 5049 13461 5083
rect 13495 5049 13507 5083
rect 13449 5043 13507 5049
rect 10704 5012 10732 5040
rect 8956 4984 10732 5012
rect 12802 4972 12808 5024
rect 12860 4972 12866 5024
rect 13354 4972 13360 5024
rect 13412 4972 13418 5024
rect 14108 5012 14136 5111
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 14366 5108 14372 5160
rect 14424 5108 14430 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15672 5148 15700 5188
rect 14875 5120 15700 5148
rect 15749 5151 15807 5157
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 15856 5148 15884 5188
rect 16485 5185 16497 5219
rect 16531 5216 16543 5219
rect 16684 5216 16712 5315
rect 16531 5188 16712 5216
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 16776 5148 16804 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18288 5324 18429 5352
rect 18288 5312 18294 5324
rect 18417 5321 18429 5324
rect 18463 5352 18475 5355
rect 18598 5352 18604 5364
rect 18463 5324 18604 5352
rect 18463 5321 18475 5324
rect 18417 5315 18475 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 20622 5352 20628 5364
rect 18708 5324 20628 5352
rect 18708 5284 18736 5324
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 21913 5355 21971 5361
rect 21913 5352 21925 5355
rect 20864 5324 21925 5352
rect 20864 5312 20870 5324
rect 21913 5321 21925 5324
rect 21959 5321 21971 5355
rect 21913 5315 21971 5321
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 23842 5352 23848 5364
rect 23256 5324 23848 5352
rect 23256 5312 23262 5324
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 24121 5355 24179 5361
rect 24121 5352 24133 5355
rect 23992 5324 24133 5352
rect 23992 5312 23998 5324
rect 24121 5321 24133 5324
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 24857 5355 24915 5361
rect 24857 5321 24869 5355
rect 24903 5352 24915 5355
rect 25130 5352 25136 5364
rect 24903 5324 25136 5352
rect 24903 5321 24915 5324
rect 24857 5315 24915 5321
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 25498 5312 25504 5364
rect 25556 5352 25562 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 25556 5324 25789 5352
rect 25556 5312 25562 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 26694 5352 26700 5364
rect 25777 5315 25835 5321
rect 25884 5324 26700 5352
rect 17052 5256 18552 5284
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 15856 5120 16804 5148
rect 16868 5148 16896 5179
rect 16942 5148 16948 5160
rect 16868 5120 16948 5148
rect 15749 5111 15807 5117
rect 14292 5080 14320 5108
rect 14844 5080 14872 5111
rect 14292 5052 14872 5080
rect 15764 5080 15792 5111
rect 16942 5108 16948 5120
rect 17000 5148 17006 5160
rect 17052 5148 17080 5256
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 18524 5225 18552 5256
rect 18616 5256 18736 5284
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17368 5188 17785 5216
rect 17368 5176 17374 5188
rect 17773 5185 17785 5188
rect 17819 5216 17831 5219
rect 18509 5219 18567 5225
rect 17819 5188 18276 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 17000 5120 17080 5148
rect 17129 5151 17187 5157
rect 17000 5108 17006 5120
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17586 5148 17592 5160
rect 17175 5120 17592 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17586 5108 17592 5120
rect 17644 5148 17650 5160
rect 17862 5148 17868 5160
rect 17644 5120 17868 5148
rect 17644 5108 17650 5120
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 17954 5108 17960 5160
rect 18012 5108 18018 5160
rect 18248 5148 18276 5188
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18616 5148 18644 5256
rect 18782 5244 18788 5296
rect 18840 5284 18846 5296
rect 19334 5284 19340 5296
rect 18840 5256 19340 5284
rect 18840 5244 18846 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 19797 5287 19855 5293
rect 19797 5284 19809 5287
rect 19576 5256 19809 5284
rect 19576 5244 19582 5256
rect 19797 5253 19809 5256
rect 19843 5253 19855 5287
rect 19797 5247 19855 5253
rect 19886 5244 19892 5296
rect 19944 5244 19950 5296
rect 20438 5244 20444 5296
rect 20496 5284 20502 5296
rect 22465 5287 22523 5293
rect 22465 5284 22477 5287
rect 20496 5256 22477 5284
rect 20496 5244 20502 5256
rect 22465 5253 22477 5256
rect 22511 5253 22523 5287
rect 22465 5247 22523 5253
rect 23008 5287 23066 5293
rect 23008 5253 23020 5287
rect 23054 5284 23066 5287
rect 25038 5284 25044 5296
rect 23054 5256 25044 5284
rect 23054 5253 23066 5256
rect 23008 5247 23066 5253
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5216 19027 5219
rect 19242 5216 19248 5228
rect 19015 5188 19248 5216
rect 19015 5185 19027 5188
rect 18969 5179 19027 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 20772 5188 21220 5216
rect 20772 5176 20778 5188
rect 18248 5120 18644 5148
rect 19153 5151 19211 5157
rect 19153 5117 19165 5151
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5148 20683 5151
rect 21082 5148 21088 5160
rect 20671 5120 21088 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 18601 5083 18659 5089
rect 18601 5080 18613 5083
rect 15764 5052 16804 5080
rect 15378 5012 15384 5024
rect 14108 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16776 5012 16804 5052
rect 16951 5052 18613 5080
rect 16951 5012 16979 5052
rect 18601 5049 18613 5052
rect 18647 5049 18659 5083
rect 19168 5080 19196 5111
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 21192 5148 21220 5188
rect 21266 5176 21272 5228
rect 21324 5176 21330 5228
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5216 21419 5219
rect 21634 5216 21640 5228
rect 21407 5188 21640 5216
rect 21407 5185 21419 5188
rect 21361 5179 21419 5185
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21744 5188 21833 5216
rect 21744 5148 21772 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 22097 5219 22155 5225
rect 22097 5216 22109 5219
rect 21968 5188 22109 5216
rect 21968 5176 21974 5188
rect 22097 5185 22109 5188
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 22381 5219 22439 5225
rect 22381 5185 22393 5219
rect 22427 5216 22439 5219
rect 22427 5188 22508 5216
rect 22427 5185 22439 5188
rect 22381 5179 22439 5185
rect 21192 5120 21772 5148
rect 22480 5148 22508 5188
rect 22646 5176 22652 5228
rect 22704 5216 22710 5228
rect 22741 5219 22799 5225
rect 22741 5216 22753 5219
rect 22704 5188 22753 5216
rect 22704 5176 22710 5188
rect 22741 5185 22753 5188
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 22848 5188 24348 5216
rect 22848 5148 22876 5188
rect 22480 5120 22876 5148
rect 24213 5151 24271 5157
rect 19168 5052 20300 5080
rect 18601 5043 18659 5049
rect 16776 4984 16979 5012
rect 17678 4972 17684 5024
rect 17736 4972 17742 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 19337 5015 19395 5021
rect 19337 5012 19349 5015
rect 18104 4984 19349 5012
rect 18104 4972 18110 4984
rect 19337 4981 19349 4984
rect 19383 4981 19395 5015
rect 20272 5012 20300 5052
rect 20346 5040 20352 5092
rect 20404 5040 20410 5092
rect 22094 5080 22100 5092
rect 20640 5052 21680 5080
rect 20640 5012 20668 5052
rect 20272 4984 20668 5012
rect 19337 4975 19395 4981
rect 21174 4972 21180 5024
rect 21232 4972 21238 5024
rect 21652 5012 21680 5052
rect 22020 5052 22100 5080
rect 22020 5012 22048 5052
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 22186 5040 22192 5092
rect 22244 5040 22250 5092
rect 22370 5040 22376 5092
rect 22428 5080 22434 5092
rect 22480 5080 22508 5120
rect 24213 5117 24225 5151
rect 24259 5117 24271 5151
rect 24213 5111 24271 5117
rect 24228 5080 24256 5111
rect 22428 5052 22508 5080
rect 23676 5052 24256 5080
rect 22428 5040 22434 5052
rect 23676 5024 23704 5052
rect 21652 4984 22048 5012
rect 23658 4972 23664 5024
rect 23716 4972 23722 5024
rect 23750 4972 23756 5024
rect 23808 5012 23814 5024
rect 24210 5012 24216 5024
rect 23808 4984 24216 5012
rect 23808 4972 23814 4984
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 24320 5012 24348 5188
rect 24394 5176 24400 5228
rect 24452 5176 24458 5228
rect 24762 5176 24768 5228
rect 24820 5216 24826 5228
rect 25884 5216 25912 5324
rect 26694 5312 26700 5324
rect 26752 5312 26758 5364
rect 28534 5312 28540 5364
rect 28592 5312 28598 5364
rect 26878 5284 26884 5296
rect 25976 5256 26884 5284
rect 25976 5225 26004 5256
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 27424 5287 27482 5293
rect 27424 5253 27436 5287
rect 27470 5284 27482 5287
rect 27522 5284 27528 5296
rect 27470 5256 27528 5284
rect 27470 5253 27482 5256
rect 27424 5247 27482 5253
rect 27522 5244 27528 5256
rect 27580 5244 27586 5296
rect 24820 5188 25912 5216
rect 25961 5219 26019 5225
rect 24820 5176 24826 5188
rect 25961 5185 25973 5219
rect 26007 5185 26019 5219
rect 25961 5179 26019 5185
rect 26234 5176 26240 5228
rect 26292 5216 26298 5228
rect 26329 5219 26387 5225
rect 26329 5216 26341 5219
rect 26292 5188 26341 5216
rect 26292 5176 26298 5188
rect 26329 5185 26341 5188
rect 26375 5185 26387 5219
rect 26329 5179 26387 5185
rect 26418 5176 26424 5228
rect 26476 5216 26482 5228
rect 27154 5216 27160 5228
rect 26476 5188 27160 5216
rect 26476 5176 26482 5188
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 25133 5151 25191 5157
rect 25133 5117 25145 5151
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 25148 5080 25176 5111
rect 25314 5108 25320 5160
rect 25372 5108 25378 5160
rect 25774 5080 25780 5092
rect 25148 5052 25780 5080
rect 25774 5040 25780 5052
rect 25832 5040 25838 5092
rect 24946 5012 24952 5024
rect 24320 4984 24952 5012
rect 24946 4972 24952 4984
rect 25004 4972 25010 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 2130 4768 2136 4820
rect 2188 4768 2194 4820
rect 3878 4768 3884 4820
rect 3936 4768 3942 4820
rect 5258 4768 5264 4820
rect 5316 4768 5322 4820
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6696 4780 7205 4808
rect 6696 4768 6702 4780
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 7193 4771 7251 4777
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 8386 4768 8392 4820
rect 8444 4768 8450 4820
rect 8478 4768 8484 4820
rect 8536 4768 8542 4820
rect 12802 4808 12808 4820
rect 11072 4780 12808 4808
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 2130 4672 2136 4684
rect 1452 4644 2136 4672
rect 1452 4632 1458 4644
rect 2130 4632 2136 4644
rect 2188 4672 2194 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2188 4644 2237 4672
rect 2188 4632 2194 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 5276 4672 5304 4768
rect 5902 4740 5908 4752
rect 4387 4644 5304 4672
rect 5644 4712 5908 4740
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 1946 4604 1952 4616
rect 1627 4576 1952 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 2372 4576 3801 4604
rect 2372 4564 2378 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4706 4604 4712 4616
rect 4203 4576 4712 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5074 4604 5080 4616
rect 4939 4576 5080 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5644 4613 5672 4712
rect 5902 4700 5908 4712
rect 5960 4740 5966 4752
rect 6825 4743 6883 4749
rect 5960 4712 6500 4740
rect 5960 4700 5966 4712
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5767 4644 6377 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6472 4672 6500 4712
rect 6825 4709 6837 4743
rect 6871 4740 6883 4743
rect 6914 4740 6920 4752
rect 6871 4712 6920 4740
rect 6871 4709 6883 4712
rect 6825 4703 6883 4709
rect 6914 4700 6920 4712
rect 6972 4740 6978 4752
rect 7576 4740 7604 4768
rect 6972 4712 7604 4740
rect 6972 4700 6978 4712
rect 6472 4644 6960 4672
rect 6365 4635 6423 4641
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5583 4576 5641 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5629 4573 5641 4576
rect 5675 4604 5687 4607
rect 5905 4607 5963 4613
rect 5905 4604 5917 4607
rect 5675 4576 5917 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 5905 4573 5917 4576
rect 5951 4573 5963 4607
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5905 4567 5963 4573
rect 6012 4576 6193 4604
rect 1964 4468 1992 4564
rect 2492 4539 2550 4545
rect 2492 4505 2504 4539
rect 2538 4536 2550 4539
rect 4246 4536 4252 4548
rect 2538 4508 4252 4536
rect 2538 4505 2550 4508
rect 2492 4499 2550 4505
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 6012 4536 6040 4576
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6932 4600 6960 4644
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 7064 4644 7389 4672
rect 7064 4632 7070 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 8297 4675 8355 4681
rect 7377 4635 7435 4641
rect 7475 4644 7696 4672
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 7015 4600 7113 4604
rect 6932 4576 7113 4600
rect 6932 4572 7043 4576
rect 7101 4573 7113 4576
rect 7147 4604 7159 4607
rect 7475 4604 7503 4644
rect 7147 4576 7503 4604
rect 7561 4607 7619 4613
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7561 4573 7573 4607
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 4816 4508 6040 4536
rect 4816 4480 4844 4508
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 1964 4440 3617 4468
rect 3605 4437 3617 4440
rect 3651 4437 3663 4471
rect 3605 4431 3663 4437
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 4982 4428 4988 4480
rect 5040 4428 5046 4480
rect 5353 4471 5411 4477
rect 5353 4437 5365 4471
rect 5399 4468 5411 4471
rect 5810 4468 5816 4480
rect 5399 4440 5816 4468
rect 5399 4437 5411 4440
rect 5353 4431 5411 4437
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 7576 4468 7604 4567
rect 7668 4536 7696 4644
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8404 4672 8432 4768
rect 8496 4740 8524 4768
rect 11072 4749 11100 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13446 4808 13452 4820
rect 13035 4780 13452 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 14366 4768 14372 4820
rect 14424 4768 14430 4820
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 16022 4808 16028 4820
rect 15804 4780 16028 4808
rect 15804 4768 15810 4780
rect 16022 4768 16028 4780
rect 16080 4808 16086 4820
rect 16942 4808 16948 4820
rect 16080 4780 16948 4808
rect 16080 4768 16086 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 18012 4780 19257 4808
rect 18012 4768 18018 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 20714 4808 20720 4820
rect 19392 4780 20720 4808
rect 19392 4768 19398 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22189 4811 22247 4817
rect 22189 4808 22201 4811
rect 22152 4780 22201 4808
rect 22152 4768 22158 4780
rect 22189 4777 22201 4780
rect 22235 4777 22247 4811
rect 22189 4771 22247 4777
rect 22370 4768 22376 4820
rect 22428 4768 22434 4820
rect 24302 4808 24308 4820
rect 22480 4780 24308 4808
rect 9401 4743 9459 4749
rect 9401 4740 9413 4743
rect 8496 4712 9413 4740
rect 9401 4709 9413 4712
rect 9447 4709 9459 4743
rect 9401 4703 9459 4709
rect 9769 4743 9827 4749
rect 9769 4709 9781 4743
rect 9815 4709 9827 4743
rect 11057 4743 11115 4749
rect 11057 4740 11069 4743
rect 9769 4703 9827 4709
rect 9876 4712 11069 4740
rect 8343 4644 8432 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 8754 4632 8760 4684
rect 8812 4632 8818 4684
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9784 4672 9812 4703
rect 9263 4644 9812 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 8067 4576 8125 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8113 4573 8125 4576
rect 8159 4604 8171 4607
rect 8570 4604 8576 4616
rect 8159 4576 8576 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 8772 4536 8800 4632
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9876 4604 9904 4712
rect 11057 4709 11069 4712
rect 11103 4709 11115 4743
rect 13078 4740 13084 4752
rect 11057 4703 11115 4709
rect 12912 4712 13084 4740
rect 10226 4672 10232 4684
rect 10060 4644 10232 4672
rect 10060 4613 10088 4644
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10459 4644 10793 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 11296 4644 11345 4672
rect 11296 4632 11302 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 9079 4576 9904 4604
rect 9953 4607 10011 4613
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9953 4573 9965 4607
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 9968 4536 9996 4567
rect 10336 4536 10364 4567
rect 10594 4564 10600 4616
rect 10652 4564 10658 4616
rect 12912 4613 12940 4712
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13648 4672 13676 4768
rect 13722 4700 13728 4752
rect 13780 4740 13786 4752
rect 13817 4743 13875 4749
rect 13817 4740 13829 4743
rect 13780 4712 13829 4740
rect 13780 4700 13786 4712
rect 13817 4709 13829 4712
rect 13863 4740 13875 4743
rect 14384 4740 14412 4768
rect 13863 4712 14412 4740
rect 17144 4740 17172 4768
rect 17144 4712 19472 4740
rect 13863 4709 13875 4712
rect 13817 4703 13875 4709
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 13311 4644 13676 4672
rect 13924 4644 14289 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 11330 4536 11336 4548
rect 7668 4508 8708 4536
rect 8772 4508 9996 4536
rect 10060 4508 11336 4536
rect 8680 4480 8708 4508
rect 6043 4440 7604 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 10060 4468 10088 4508
rect 11330 4496 11336 4508
rect 11388 4496 11394 4548
rect 11600 4539 11658 4545
rect 11600 4505 11612 4539
rect 11646 4536 11658 4539
rect 12802 4536 12808 4548
rect 11646 4508 12808 4536
rect 11646 4505 11658 4508
rect 11600 4499 11658 4505
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 13350 4539 13408 4545
rect 13350 4505 13362 4539
rect 13396 4505 13408 4539
rect 13350 4499 13408 4505
rect 8720 4440 10088 4468
rect 8720 4428 8726 4440
rect 10134 4428 10140 4480
rect 10192 4428 10198 4480
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 11848 4440 12725 4468
rect 11848 4428 11854 4440
rect 12713 4437 12725 4440
rect 12759 4437 12771 4471
rect 13372 4468 13400 4499
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 13924 4536 13952 4644
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 14277 4635 14335 4641
rect 15286 4632 15292 4684
rect 15344 4632 15350 4684
rect 16114 4632 16120 4684
rect 16172 4632 16178 4684
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16264 4644 17049 4672
rect 16264 4632 16270 4644
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 18138 4672 18144 4684
rect 17635 4644 18144 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18248 4644 19196 4672
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 13504 4508 13952 4536
rect 14108 4536 14136 4567
rect 16316 4536 16344 4567
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16632 4576 16865 4604
rect 16632 4564 16638 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17770 4564 17776 4616
rect 17828 4564 17834 4616
rect 18248 4604 18276 4644
rect 17880 4576 18276 4604
rect 17880 4536 17908 4576
rect 14108 4508 15884 4536
rect 16316 4508 17908 4536
rect 13504 4496 13510 4508
rect 14090 4468 14096 4480
rect 13372 4440 14096 4468
rect 12713 4431 12771 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 15856 4468 15884 4508
rect 18046 4496 18052 4548
rect 18104 4496 18110 4548
rect 18138 4496 18144 4548
rect 18196 4536 18202 4548
rect 18196 4508 18368 4536
rect 18196 4496 18202 4508
rect 16761 4471 16819 4477
rect 16761 4468 16773 4471
rect 15856 4440 16773 4468
rect 16761 4437 16773 4440
rect 16807 4468 16819 4471
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 16807 4440 17509 4468
rect 16807 4437 16819 4440
rect 16761 4431 16819 4437
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 18064 4468 18092 4496
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 18064 4440 18245 4468
rect 17497 4431 17555 4437
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18340 4468 18368 4508
rect 18414 4496 18420 4548
rect 18472 4496 18478 4548
rect 18509 4539 18567 4545
rect 18509 4505 18521 4539
rect 18555 4505 18567 4539
rect 18509 4499 18567 4505
rect 18524 4468 18552 4499
rect 18782 4496 18788 4548
rect 18840 4536 18846 4548
rect 19061 4539 19119 4545
rect 19061 4536 19073 4539
rect 18840 4508 19073 4536
rect 18840 4496 18846 4508
rect 19061 4505 19073 4508
rect 19107 4505 19119 4539
rect 19168 4536 19196 4644
rect 19444 4613 19472 4712
rect 21082 4700 21088 4752
rect 21140 4740 21146 4752
rect 21177 4743 21235 4749
rect 21177 4740 21189 4743
rect 21140 4712 21189 4740
rect 21140 4700 21146 4712
rect 21177 4709 21189 4712
rect 21223 4740 21235 4743
rect 22388 4740 22416 4768
rect 21223 4712 22416 4740
rect 21223 4709 21235 4712
rect 21177 4703 21235 4709
rect 20824 4644 22416 4672
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19702 4564 19708 4616
rect 19760 4564 19766 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 19843 4576 20300 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 20272 4548 20300 4576
rect 20622 4564 20628 4616
rect 20680 4604 20686 4616
rect 20824 4604 20852 4644
rect 22388 4613 22416 4644
rect 20680 4576 20852 4604
rect 21545 4607 21603 4613
rect 20680 4564 20686 4576
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 22373 4607 22431 4613
rect 21591 4576 22094 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 20064 4539 20122 4545
rect 19168 4508 19564 4536
rect 19061 4499 19119 4505
rect 19536 4477 19564 4508
rect 20064 4505 20076 4539
rect 20110 4505 20122 4539
rect 20064 4499 20122 4505
rect 18340 4440 18552 4468
rect 19521 4471 19579 4477
rect 18233 4431 18291 4437
rect 19521 4437 19533 4471
rect 19567 4437 19579 4471
rect 20079 4468 20107 4499
rect 20254 4496 20260 4548
rect 20312 4496 20318 4548
rect 22066 4536 22094 4576
rect 22373 4573 22385 4607
rect 22419 4573 22431 4607
rect 22480 4604 22508 4780
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 25041 4811 25099 4817
rect 25041 4777 25053 4811
rect 25087 4808 25099 4811
rect 25130 4808 25136 4820
rect 25087 4780 25136 4808
rect 25087 4777 25099 4780
rect 25041 4771 25099 4777
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 25774 4768 25780 4820
rect 25832 4808 25838 4820
rect 26513 4811 26571 4817
rect 26513 4808 26525 4811
rect 25832 4780 26525 4808
rect 25832 4768 25838 4780
rect 26513 4777 26525 4780
rect 26559 4777 26571 4811
rect 26513 4771 26571 4777
rect 27798 4768 27804 4820
rect 27856 4808 27862 4820
rect 28261 4811 28319 4817
rect 28261 4808 28273 4811
rect 27856 4780 28273 4808
rect 27856 4768 27862 4780
rect 28261 4777 28273 4780
rect 28307 4777 28319 4811
rect 28261 4771 28319 4777
rect 23201 4743 23259 4749
rect 23201 4709 23213 4743
rect 23247 4740 23259 4743
rect 23658 4740 23664 4752
rect 23247 4712 23664 4740
rect 23247 4709 23259 4712
rect 23201 4703 23259 4709
rect 23658 4700 23664 4712
rect 23716 4700 23722 4752
rect 23842 4700 23848 4752
rect 23900 4740 23906 4752
rect 24029 4743 24087 4749
rect 24029 4740 24041 4743
rect 23900 4712 24041 4740
rect 23900 4700 23906 4712
rect 24029 4709 24041 4712
rect 24075 4709 24087 4743
rect 24029 4703 24087 4709
rect 24578 4700 24584 4752
rect 24636 4740 24642 4752
rect 24636 4712 28120 4740
rect 24636 4700 24642 4712
rect 22557 4675 22615 4681
rect 22557 4641 22569 4675
rect 22603 4672 22615 4675
rect 23750 4672 23756 4684
rect 22603 4644 23756 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 26973 4675 27031 4681
rect 26973 4672 26985 4675
rect 24136 4644 26985 4672
rect 22741 4607 22799 4613
rect 22741 4604 22753 4607
rect 22480 4576 22753 4604
rect 22373 4567 22431 4573
rect 22741 4573 22753 4576
rect 22787 4573 22799 4607
rect 22741 4567 22799 4573
rect 23198 4564 23204 4616
rect 23256 4564 23262 4616
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 23477 4607 23535 4613
rect 23477 4573 23489 4607
rect 23523 4604 23535 4607
rect 24136 4604 24164 4644
rect 26973 4641 26985 4644
rect 27019 4641 27031 4675
rect 26973 4635 27031 4641
rect 27062 4632 27068 4684
rect 27120 4672 27126 4684
rect 27157 4675 27215 4681
rect 27157 4672 27169 4675
rect 27120 4644 27169 4672
rect 27120 4632 27126 4644
rect 27157 4641 27169 4644
rect 27203 4641 27215 4675
rect 27157 4635 27215 4641
rect 27246 4632 27252 4684
rect 27304 4672 27310 4684
rect 27341 4675 27399 4681
rect 27341 4672 27353 4675
rect 27304 4644 27353 4672
rect 27304 4632 27310 4644
rect 27341 4641 27353 4644
rect 27387 4641 27399 4675
rect 27341 4635 27399 4641
rect 27614 4632 27620 4684
rect 27672 4672 27678 4684
rect 28092 4681 28120 4712
rect 27893 4675 27951 4681
rect 27893 4672 27905 4675
rect 27672 4644 27905 4672
rect 27672 4632 27678 4644
rect 27893 4641 27905 4644
rect 27939 4641 27951 4675
rect 27893 4635 27951 4641
rect 28077 4675 28135 4681
rect 28077 4641 28089 4675
rect 28123 4641 28135 4675
rect 28077 4635 28135 4641
rect 23523 4576 24164 4604
rect 24213 4607 24271 4613
rect 23523 4573 23535 4576
rect 23477 4567 23535 4573
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 23216 4536 23244 4564
rect 22066 4508 23244 4536
rect 23308 4536 23336 4567
rect 23566 4536 23572 4548
rect 23308 4508 23572 4536
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 24228 4536 24256 4567
rect 24394 4564 24400 4616
rect 24452 4564 24458 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 23952 4508 24256 4536
rect 22097 4471 22155 4477
rect 22097 4468 22109 4471
rect 20079 4440 22109 4468
rect 19521 4431 19579 4437
rect 22097 4437 22109 4440
rect 22143 4437 22155 4471
rect 22097 4431 22155 4437
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 23952 4468 23980 4508
rect 24302 4496 24308 4548
rect 24360 4536 24366 4548
rect 24596 4536 24624 4567
rect 24854 4564 24860 4616
rect 24912 4564 24918 4616
rect 24946 4564 24952 4616
rect 25004 4604 25010 4616
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 25004 4576 25329 4604
rect 25004 4564 25010 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 25409 4607 25467 4613
rect 25409 4573 25421 4607
rect 25455 4573 25467 4607
rect 25409 4567 25467 4573
rect 24360 4508 24624 4536
rect 24360 4496 24366 4508
rect 23348 4440 23980 4468
rect 24872 4468 24900 4564
rect 25424 4536 25452 4567
rect 25498 4564 25504 4616
rect 25556 4604 25562 4616
rect 25593 4607 25651 4613
rect 25593 4604 25605 4607
rect 25556 4576 25605 4604
rect 25556 4564 25562 4576
rect 25593 4573 25605 4576
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 26142 4564 26148 4616
rect 26200 4564 26206 4616
rect 26326 4564 26332 4616
rect 26384 4564 26390 4616
rect 26786 4564 26792 4616
rect 26844 4604 26850 4616
rect 26881 4607 26939 4613
rect 26881 4604 26893 4607
rect 26844 4576 26893 4604
rect 26844 4564 26850 4576
rect 26881 4573 26893 4576
rect 26927 4573 26939 4607
rect 26881 4567 26939 4573
rect 27614 4536 27620 4548
rect 25424 4508 27620 4536
rect 27614 4496 27620 4508
rect 27672 4536 27678 4548
rect 27801 4539 27859 4545
rect 27801 4536 27813 4539
rect 27672 4508 27813 4536
rect 27672 4496 27678 4508
rect 27801 4505 27813 4508
rect 27847 4505 27859 4539
rect 27801 4499 27859 4505
rect 25133 4471 25191 4477
rect 25133 4468 25145 4471
rect 24872 4440 25145 4468
rect 23348 4428 23354 4440
rect 25133 4437 25145 4440
rect 25179 4437 25191 4471
rect 25133 4431 25191 4437
rect 25406 4428 25412 4480
rect 25464 4468 25470 4480
rect 26234 4468 26240 4480
rect 25464 4440 26240 4468
rect 25464 4428 25470 4440
rect 26234 4428 26240 4440
rect 26292 4468 26298 4480
rect 26786 4468 26792 4480
rect 26292 4440 26792 4468
rect 26292 4428 26298 4440
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 4246 4224 4252 4276
rect 4304 4224 4310 4276
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 4764 4236 5273 4264
rect 4764 4224 4770 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 5442 4224 5448 4276
rect 5500 4224 5506 4276
rect 5810 4224 5816 4276
rect 5868 4224 5874 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7009 4267 7067 4273
rect 7009 4264 7021 4267
rect 6972 4236 7021 4264
rect 6972 4224 6978 4236
rect 7009 4233 7021 4236
rect 7055 4233 7067 4267
rect 11149 4267 11207 4273
rect 7009 4227 7067 4233
rect 7116 4236 9674 4264
rect 5552 4168 5764 4196
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 1394 3884 1400 3936
rect 1452 3884 1458 3936
rect 1596 3924 1624 4091
rect 2130 4088 2136 4140
rect 2188 4088 2194 4140
rect 2400 4131 2458 4137
rect 2400 4097 2412 4131
rect 2446 4128 2458 4131
rect 3234 4128 3240 4140
rect 2446 4100 3240 4128
rect 2446 4097 2458 4100
rect 2400 4091 2458 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4525 4131 4583 4137
rect 3743 4100 4476 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 3712 3992 3740 4091
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 4448 4060 4476 4100
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4982 4128 4988 4140
rect 4571 4100 4988 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5184 4060 5212 4091
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5552 4128 5580 4168
rect 5500 4100 5580 4128
rect 5500 4088 5506 4100
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5736 4137 5764 4168
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5828 4128 5856 4224
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 7116 4196 7144 4236
rect 6788 4168 7144 4196
rect 9646 4196 9674 4236
rect 11149 4233 11161 4267
rect 11195 4233 11207 4267
rect 11149 4227 11207 4233
rect 11164 4196 11192 4227
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13173 4267 13231 4273
rect 13173 4264 13185 4267
rect 13136 4236 13185 4264
rect 13136 4224 13142 4236
rect 13173 4233 13185 4236
rect 13219 4233 13231 4267
rect 13173 4227 13231 4233
rect 13354 4224 13360 4276
rect 13412 4264 13418 4276
rect 13412 4236 13492 4264
rect 13412 4224 13418 4236
rect 13464 4205 13492 4236
rect 16206 4224 16212 4276
rect 16264 4224 16270 4276
rect 17405 4267 17463 4273
rect 17405 4233 17417 4267
rect 17451 4264 17463 4267
rect 19702 4264 19708 4276
rect 17451 4236 19708 4264
rect 17451 4233 17463 4236
rect 17405 4227 17463 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 19812 4236 21312 4264
rect 13449 4199 13507 4205
rect 9646 4168 9996 4196
rect 11164 4168 11468 4196
rect 6788 4156 6794 4168
rect 8113 4140 8171 4141
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 5828 4100 6193 4128
rect 5721 4091 5779 4097
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 8110 4088 8116 4140
rect 8168 4132 8174 4140
rect 8168 4104 8209 4132
rect 8168 4088 8174 4104
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 9968 4137 9996 4168
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 8389 4091 8447 4097
rect 8864 4100 9873 4128
rect 4448 4032 5212 4060
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5408 4032 6377 4060
rect 5408 4020 5414 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6549 4063 6607 4069
rect 6549 4029 6561 4063
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 3559 3964 3740 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 4798 3952 4804 4004
rect 4856 3952 4862 4004
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6564 3992 6592 4023
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 7101 4063 7159 4069
rect 7101 4060 7113 4063
rect 6696 4032 7113 4060
rect 6696 4020 6702 4032
rect 7101 4029 7113 4032
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7282 4020 7288 4072
rect 7340 4020 7346 4072
rect 8202 4020 8208 4072
rect 8260 4020 8266 4072
rect 8864 4060 8892 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 8312 4032 8892 4060
rect 8941 4063 8999 4069
rect 6043 3964 6592 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 7469 3995 7527 4001
rect 7469 3992 7481 3995
rect 7064 3964 7481 3992
rect 7064 3952 7070 3964
rect 7469 3961 7481 3964
rect 7515 3961 7527 3995
rect 7469 3955 7527 3961
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8312 3992 8340 4032
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 8956 3992 8984 4023
rect 9122 4020 9128 4072
rect 9180 4020 9186 4072
rect 7975 3964 8340 3992
rect 8404 3964 8984 3992
rect 9968 3992 9996 4091
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 10192 4100 10241 4128
rect 10192 4088 10198 4100
rect 10229 4097 10241 4100
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 11238 4088 11244 4140
rect 11296 4088 11302 4140
rect 11330 4088 11336 4140
rect 11388 4088 11394 4140
rect 11440 4128 11468 4168
rect 13449 4165 13461 4199
rect 13495 4165 13507 4199
rect 13449 4159 13507 4165
rect 13538 4156 13544 4208
rect 13596 4196 13602 4208
rect 13596 4168 15424 4196
rect 13596 4156 13602 4168
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11440 4100 11713 4128
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 12060 4131 12118 4137
rect 12060 4097 12072 4131
rect 12106 4128 12118 4131
rect 15286 4128 15292 4140
rect 12106 4100 13216 4128
rect 12106 4097 12118 4100
rect 12060 4091 12118 4097
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10091 4032 10425 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 10502 4020 10508 4072
rect 10560 4020 10566 4072
rect 11256 4060 11284 4088
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11256 4032 11805 4060
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 10520 3992 10548 4020
rect 9968 3964 10548 3992
rect 13188 3992 13216 4100
rect 15120 4100 15292 4128
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13722 4060 13728 4072
rect 13311 4032 13728 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 15120 4060 15148 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15396 4128 15424 4168
rect 17954 4156 17960 4208
rect 18012 4156 18018 4208
rect 19150 4156 19156 4208
rect 19208 4196 19214 4208
rect 19812 4196 19840 4236
rect 20254 4196 20260 4208
rect 19208 4168 19840 4196
rect 19904 4168 20260 4196
rect 19208 4156 19214 4168
rect 16114 4128 16120 4140
rect 15396 4100 16120 4128
rect 13872 4032 15148 4060
rect 15197 4063 15255 4069
rect 13872 4020 13878 4032
rect 15197 4029 15209 4063
rect 15243 4060 15255 4063
rect 15396 4060 15424 4100
rect 16114 4088 16120 4100
rect 16172 4128 16178 4140
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 16172 4100 17601 4128
rect 16172 4088 16178 4100
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 19518 4128 19524 4140
rect 19168 4100 19524 4128
rect 15243 4032 15424 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 16758 4020 16764 4072
rect 16816 4020 16822 4072
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 18046 4060 18052 4072
rect 17911 4032 18052 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 19168 4060 19196 4100
rect 19518 4088 19524 4100
rect 19576 4088 19582 4140
rect 19904 4137 19932 4168
rect 20254 4156 20260 4168
rect 20312 4156 20318 4208
rect 21174 4156 21180 4208
rect 21232 4156 21238 4208
rect 21284 4196 21312 4236
rect 21450 4224 21456 4276
rect 21508 4264 21514 4276
rect 24302 4264 24308 4276
rect 21508 4236 24308 4264
rect 21508 4224 21514 4236
rect 24302 4224 24308 4236
rect 24360 4224 24366 4276
rect 24394 4224 24400 4276
rect 24452 4264 24458 4276
rect 24673 4267 24731 4273
rect 24673 4264 24685 4267
rect 24452 4236 24685 4264
rect 24452 4224 24458 4236
rect 24673 4233 24685 4236
rect 24719 4233 24731 4267
rect 24673 4227 24731 4233
rect 24762 4224 24768 4276
rect 24820 4224 24826 4276
rect 24872 4236 25544 4264
rect 24872 4196 24900 4236
rect 25516 4208 25544 4236
rect 27614 4224 27620 4276
rect 27672 4264 27678 4276
rect 27709 4267 27767 4273
rect 27709 4264 27721 4267
rect 27672 4236 27721 4264
rect 27672 4224 27678 4236
rect 27709 4233 27721 4236
rect 27755 4233 27767 4267
rect 27709 4227 27767 4233
rect 21284 4168 24900 4196
rect 25498 4156 25504 4208
rect 25556 4156 25562 4208
rect 26804 4168 28212 4196
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 18340 4032 19196 4060
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 13188 3964 15853 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 4246 3924 4252 3936
rect 1596 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 8404 3924 8432 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 18340 3992 18368 4032
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 19628 4060 19656 4091
rect 19978 4088 19984 4140
rect 20036 4088 20042 4140
rect 20156 4131 20214 4137
rect 20156 4097 20168 4131
rect 20202 4128 20214 4131
rect 21192 4128 21220 4156
rect 26804 4140 26832 4168
rect 20202 4100 21220 4128
rect 20202 4097 20214 4100
rect 20156 4091 20214 4097
rect 21542 4088 21548 4140
rect 21600 4088 21606 4140
rect 22088 4131 22146 4137
rect 22088 4097 22100 4131
rect 22134 4128 22146 4131
rect 22134 4100 23060 4128
rect 22134 4097 22146 4100
rect 22088 4091 22146 4097
rect 19996 4060 20024 4088
rect 19628 4032 20024 4060
rect 21821 4063 21879 4069
rect 21821 4029 21833 4063
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 15841 3955 15899 3961
rect 17236 3964 18368 3992
rect 18417 3995 18475 4001
rect 6512 3896 8432 3924
rect 6512 3884 6518 3896
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 10594 3924 10600 3936
rect 9916 3896 10600 3924
rect 9916 3884 9922 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 12526 3924 12532 3936
rect 11563 3896 12532 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 17236 3924 17264 3964
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 19334 3992 19340 4004
rect 18463 3964 19340 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 21269 3995 21327 4001
rect 21269 3961 21281 3995
rect 21315 3992 21327 3995
rect 21315 3964 21496 3992
rect 21315 3961 21327 3964
rect 21269 3955 21327 3961
rect 21468 3936 21496 3964
rect 15712 3896 17264 3924
rect 15712 3884 15718 3896
rect 17310 3884 17316 3936
rect 17368 3884 17374 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 18506 3924 18512 3936
rect 17460 3896 18512 3924
rect 17460 3884 17466 3896
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 20622 3924 20628 3936
rect 19475 3896 20628 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 21358 3884 21364 3936
rect 21416 3884 21422 3936
rect 21450 3884 21456 3936
rect 21508 3884 21514 3936
rect 21836 3924 21864 4023
rect 23032 3992 23060 4100
rect 23382 4088 23388 4140
rect 23440 4128 23446 4140
rect 24949 4131 25007 4137
rect 24949 4128 24961 4131
rect 23440 4100 24961 4128
rect 23440 4088 23446 4100
rect 24949 4097 24961 4100
rect 24995 4097 25007 4131
rect 24949 4091 25007 4097
rect 25130 4088 25136 4140
rect 25188 4128 25194 4140
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 25188 4100 25237 4128
rect 25188 4088 25194 4100
rect 25225 4097 25237 4100
rect 25271 4128 25283 4131
rect 25406 4128 25412 4140
rect 25271 4100 25412 4128
rect 25271 4097 25283 4100
rect 25225 4091 25283 4097
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 25682 4088 25688 4140
rect 25740 4088 25746 4140
rect 26786 4088 26792 4140
rect 26844 4088 26850 4140
rect 26970 4088 26976 4140
rect 27028 4128 27034 4140
rect 27249 4131 27307 4137
rect 27249 4128 27261 4131
rect 27028 4100 27261 4128
rect 27028 4088 27034 4100
rect 27249 4097 27261 4100
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 27706 4088 27712 4140
rect 27764 4088 27770 4140
rect 28184 4137 28212 4168
rect 28169 4131 28227 4137
rect 28169 4097 28181 4131
rect 28215 4097 28227 4131
rect 28169 4091 28227 4097
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4060 23351 4063
rect 23658 4060 23664 4072
rect 23339 4032 23664 4060
rect 23339 4029 23351 4032
rect 23293 4023 23351 4029
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 24026 4020 24032 4072
rect 24084 4020 24090 4072
rect 24210 4020 24216 4072
rect 24268 4020 24274 4072
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 25317 4063 25375 4069
rect 25317 4060 25329 4063
rect 24912 4032 25329 4060
rect 24912 4020 24918 4032
rect 25317 4029 25329 4032
rect 25363 4029 25375 4063
rect 25317 4023 25375 4029
rect 23937 3995 23995 4001
rect 23937 3992 23949 3995
rect 23032 3964 23949 3992
rect 23937 3961 23949 3964
rect 23983 3961 23995 3995
rect 23937 3955 23995 3961
rect 25041 3995 25099 4001
rect 25041 3961 25053 3995
rect 25087 3992 25099 3995
rect 25700 3992 25728 4088
rect 25774 4020 25780 4072
rect 25832 4060 25838 4072
rect 26053 4063 26111 4069
rect 26053 4060 26065 4063
rect 25832 4032 26065 4060
rect 25832 4020 25838 4032
rect 26053 4029 26065 4032
rect 26099 4029 26111 4063
rect 26053 4023 26111 4029
rect 26142 4020 26148 4072
rect 26200 4020 26206 4072
rect 26237 4063 26295 4069
rect 26237 4029 26249 4063
rect 26283 4060 26295 4063
rect 26326 4060 26332 4072
rect 26283 4032 26332 4060
rect 26283 4029 26295 4032
rect 26237 4023 26295 4029
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 26510 4020 26516 4072
rect 26568 4060 26574 4072
rect 27065 4063 27123 4069
rect 27065 4060 27077 4063
rect 26568 4032 27077 4060
rect 26568 4020 26574 4032
rect 27065 4029 27077 4032
rect 27111 4029 27123 4063
rect 27724 4060 27752 4088
rect 28261 4063 28319 4069
rect 28261 4060 28273 4063
rect 27724 4032 28273 4060
rect 27065 4023 27123 4029
rect 28261 4029 28273 4032
rect 28307 4029 28319 4063
rect 28261 4023 28319 4029
rect 25087 3964 25728 3992
rect 26160 3992 26188 4020
rect 26421 3995 26479 4001
rect 26421 3992 26433 3995
rect 26160 3964 26433 3992
rect 25087 3961 25099 3964
rect 25041 3955 25099 3961
rect 26421 3961 26433 3964
rect 26467 3961 26479 3995
rect 27080 3992 27108 4023
rect 27985 3995 28043 4001
rect 27985 3992 27997 3995
rect 27080 3964 27997 3992
rect 26421 3955 26479 3961
rect 27985 3961 27997 3964
rect 28031 3961 28043 3995
rect 27985 3955 28043 3961
rect 22738 3924 22744 3936
rect 21836 3896 22744 3924
rect 22738 3884 22744 3896
rect 22796 3884 22802 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 23382 3924 23388 3936
rect 23256 3896 23388 3924
rect 23256 3884 23262 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 25188 3896 25973 3924
rect 25188 3884 25194 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 25961 3887 26019 3893
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 3142 3720 3148 3732
rect 1903 3692 3148 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 4338 3680 4344 3732
rect 4396 3680 4402 3732
rect 4525 3723 4583 3729
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 5350 3720 5356 3732
rect 4571 3692 5356 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3720 5503 3723
rect 7282 3720 7288 3732
rect 5491 3692 7288 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8260 3692 8585 3720
rect 8260 3680 8266 3692
rect 8573 3689 8585 3692
rect 8619 3720 8631 3723
rect 9306 3720 9312 3732
rect 8619 3692 9312 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 12434 3720 12440 3732
rect 11808 3692 12440 3720
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 4356 3652 4384 3680
rect 2179 3624 4384 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 4706 3612 4712 3664
rect 4764 3652 4770 3664
rect 5166 3652 5172 3664
rect 4764 3624 5172 3652
rect 4764 3612 4770 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 5721 3655 5779 3661
rect 5721 3652 5733 3655
rect 5684 3624 5733 3652
rect 5684 3612 5690 3624
rect 5721 3621 5733 3624
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 5994 3612 6000 3664
rect 6052 3612 6058 3664
rect 6273 3655 6331 3661
rect 6273 3621 6285 3655
rect 6319 3652 6331 3655
rect 6319 3624 8156 3652
rect 6319 3621 6331 3624
rect 6273 3615 6331 3621
rect 2593 3587 2651 3593
rect 2593 3584 2605 3587
rect 1504 3556 2605 3584
rect 1504 3525 1532 3556
rect 2593 3553 2605 3556
rect 2639 3553 2651 3587
rect 2593 3547 2651 3553
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 6638 3584 6644 3596
rect 3559 3556 6644 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1728 3488 1777 3516
rect 1728 3476 1734 3488
rect 1765 3485 1777 3488
rect 1811 3516 1823 3519
rect 1854 3516 1860 3528
rect 1811 3488 1860 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 2004 3488 2053 3516
rect 2004 3476 2010 3488
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2498 3476 2504 3528
rect 2556 3476 2562 3528
rect 2608 3518 2636 3547
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 8128 3593 8156 3624
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 6963 3556 7941 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7929 3553 7941 3556
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3584 9459 3587
rect 9692 3584 9720 3680
rect 11808 3661 11836 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12802 3680 12808 3732
rect 12860 3680 12866 3732
rect 13814 3720 13820 3732
rect 12912 3692 13820 3720
rect 11333 3655 11391 3661
rect 11333 3621 11345 3655
rect 11379 3652 11391 3655
rect 11793 3655 11851 3661
rect 11793 3652 11805 3655
rect 11379 3624 11805 3652
rect 11379 3621 11391 3624
rect 11333 3615 11391 3621
rect 11793 3621 11805 3624
rect 11839 3621 11851 3655
rect 12912 3652 12940 3692
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14090 3680 14096 3732
rect 14148 3680 14154 3732
rect 16758 3720 16764 3732
rect 14200 3692 16764 3720
rect 11793 3615 11851 3621
rect 12406 3624 12940 3652
rect 12989 3655 13047 3661
rect 9447 3556 9720 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 12406 3584 12434 3624
rect 12989 3621 13001 3655
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 11756 3556 12434 3584
rect 13004 3584 13032 3615
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14200 3652 14228 3692
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17218 3720 17224 3732
rect 16899 3692 17224 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 19610 3680 19616 3732
rect 19668 3720 19674 3732
rect 21358 3720 21364 3732
rect 19668 3692 21364 3720
rect 19668 3680 19674 3692
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 21450 3680 21456 3732
rect 21508 3720 21514 3732
rect 21508 3692 22223 3720
rect 21508 3680 21514 3692
rect 14056 3624 14228 3652
rect 15749 3655 15807 3661
rect 14056 3612 14062 3624
rect 15749 3621 15761 3655
rect 15795 3652 15807 3655
rect 15795 3624 16068 3652
rect 15795 3621 15807 3624
rect 15749 3615 15807 3621
rect 13004 3556 14320 3584
rect 11756 3544 11762 3556
rect 2608 3516 2774 3518
rect 3234 3516 3240 3528
rect 2608 3490 3240 3516
rect 2746 3488 3240 3490
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3418 3476 3424 3528
rect 3476 3476 3482 3528
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3660 3488 3893 3516
rect 3660 3476 3666 3488
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4304 3488 4721 3516
rect 4304 3476 4310 3488
rect 4709 3485 4721 3488
rect 4755 3516 4767 3519
rect 4755 3488 5580 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 3142 3448 3148 3460
rect 1627 3420 3148 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 3142 3408 3148 3420
rect 3200 3408 3206 3460
rect 5166 3408 5172 3460
rect 5224 3408 5230 3460
rect 5552 3448 5580 3488
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5776 3488 5917 3516
rect 5776 3476 5782 3488
rect 5905 3485 5917 3488
rect 5951 3516 5963 3519
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5951 3488 6193 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6181 3485 6193 3488
rect 6227 3516 6239 3519
rect 6270 3516 6276 3528
rect 6227 3488 6276 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6748 3516 6776 3544
rect 6595 3488 6776 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 5736 3448 5764 3476
rect 5552 3420 5764 3448
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 6472 3448 6500 3479
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6932 3488 7113 3516
rect 6052 3420 6500 3448
rect 6052 3408 6058 3420
rect 6638 3408 6644 3460
rect 6696 3408 6702 3460
rect 2314 3340 2320 3392
rect 2372 3340 2378 3392
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 6932 3380 6960 3488
rect 7101 3485 7113 3488
rect 7147 3516 7159 3519
rect 8662 3516 8668 3528
rect 7147 3488 8668 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3516 9091 3519
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 9079 3488 9229 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 8956 3448 8984 3479
rect 9674 3448 9680 3460
rect 8956 3420 9680 3448
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 9968 3448 9996 3479
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10100 3488 10701 3516
rect 10100 3476 10106 3488
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 10870 3476 10876 3528
rect 10928 3476 10934 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 13078 3516 13084 3528
rect 12299 3488 13084 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 10318 3448 10324 3460
rect 9968 3420 10324 3448
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11624 3448 11652 3479
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14182 3516 14188 3528
rect 13403 3488 14188 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 11204 3420 11652 3448
rect 13188 3448 13216 3479
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14292 3525 14320 3556
rect 16040 3528 16068 3624
rect 16666 3612 16672 3664
rect 16724 3612 16730 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 20622 3652 20628 3664
rect 18748 3624 20628 3652
rect 18748 3612 18754 3624
rect 20622 3612 20628 3624
rect 20680 3612 20686 3664
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14415 3488 15884 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 13538 3448 13544 3460
rect 13188 3420 13544 3448
rect 11204 3408 11210 3420
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 13909 3451 13967 3457
rect 13909 3417 13921 3451
rect 13955 3448 13967 3451
rect 14614 3451 14672 3457
rect 14614 3448 14626 3451
rect 13955 3420 14626 3448
rect 13955 3417 13967 3420
rect 13909 3411 13967 3417
rect 14614 3417 14626 3420
rect 14660 3417 14672 3451
rect 15856 3448 15884 3488
rect 16022 3476 16028 3528
rect 16080 3476 16086 3528
rect 16684 3525 16712 3612
rect 19426 3584 19432 3596
rect 18248 3556 19432 3584
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 16908 3488 17141 3516
rect 16908 3476 16914 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3516 17279 3519
rect 18248 3516 18276 3556
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 19705 3587 19763 3593
rect 19705 3584 19717 3587
rect 19576 3556 19717 3584
rect 19576 3544 19582 3556
rect 19705 3553 19717 3556
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 20312 3556 21189 3584
rect 20312 3544 20318 3556
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 22195 3584 22223 3692
rect 24302 3680 24308 3732
rect 24360 3680 24366 3732
rect 24394 3680 24400 3732
rect 24452 3720 24458 3732
rect 24765 3723 24823 3729
rect 24765 3720 24777 3723
rect 24452 3692 24777 3720
rect 24452 3680 24458 3692
rect 24765 3689 24777 3692
rect 24811 3689 24823 3723
rect 24765 3683 24823 3689
rect 25866 3680 25872 3732
rect 25924 3680 25930 3732
rect 26142 3680 26148 3732
rect 26200 3720 26206 3732
rect 26237 3723 26295 3729
rect 26237 3720 26249 3723
rect 26200 3692 26249 3720
rect 26200 3680 26206 3692
rect 26237 3689 26249 3692
rect 26283 3689 26295 3723
rect 26237 3683 26295 3689
rect 26602 3680 26608 3732
rect 26660 3680 26666 3732
rect 26786 3680 26792 3732
rect 26844 3720 26850 3732
rect 26973 3723 27031 3729
rect 26844 3692 26924 3720
rect 26844 3680 26850 3692
rect 22557 3655 22615 3661
rect 22557 3621 22569 3655
rect 22603 3652 22615 3655
rect 23658 3652 23664 3664
rect 22603 3624 23664 3652
rect 22603 3621 22615 3624
rect 22557 3615 22615 3621
rect 23658 3612 23664 3624
rect 23716 3612 23722 3664
rect 23934 3652 23940 3664
rect 23760 3624 23940 3652
rect 22195 3556 22784 3584
rect 21177 3547 21235 3553
rect 18966 3516 18972 3528
rect 17267 3488 18276 3516
rect 18524 3488 18972 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 16758 3448 16764 3460
rect 15856 3420 16764 3448
rect 14614 3411 14672 3417
rect 16758 3408 16764 3420
rect 16816 3448 16822 3460
rect 17236 3448 17264 3479
rect 16816 3420 17264 3448
rect 17488 3451 17546 3457
rect 16816 3408 16822 3420
rect 17488 3417 17500 3451
rect 17534 3448 17546 3451
rect 17862 3448 17868 3460
rect 17534 3420 17868 3448
rect 17534 3417 17546 3420
rect 17488 3411 17546 3417
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 18524 3448 18552 3488
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 22756 3525 22784 3556
rect 23382 3544 23388 3596
rect 23440 3544 23446 3596
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3516 22799 3519
rect 23760 3516 23788 3624
rect 23934 3612 23940 3624
rect 23992 3612 23998 3664
rect 24320 3652 24348 3680
rect 25682 3652 25688 3664
rect 24320 3624 25688 3652
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 25884 3652 25912 3680
rect 25884 3624 26832 3652
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 23900 3556 25789 3584
rect 23900 3544 23906 3556
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 25866 3544 25872 3596
rect 25924 3544 25930 3596
rect 26050 3544 26056 3596
rect 26108 3544 26114 3596
rect 22787 3488 23788 3516
rect 22787 3485 22799 3488
rect 22741 3479 22799 3485
rect 19150 3448 19156 3460
rect 18156 3420 18552 3448
rect 18616 3420 19156 3448
rect 3476 3352 6960 3380
rect 3476 3340 3482 3352
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 16574 3340 16580 3392
rect 16632 3340 16638 3392
rect 16945 3383 17003 3389
rect 16945 3349 16957 3383
rect 16991 3380 17003 3383
rect 18156 3380 18184 3420
rect 16991 3352 18184 3380
rect 16991 3349 17003 3352
rect 16945 3343 17003 3349
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 18616 3389 18644 3420
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18288 3352 18613 3380
rect 18288 3340 18294 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 19260 3380 19288 3479
rect 24394 3476 24400 3528
rect 24452 3476 24458 3528
rect 24486 3476 24492 3528
rect 24544 3476 24550 3528
rect 24578 3476 24584 3528
rect 24636 3476 24642 3528
rect 26804 3525 26832 3624
rect 26896 3525 26924 3692
rect 26973 3689 26985 3723
rect 27019 3720 27031 3723
rect 27338 3720 27344 3732
rect 27019 3692 27344 3720
rect 27019 3689 27031 3692
rect 26973 3683 27031 3689
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 27154 3544 27160 3596
rect 27212 3544 27218 3596
rect 25133 3519 25191 3525
rect 25133 3485 25145 3519
rect 25179 3485 25191 3519
rect 25133 3479 25191 3485
rect 26789 3519 26847 3525
rect 26789 3485 26801 3519
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 26881 3519 26939 3525
rect 26881 3485 26893 3519
rect 26927 3485 26939 3519
rect 26881 3479 26939 3485
rect 19429 3451 19487 3457
rect 19429 3417 19441 3451
rect 19475 3448 19487 3451
rect 20438 3448 20444 3460
rect 19475 3420 20444 3448
rect 19475 3417 19487 3420
rect 19429 3411 19487 3417
rect 20438 3408 20444 3420
rect 20496 3408 20502 3460
rect 21444 3451 21502 3457
rect 21444 3417 21456 3451
rect 21490 3448 21502 3451
rect 24029 3451 24087 3457
rect 24029 3448 24041 3451
rect 21490 3420 24041 3448
rect 21490 3417 21502 3420
rect 21444 3411 21502 3417
rect 24029 3417 24041 3420
rect 24075 3417 24087 3451
rect 24504 3448 24532 3476
rect 24670 3448 24676 3460
rect 24504 3420 24676 3448
rect 24029 3411 24087 3417
rect 24670 3408 24676 3420
rect 24728 3448 24734 3460
rect 25148 3448 25176 3479
rect 24728 3420 25176 3448
rect 27424 3451 27482 3457
rect 24728 3408 24734 3420
rect 27424 3417 27436 3451
rect 27470 3448 27482 3451
rect 27982 3448 27988 3460
rect 27470 3420 27988 3448
rect 27470 3417 27482 3420
rect 27424 3411 27482 3417
rect 27982 3408 27988 3420
rect 28040 3408 28046 3460
rect 19334 3380 19340 3392
rect 19260 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3380 19398 3392
rect 20346 3380 20352 3392
rect 19392 3352 20352 3380
rect 19392 3340 19398 3352
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 21324 3352 23305 3380
rect 21324 3340 21330 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23293 3343 23351 3349
rect 25682 3340 25688 3392
rect 25740 3380 25746 3392
rect 28537 3383 28595 3389
rect 28537 3380 28549 3383
rect 25740 3352 28549 3380
rect 25740 3340 25746 3352
rect 28537 3349 28549 3352
rect 28583 3349 28595 3383
rect 28537 3343 28595 3349
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 3234 3176 3240 3188
rect 2056 3148 3240 3176
rect 2056 3108 2084 3148
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3384 3148 4077 3176
rect 3384 3136 3390 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 5258 3176 5264 3188
rect 4571 3148 5264 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6454 3136 6460 3188
rect 6512 3136 6518 3188
rect 7742 3136 7748 3188
rect 7800 3136 7806 3188
rect 8570 3176 8576 3188
rect 7852 3148 8576 3176
rect 1412 3080 2084 3108
rect 1412 3049 1440 3080
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3040 1823 3043
rect 1811 3012 1992 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 1535 2944 1900 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 1872 2836 1900 2944
rect 1964 2904 1992 3012
rect 2056 2981 2084 3080
rect 2130 3068 2136 3120
rect 2188 3108 2194 3120
rect 5068 3111 5126 3117
rect 2188 3080 4844 3108
rect 2188 3068 2194 3080
rect 2608 3040 2636 3080
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2608 3012 2697 3040
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2941 3043 2999 3049
rect 2941 3040 2953 3043
rect 2685 3003 2743 3009
rect 2792 3012 2953 3040
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2941 2099 2975
rect 2041 2935 2099 2941
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 2792 2972 2820 3012
rect 2941 3009 2953 3012
rect 2987 3009 2999 3043
rect 2941 3003 2999 3009
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4522 3040 4528 3052
rect 4295 3012 4528 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4706 3000 4712 3052
rect 4764 3000 4770 3052
rect 4816 3049 4844 3080
rect 5068 3077 5080 3111
rect 5114 3108 5126 3111
rect 7760 3108 7788 3136
rect 5114 3080 7788 3108
rect 5114 3077 5126 3080
rect 5068 3071 5126 3077
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6411 3012 6745 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6733 3009 6745 3012
rect 6779 3040 6791 3043
rect 7852 3040 7880 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 8720 3148 9505 3176
rect 8720 3136 8726 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11480 3148 11805 3176
rect 11480 3136 11486 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 13998 3176 14004 3188
rect 11793 3139 11851 3145
rect 12084 3148 14004 3176
rect 8202 3108 8208 3120
rect 8128 3080 8208 3108
rect 6779 3012 7880 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 8018 3000 8024 3052
rect 8076 3000 8082 3052
rect 8128 3049 8156 3080
rect 8202 3068 8208 3080
rect 8260 3108 8266 3120
rect 8260 3080 12020 3108
rect 8260 3068 8266 3080
rect 9784 3049 9812 3080
rect 11256 3052 11284 3080
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3009 8171 3043
rect 8369 3043 8427 3049
rect 8369 3040 8381 3043
rect 8113 3003 8171 3009
rect 8220 3012 8381 3040
rect 2639 2944 2820 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 4080 2904 4108 3000
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6880 2944 7389 2972
rect 6880 2932 6886 2944
rect 1964 2876 2636 2904
rect 2498 2836 2504 2848
rect 1872 2808 2504 2836
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 2608 2836 2636 2876
rect 3620 2876 4108 2904
rect 3620 2836 3648 2876
rect 4338 2864 4344 2916
rect 4396 2864 4402 2916
rect 4448 2876 4844 2904
rect 2608 2808 3648 2836
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4448 2836 4476 2876
rect 4212 2808 4476 2836
rect 4816 2836 4844 2876
rect 5442 2836 5448 2848
rect 4816 2808 5448 2836
rect 4212 2796 4218 2808
rect 5442 2796 5448 2808
rect 5500 2836 5506 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5500 2808 6193 2836
rect 5500 2796 5506 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 7208 2836 7236 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 8220 2972 8248 3012
rect 8369 3009 8381 3012
rect 8415 3009 8427 3043
rect 8369 3003 8427 3009
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10036 3043 10094 3049
rect 10036 3009 10048 3043
rect 10082 3040 10094 3043
rect 10594 3040 10600 3052
rect 10082 3012 10600 3040
rect 10082 3009 10094 3012
rect 10036 3003 10094 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11238 3000 11244 3052
rect 11296 3000 11302 3052
rect 11992 3049 12020 3080
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 7377 2935 7435 2941
rect 7944 2944 8248 2972
rect 11716 2972 11744 3003
rect 12084 2972 12112 3148
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 14240 3148 14841 3176
rect 14240 3136 14246 3148
rect 14829 3145 14841 3148
rect 14875 3176 14887 3179
rect 14918 3176 14924 3188
rect 14875 3148 14924 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 16172 3148 16313 3176
rect 16172 3136 16178 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16301 3139 16359 3145
rect 17402 3136 17408 3188
rect 17460 3136 17466 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 17770 3176 17776 3188
rect 17543 3148 17776 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 18690 3176 18696 3188
rect 18104 3148 18696 3176
rect 18104 3136 18110 3148
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 18782 3136 18788 3188
rect 18840 3136 18846 3188
rect 19168 3148 20392 3176
rect 12244 3111 12302 3117
rect 12244 3077 12256 3111
rect 12290 3108 12302 3111
rect 12342 3108 12348 3120
rect 12290 3080 12348 3108
rect 12290 3077 12302 3080
rect 12244 3071 12302 3077
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 16758 3108 16764 3120
rect 13464 3080 16764 3108
rect 13464 3049 13492 3080
rect 14936 3049 14964 3080
rect 16758 3068 16764 3080
rect 16816 3068 16822 3120
rect 18800 3108 18828 3136
rect 19168 3120 19196 3148
rect 17604 3080 18828 3108
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 13716 3043 13774 3049
rect 13716 3009 13728 3043
rect 13762 3040 13774 3043
rect 14921 3043 14979 3049
rect 13762 3012 14872 3040
rect 13762 3009 13774 3012
rect 13716 3003 13774 3009
rect 11716 2944 12112 2972
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 7944 2904 7972 2944
rect 7331 2876 7972 2904
rect 14844 2904 14872 3012
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15188 3043 15246 3049
rect 15188 3009 15200 3043
rect 15234 3040 15246 3043
rect 16574 3040 16580 3052
rect 15234 3012 16580 3040
rect 15234 3009 15246 3012
rect 15188 3003 15246 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 17604 3040 17632 3080
rect 19150 3068 19156 3120
rect 19208 3068 19214 3120
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19889 3111 19947 3117
rect 19889 3108 19901 3111
rect 19484 3080 19901 3108
rect 19484 3068 19490 3080
rect 19889 3077 19901 3080
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 20162 3068 20168 3120
rect 20220 3068 20226 3120
rect 20364 3108 20392 3148
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 21545 3179 21603 3185
rect 21545 3176 21557 3179
rect 20496 3148 21557 3176
rect 20496 3136 20502 3148
rect 21545 3145 21557 3148
rect 21591 3145 21603 3179
rect 22646 3176 22652 3188
rect 21545 3139 21603 3145
rect 21928 3148 22652 3176
rect 20364 3080 21496 3108
rect 16776 3012 17632 3040
rect 17681 3043 17739 3049
rect 16776 2981 16804 3012
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3009 18015 3043
rect 17957 3003 18015 3009
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 16942 2932 16948 2984
rect 17000 2932 17006 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 17696 2972 17724 3003
rect 17644 2944 17724 2972
rect 17644 2932 17650 2944
rect 17972 2904 18000 3003
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 20180 3040 20208 3068
rect 20027 3012 20208 3040
rect 20248 3043 20306 3049
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20248 3009 20260 3043
rect 20294 3040 20306 3043
rect 21266 3040 21272 3052
rect 20294 3012 21272 3040
rect 20294 3009 20306 3012
rect 20248 3003 20306 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 21468 3049 21496 3080
rect 21928 3049 21956 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23750 3136 23756 3188
rect 23808 3136 23814 3188
rect 23842 3136 23848 3188
rect 23900 3136 23906 3188
rect 24854 3136 24860 3188
rect 24912 3176 24918 3188
rect 26789 3179 26847 3185
rect 26789 3176 26801 3179
rect 24912 3148 26801 3176
rect 24912 3136 24918 3148
rect 26789 3145 26801 3148
rect 26835 3145 26847 3179
rect 26789 3139 26847 3145
rect 27154 3136 27160 3188
rect 27212 3136 27218 3188
rect 23860 3108 23888 3136
rect 23492 3080 23888 3108
rect 23952 3080 25452 3108
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3009 21971 3043
rect 21913 3003 21971 3009
rect 22180 3043 22238 3049
rect 23492 3044 23520 3080
rect 22180 3009 22192 3043
rect 22226 3040 22238 3043
rect 23308 3040 23520 3044
rect 22226 3016 23520 3040
rect 23569 3043 23627 3049
rect 22226 3012 23336 3016
rect 22226 3009 22238 3012
rect 22180 3003 22238 3009
rect 23569 3009 23581 3043
rect 23615 3009 23627 3043
rect 23569 3003 23627 3009
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2972 18291 2975
rect 19794 2972 19800 2984
rect 18279 2944 19800 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 19978 2904 19984 2916
rect 14844 2876 14964 2904
rect 17972 2876 19984 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 7208 2808 11161 2836
rect 6181 2799 6239 2805
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 13354 2796 13360 2848
rect 13412 2796 13418 2848
rect 14936 2836 14964 2876
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 20990 2864 20996 2916
rect 21048 2904 21054 2916
rect 21361 2907 21419 2913
rect 21361 2904 21373 2907
rect 21048 2876 21373 2904
rect 21048 2864 21054 2876
rect 21361 2873 21373 2876
rect 21407 2873 21419 2907
rect 21361 2867 21419 2873
rect 15286 2836 15292 2848
rect 14936 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 17773 2839 17831 2845
rect 17773 2805 17785 2839
rect 17819 2836 17831 2839
rect 18138 2836 18144 2848
rect 17819 2808 18144 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 20898 2836 20904 2848
rect 18748 2808 20904 2836
rect 18748 2796 18754 2808
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 21468 2836 21496 3003
rect 23584 2972 23612 3003
rect 23658 3000 23664 3052
rect 23716 3000 23722 3052
rect 23952 2981 23980 3080
rect 24204 3043 24262 3049
rect 24204 3009 24216 3043
rect 24250 3040 24262 3043
rect 25130 3040 25136 3052
rect 24250 3012 25136 3040
rect 24250 3009 24262 3012
rect 24204 3003 24262 3009
rect 25130 3000 25136 3012
rect 25188 3000 25194 3052
rect 25424 3049 25452 3080
rect 25409 3043 25467 3049
rect 25409 3009 25421 3043
rect 25455 3009 25467 3043
rect 25409 3003 25467 3009
rect 25676 3043 25734 3049
rect 25676 3009 25688 3043
rect 25722 3040 25734 3043
rect 26694 3040 26700 3052
rect 25722 3012 26700 3040
rect 25722 3009 25734 3012
rect 25676 3003 25734 3009
rect 23216 2944 23612 2972
rect 23937 2975 23995 2981
rect 23216 2836 23244 2944
rect 23937 2941 23949 2975
rect 23983 2941 23995 2975
rect 23937 2935 23995 2941
rect 23290 2864 23296 2916
rect 23348 2864 23354 2916
rect 21468 2808 23244 2836
rect 23382 2796 23388 2848
rect 23440 2796 23446 2848
rect 24670 2796 24676 2848
rect 24728 2836 24734 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 24728 2808 25329 2836
rect 24728 2796 24734 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25424 2836 25452 3003
rect 26694 3000 26700 3012
rect 26752 3000 26758 3052
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3040 27031 3043
rect 27172 3040 27200 3136
rect 27246 3049 27252 3052
rect 27019 3012 27200 3040
rect 27019 3009 27031 3012
rect 26973 3003 27031 3009
rect 27240 3003 27252 3049
rect 26988 2836 27016 3003
rect 27246 3000 27252 3003
rect 27304 3000 27310 3052
rect 25424 2808 27016 2836
rect 25317 2799 25375 2805
rect 27154 2796 27160 2848
rect 27212 2836 27218 2848
rect 28353 2839 28411 2845
rect 28353 2836 28365 2839
rect 27212 2808 28365 2836
rect 27212 2796 27218 2808
rect 28353 2805 28365 2808
rect 28399 2805 28411 2839
rect 28353 2799 28411 2805
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 2130 2592 2136 2644
rect 2188 2592 2194 2644
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2556 2604 3188 2632
rect 2556 2592 2562 2604
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2038 2564 2044 2576
rect 1995 2536 2044 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2038 2524 2044 2536
rect 2096 2524 2102 2576
rect 2148 2496 2176 2592
rect 3160 2564 3188 2604
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 3605 2635 3663 2641
rect 3605 2632 3617 2635
rect 3292 2604 3617 2632
rect 3292 2592 3298 2604
rect 3605 2601 3617 2604
rect 3651 2601 3663 2635
rect 3605 2595 3663 2601
rect 5350 2592 5356 2644
rect 5408 2592 5414 2644
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 8570 2592 8576 2644
rect 8628 2592 8634 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 10042 2632 10048 2644
rect 9171 2604 10048 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10376 2604 10701 2632
rect 10376 2592 10382 2604
rect 10689 2601 10701 2604
rect 10735 2601 10747 2635
rect 10689 2595 10747 2601
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10928 2604 10977 2632
rect 10928 2592 10934 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11146 2592 11152 2644
rect 11204 2592 11210 2644
rect 11256 2604 14412 2632
rect 3160 2536 4752 2564
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 2148 2468 2237 2496
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 3510 2456 3516 2508
rect 3568 2496 3574 2508
rect 4065 2499 4123 2505
rect 3568 2468 4016 2496
rect 3568 2456 3574 2468
rect 1394 2388 1400 2440
rect 1452 2428 1458 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1452 2400 1593 2428
rect 1452 2388 1458 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2130 2388 2136 2440
rect 2188 2388 2194 2440
rect 3234 2428 3240 2440
rect 2424 2400 3240 2428
rect 2424 2360 2452 2400
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3988 2428 4016 2468
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4154 2496 4160 2508
rect 4111 2468 4160 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4724 2505 4752 2536
rect 4816 2536 6592 2564
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 4816 2428 4844 2536
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6564 2505 6592 2536
rect 10410 2524 10416 2576
rect 10468 2564 10474 2576
rect 11256 2564 11284 2604
rect 10468 2536 11284 2564
rect 10468 2524 10474 2536
rect 13078 2524 13084 2576
rect 13136 2564 13142 2576
rect 14384 2564 14412 2604
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14516 2604 15025 2632
rect 14516 2592 14522 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15013 2595 15071 2601
rect 15194 2592 15200 2644
rect 15252 2592 15258 2644
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 15344 2604 16497 2632
rect 15344 2592 15350 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 18141 2635 18199 2641
rect 18141 2632 18153 2635
rect 17000 2604 18153 2632
rect 17000 2592 17006 2604
rect 18141 2601 18153 2604
rect 18187 2601 18199 2635
rect 18141 2595 18199 2601
rect 19245 2635 19303 2641
rect 19245 2601 19257 2635
rect 19291 2632 19303 2635
rect 19886 2632 19892 2644
rect 19291 2604 19892 2632
rect 19291 2601 19303 2604
rect 19245 2595 19303 2601
rect 19886 2592 19892 2604
rect 19944 2592 19950 2644
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 21269 2635 21327 2641
rect 21269 2632 21281 2635
rect 20036 2604 21281 2632
rect 20036 2592 20042 2604
rect 21269 2601 21281 2604
rect 21315 2601 21327 2635
rect 21269 2595 21327 2601
rect 24489 2635 24547 2641
rect 24489 2601 24501 2635
rect 24535 2632 24547 2635
rect 24578 2632 24584 2644
rect 24535 2604 24584 2632
rect 24535 2601 24547 2604
rect 24489 2595 24547 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 25501 2635 25559 2641
rect 24688 2604 25176 2632
rect 13136 2536 14136 2564
rect 14384 2536 16068 2564
rect 13136 2524 13142 2536
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5868 2468 6377 2496
rect 5868 2456 5874 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 8260 2468 9321 2496
rect 8260 2456 8266 2468
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11296 2468 11713 2496
rect 11296 2456 11302 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 13096 2468 13952 2496
rect 3476 2400 3832 2428
rect 3988 2400 4844 2428
rect 4893 2431 4951 2437
rect 3476 2388 3482 2400
rect 1412 2332 2452 2360
rect 2492 2363 2550 2369
rect 1412 2301 1440 2332
rect 2492 2329 2504 2363
rect 2538 2360 2550 2363
rect 3804 2360 3832 2400
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5767 2400 6193 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 6181 2397 6193 2400
rect 6227 2428 6239 2431
rect 6270 2428 6276 2440
rect 6227 2400 6276 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 4908 2360 4936 2391
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2428 7251 2431
rect 8220 2428 8248 2456
rect 7239 2400 8248 2428
rect 9033 2431 9091 2437
rect 7239 2397 7251 2400
rect 7193 2391 7251 2397
rect 9033 2397 9045 2431
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9576 2431 9634 2437
rect 9576 2397 9588 2431
rect 9622 2428 9634 2431
rect 9622 2400 10456 2428
rect 9622 2397 9634 2400
rect 9576 2391 9634 2397
rect 2538 2332 3280 2360
rect 3804 2332 4936 2360
rect 7460 2363 7518 2369
rect 2538 2329 2550 2332
rect 2492 2323 2550 2329
rect 1397 2295 1455 2301
rect 1397 2261 1409 2295
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 1765 2295 1823 2301
rect 1765 2261 1777 2295
rect 1811 2292 1823 2295
rect 3142 2292 3148 2304
rect 1811 2264 3148 2292
rect 1811 2261 1823 2264
rect 1765 2255 1823 2261
rect 3142 2252 3148 2264
rect 3200 2252 3206 2304
rect 3252 2292 3280 2332
rect 7460 2329 7472 2363
rect 7506 2360 7518 2363
rect 8018 2360 8024 2372
rect 7506 2332 8024 2360
rect 7506 2329 7518 2332
rect 7460 2323 7518 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 3252 2264 4629 2292
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 4617 2255 4675 2261
rect 5994 2252 6000 2304
rect 6052 2252 6058 2304
rect 9048 2292 9076 2391
rect 10428 2360 10456 2400
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10560 2400 10885 2428
rect 10560 2388 10566 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 13096 2428 13124 2468
rect 11440 2400 13124 2428
rect 11440 2360 11468 2400
rect 13170 2388 13176 2440
rect 13228 2388 13234 2440
rect 10428 2332 11468 2360
rect 11968 2363 12026 2369
rect 11968 2329 11980 2363
rect 12014 2360 12026 2363
rect 13817 2363 13875 2369
rect 13817 2360 13829 2363
rect 12014 2332 13829 2360
rect 12014 2329 12026 2332
rect 11968 2323 12026 2329
rect 13817 2329 13829 2332
rect 13863 2329 13875 2363
rect 13924 2360 13952 2468
rect 14108 2437 14136 2536
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14752 2360 14780 2391
rect 13924 2332 14780 2360
rect 13817 2323 13875 2329
rect 13170 2292 13176 2304
rect 9048 2264 13176 2292
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 14844 2292 14872 2391
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15381 2431 15439 2437
rect 15381 2428 15393 2431
rect 14976 2400 15393 2428
rect 14976 2388 14982 2400
rect 15381 2397 15393 2400
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2397 15991 2431
rect 16040 2428 16068 2536
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 19061 2567 19119 2573
rect 19061 2564 19073 2567
rect 17920 2536 19073 2564
rect 17920 2524 17926 2536
rect 19061 2533 19073 2536
rect 19107 2533 19119 2567
rect 21542 2564 21548 2576
rect 19061 2527 19119 2533
rect 19812 2536 21548 2564
rect 16666 2456 16672 2508
rect 16724 2456 16730 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 18012 2468 19717 2496
rect 18012 2456 18018 2468
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 16758 2428 16764 2440
rect 16040 2400 16764 2428
rect 15933 2391 15991 2397
rect 15948 2360 15976 2391
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16936 2431 16994 2437
rect 16936 2397 16948 2431
rect 16982 2428 16994 2431
rect 17678 2428 17684 2440
rect 16982 2400 17684 2428
rect 16982 2397 16994 2400
rect 16936 2391 16994 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17828 2400 18337 2428
rect 17828 2388 17834 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2430 19487 2431
rect 19518 2430 19524 2440
rect 19475 2402 19524 2430
rect 19475 2397 19487 2402
rect 19429 2391 19487 2397
rect 18230 2360 18236 2372
rect 15948 2332 18236 2360
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 18432 2360 18460 2391
rect 19518 2388 19524 2402
rect 19576 2388 19582 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2424 19671 2431
rect 19812 2430 19840 2536
rect 21542 2524 21548 2536
rect 21600 2564 21606 2576
rect 21600 2536 22094 2564
rect 21600 2524 21606 2536
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2496 20039 2499
rect 20346 2496 20352 2508
rect 20027 2468 20352 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 20622 2456 20628 2508
rect 20680 2456 20686 2508
rect 21082 2456 21088 2508
rect 21140 2456 21146 2508
rect 19720 2424 19840 2430
rect 19659 2402 19840 2424
rect 19659 2397 19748 2402
rect 19613 2396 19748 2397
rect 19613 2391 19671 2396
rect 19812 2360 19840 2402
rect 20806 2388 20812 2440
rect 20864 2388 20870 2440
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 21560 2428 21588 2524
rect 21910 2456 21916 2508
rect 21968 2456 21974 2508
rect 22066 2496 22094 2536
rect 23566 2524 23572 2576
rect 23624 2564 23630 2576
rect 24688 2564 24716 2604
rect 23624 2536 24716 2564
rect 23624 2524 23630 2536
rect 24762 2524 24768 2576
rect 24820 2524 24826 2576
rect 22066 2468 22784 2496
rect 21499 2400 21588 2428
rect 22756 2428 22784 2468
rect 22830 2456 22836 2508
rect 22888 2456 22894 2508
rect 23106 2456 23112 2508
rect 23164 2496 23170 2508
rect 23164 2468 25084 2496
rect 23164 2456 23170 2468
rect 23017 2431 23075 2437
rect 23017 2428 23029 2431
rect 22756 2400 23029 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 23017 2397 23029 2400
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 23750 2388 23756 2440
rect 23808 2388 23814 2440
rect 23842 2388 23848 2440
rect 23900 2388 23906 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 24946 2430 24952 2440
rect 24872 2428 24952 2430
rect 24443 2402 24952 2428
rect 24443 2400 24900 2402
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 24946 2388 24952 2402
rect 25004 2388 25010 2440
rect 18432 2332 19334 2360
rect 13688 2264 14872 2292
rect 13688 2252 13694 2264
rect 15470 2252 15476 2304
rect 15528 2252 15534 2304
rect 18049 2295 18107 2301
rect 18049 2261 18061 2295
rect 18095 2292 18107 2295
rect 18432 2292 18460 2332
rect 18095 2264 18460 2292
rect 19306 2292 19334 2332
rect 19619 2332 19840 2360
rect 20073 2363 20131 2369
rect 19619 2292 19647 2332
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 20119 2332 21404 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 19306 2264 19647 2292
rect 21376 2292 21404 2332
rect 21542 2320 21548 2372
rect 21600 2360 21606 2372
rect 22005 2363 22063 2369
rect 22005 2360 22017 2363
rect 21600 2332 22017 2360
rect 21600 2320 21606 2332
rect 22005 2329 22017 2332
rect 22051 2329 22063 2363
rect 22005 2323 22063 2329
rect 23382 2320 23388 2372
rect 23440 2360 23446 2372
rect 24762 2360 24768 2372
rect 23440 2332 24768 2360
rect 23440 2320 23446 2332
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 25056 2360 25084 2468
rect 25148 2437 25176 2604
rect 25501 2601 25513 2635
rect 25547 2632 25559 2635
rect 25590 2632 25596 2644
rect 25547 2604 25596 2632
rect 25547 2601 25559 2604
rect 25501 2595 25559 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25961 2635 26019 2641
rect 25961 2601 25973 2635
rect 26007 2632 26019 2635
rect 26050 2632 26056 2644
rect 26007 2604 26056 2632
rect 26007 2601 26019 2604
rect 25961 2595 26019 2601
rect 26050 2592 26056 2604
rect 26108 2592 26114 2644
rect 26694 2592 26700 2644
rect 26752 2592 26758 2644
rect 26789 2635 26847 2641
rect 26789 2601 26801 2635
rect 26835 2632 26847 2635
rect 27246 2632 27252 2644
rect 26835 2604 27252 2632
rect 26835 2601 26847 2604
rect 26789 2595 26847 2601
rect 27246 2592 27252 2604
rect 27304 2592 27310 2644
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 28040 2604 28549 2632
rect 28040 2592 28046 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 28537 2595 28595 2601
rect 26712 2564 26740 2592
rect 27617 2567 27675 2573
rect 27617 2564 27629 2567
rect 26712 2536 27629 2564
rect 27617 2533 27629 2536
rect 27663 2533 27675 2567
rect 27617 2527 27675 2533
rect 25682 2456 25688 2508
rect 25740 2496 25746 2508
rect 26145 2499 26203 2505
rect 26145 2496 26157 2499
rect 25740 2468 26157 2496
rect 25740 2456 25746 2468
rect 26145 2465 26157 2468
rect 26191 2465 26203 2499
rect 26145 2459 26203 2465
rect 27062 2456 27068 2508
rect 27120 2456 27126 2508
rect 27985 2499 28043 2505
rect 27985 2465 27997 2499
rect 28031 2496 28043 2499
rect 28534 2496 28540 2508
rect 28031 2468 28540 2496
rect 28031 2465 28043 2468
rect 27985 2459 28043 2465
rect 28534 2456 28540 2468
rect 28592 2456 28598 2508
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2428 25927 2431
rect 28350 2428 28356 2440
rect 25915 2400 28356 2428
rect 25915 2397 25927 2400
rect 25869 2391 25927 2397
rect 25424 2360 25452 2391
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 25056 2332 25452 2360
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 21376 2264 23121 2292
rect 18095 2261 18107 2264
rect 18049 2255 18107 2261
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23474 2252 23480 2304
rect 23532 2252 23538 2304
rect 23566 2252 23572 2304
rect 23624 2252 23630 2304
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 25225 2295 25283 2301
rect 25225 2292 25237 2295
rect 23716 2264 25237 2292
rect 23716 2252 23722 2264
rect 25225 2261 25237 2264
rect 25271 2261 25283 2295
rect 25225 2255 25283 2261
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 2038 2048 2044 2100
rect 2096 2048 2102 2100
rect 2130 2048 2136 2100
rect 2188 2088 2194 2100
rect 23382 2088 23388 2100
rect 2188 2060 23388 2088
rect 2188 2048 2194 2060
rect 23382 2048 23388 2060
rect 23440 2048 23446 2100
rect 23474 2048 23480 2100
rect 23532 2048 23538 2100
rect 23566 2048 23572 2100
rect 23624 2048 23630 2100
rect 2056 2020 2084 2048
rect 2056 1992 2774 2020
rect 2746 1884 2774 1992
rect 4798 1980 4804 2032
rect 4856 2020 4862 2032
rect 10410 2020 10416 2032
rect 4856 1992 10416 2020
rect 4856 1980 4862 1992
rect 10410 1980 10416 1992
rect 10468 1980 10474 2032
rect 11330 1980 11336 2032
rect 11388 1980 11394 2032
rect 11606 1980 11612 2032
rect 11664 2020 11670 2032
rect 13630 2020 13636 2032
rect 11664 1992 13636 2020
rect 11664 1980 11670 1992
rect 13630 1980 13636 1992
rect 13688 1980 13694 2032
rect 15470 1980 15476 2032
rect 15528 1980 15534 2032
rect 19794 1980 19800 2032
rect 19852 2020 19858 2032
rect 23492 2020 23520 2048
rect 19852 1992 23520 2020
rect 19852 1980 19858 1992
rect 11348 1952 11376 1980
rect 15488 1952 15516 1980
rect 11348 1924 15516 1952
rect 17494 1912 17500 1964
rect 17552 1952 17558 1964
rect 21542 1952 21548 1964
rect 17552 1924 21548 1952
rect 17552 1912 17558 1924
rect 21542 1912 21548 1924
rect 21600 1912 21606 1964
rect 23198 1952 23204 1964
rect 21744 1924 23204 1952
rect 2746 1856 15700 1884
rect 9858 1776 9864 1828
rect 9916 1816 9922 1828
rect 13078 1816 13084 1828
rect 9916 1788 13084 1816
rect 9916 1776 9922 1788
rect 13078 1776 13084 1788
rect 13136 1776 13142 1828
rect 15672 1680 15700 1856
rect 16758 1776 16764 1828
rect 16816 1816 16822 1828
rect 21744 1816 21772 1924
rect 23198 1912 23204 1924
rect 23256 1912 23262 1964
rect 16816 1788 21772 1816
rect 16816 1776 16822 1788
rect 18782 1708 18788 1760
rect 18840 1748 18846 1760
rect 23584 1748 23612 2048
rect 18840 1720 23612 1748
rect 18840 1708 18846 1720
rect 24210 1680 24216 1692
rect 15672 1652 24216 1680
rect 24210 1640 24216 1652
rect 24268 1640 24274 1692
<< via1 >>
rect 9680 27820 9732 27872
rect 11980 27820 12032 27872
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 23664 27659 23716 27668
rect 23664 27625 23673 27659
rect 23673 27625 23707 27659
rect 23707 27625 23716 27659
rect 23664 27616 23716 27625
rect 3792 27548 3844 27600
rect 5356 27480 5408 27532
rect 8484 27548 8536 27600
rect 9680 27548 9732 27600
rect 1492 27387 1544 27396
rect 1492 27353 1501 27387
rect 1501 27353 1535 27387
rect 1535 27353 1544 27387
rect 1492 27344 1544 27353
rect 5080 27412 5132 27464
rect 940 27276 992 27328
rect 4620 27319 4672 27328
rect 4620 27285 4629 27319
rect 4629 27285 4663 27319
rect 4663 27285 4672 27319
rect 4620 27276 4672 27285
rect 4804 27276 4856 27328
rect 4896 27319 4948 27328
rect 4896 27285 4905 27319
rect 4905 27285 4939 27319
rect 4939 27285 4948 27319
rect 4896 27276 4948 27285
rect 5448 27319 5500 27328
rect 5448 27285 5457 27319
rect 5457 27285 5491 27319
rect 5491 27285 5500 27319
rect 5448 27276 5500 27285
rect 5724 27319 5776 27328
rect 5724 27285 5733 27319
rect 5733 27285 5767 27319
rect 5767 27285 5776 27319
rect 5724 27276 5776 27285
rect 6000 27276 6052 27328
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 8944 27480 8996 27532
rect 11428 27480 11480 27532
rect 6276 27344 6328 27396
rect 10140 27412 10192 27464
rect 10416 27412 10468 27464
rect 11152 27412 11204 27464
rect 15384 27548 15436 27600
rect 15752 27548 15804 27600
rect 19156 27548 19208 27600
rect 21364 27548 21416 27600
rect 11980 27455 12032 27464
rect 11980 27421 11989 27455
rect 11989 27421 12023 27455
rect 12023 27421 12032 27455
rect 11980 27412 12032 27421
rect 16856 27523 16908 27532
rect 16856 27489 16865 27523
rect 16865 27489 16899 27523
rect 16899 27489 16908 27523
rect 16856 27480 16908 27489
rect 6644 27276 6696 27328
rect 6828 27319 6880 27328
rect 6828 27285 6837 27319
rect 6837 27285 6871 27319
rect 6871 27285 6880 27319
rect 6828 27276 6880 27285
rect 6920 27276 6972 27328
rect 8300 27276 8352 27328
rect 8392 27319 8444 27328
rect 8392 27285 8401 27319
rect 8401 27285 8435 27319
rect 8435 27285 8444 27319
rect 8392 27276 8444 27285
rect 8576 27276 8628 27328
rect 9036 27276 9088 27328
rect 9588 27276 9640 27328
rect 9772 27319 9824 27328
rect 9772 27285 9781 27319
rect 9781 27285 9815 27319
rect 9815 27285 9824 27319
rect 9772 27276 9824 27285
rect 10508 27276 10560 27328
rect 10968 27319 11020 27328
rect 10968 27285 10977 27319
rect 10977 27285 11011 27319
rect 11011 27285 11020 27319
rect 10968 27276 11020 27285
rect 11060 27319 11112 27328
rect 11060 27285 11069 27319
rect 11069 27285 11103 27319
rect 11103 27285 11112 27319
rect 11060 27276 11112 27285
rect 13912 27412 13964 27464
rect 12900 27344 12952 27396
rect 14648 27412 14700 27464
rect 15844 27412 15896 27464
rect 18696 27480 18748 27532
rect 18328 27455 18380 27464
rect 18328 27421 18337 27455
rect 18337 27421 18371 27455
rect 18371 27421 18380 27455
rect 18328 27412 18380 27421
rect 19524 27455 19576 27464
rect 26240 27548 26292 27600
rect 26608 27548 26660 27600
rect 19524 27421 19557 27455
rect 19557 27421 19576 27455
rect 19524 27412 19576 27421
rect 16488 27344 16540 27396
rect 21088 27455 21140 27464
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 22836 27412 22888 27464
rect 24124 27412 24176 27464
rect 25044 27412 25096 27464
rect 26056 27455 26108 27464
rect 26056 27421 26065 27455
rect 26065 27421 26099 27455
rect 26099 27421 26108 27455
rect 26056 27412 26108 27421
rect 28172 27412 28224 27464
rect 24032 27344 24084 27396
rect 27804 27344 27856 27396
rect 12992 27319 13044 27328
rect 12992 27285 13001 27319
rect 13001 27285 13035 27319
rect 13035 27285 13044 27319
rect 12992 27276 13044 27285
rect 13728 27319 13780 27328
rect 13728 27285 13737 27319
rect 13737 27285 13771 27319
rect 13771 27285 13780 27319
rect 13728 27276 13780 27285
rect 14740 27276 14792 27328
rect 15200 27276 15252 27328
rect 16304 27319 16356 27328
rect 16304 27285 16313 27319
rect 16313 27285 16347 27319
rect 16347 27285 16356 27319
rect 16304 27276 16356 27285
rect 17408 27319 17460 27328
rect 17408 27285 17417 27319
rect 17417 27285 17451 27319
rect 17451 27285 17460 27319
rect 17408 27276 17460 27285
rect 17684 27276 17736 27328
rect 18880 27319 18932 27328
rect 18880 27285 18889 27319
rect 18889 27285 18923 27319
rect 18923 27285 18932 27319
rect 18880 27276 18932 27285
rect 19340 27319 19392 27328
rect 19340 27285 19349 27319
rect 19349 27285 19383 27319
rect 19383 27285 19392 27319
rect 19340 27276 19392 27285
rect 19616 27319 19668 27328
rect 19616 27285 19625 27319
rect 19625 27285 19659 27319
rect 19659 27285 19668 27319
rect 19616 27276 19668 27285
rect 20812 27319 20864 27328
rect 20812 27285 20821 27319
rect 20821 27285 20855 27319
rect 20855 27285 20864 27319
rect 20812 27276 20864 27285
rect 21272 27276 21324 27328
rect 22744 27276 22796 27328
rect 26516 27276 26568 27328
rect 28448 27319 28500 27328
rect 28448 27285 28457 27319
rect 28457 27285 28491 27319
rect 28491 27285 28500 27319
rect 28448 27276 28500 27285
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 1492 27072 1544 27124
rect 2596 27047 2648 27056
rect 2596 27013 2605 27047
rect 2605 27013 2639 27047
rect 2639 27013 2648 27047
rect 2596 27004 2648 27013
rect 2688 27047 2740 27056
rect 2688 27013 2697 27047
rect 2697 27013 2731 27047
rect 2731 27013 2740 27047
rect 2688 27004 2740 27013
rect 4620 27072 4672 27124
rect 4896 27072 4948 27124
rect 5448 27072 5500 27124
rect 5724 27072 5776 27124
rect 6736 27072 6788 27124
rect 8300 27072 8352 27124
rect 8392 27072 8444 27124
rect 2320 26936 2372 26988
rect 2228 26775 2280 26784
rect 2228 26741 2237 26775
rect 2237 26741 2271 26775
rect 2271 26741 2280 26775
rect 2228 26732 2280 26741
rect 3792 26936 3844 26988
rect 6644 27004 6696 27056
rect 7012 27004 7064 27056
rect 6000 26979 6052 26988
rect 6000 26945 6009 26979
rect 6009 26945 6043 26979
rect 6043 26945 6052 26979
rect 6000 26936 6052 26945
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 9036 27004 9088 27056
rect 3516 26911 3568 26920
rect 3516 26877 3525 26911
rect 3525 26877 3559 26911
rect 3559 26877 3568 26911
rect 3516 26868 3568 26877
rect 5264 26843 5316 26852
rect 5264 26809 5273 26843
rect 5273 26809 5307 26843
rect 5307 26809 5316 26843
rect 5264 26800 5316 26809
rect 6276 26868 6328 26920
rect 6368 26911 6420 26920
rect 6368 26877 6377 26911
rect 6377 26877 6411 26911
rect 6411 26877 6420 26911
rect 6368 26868 6420 26877
rect 9864 26979 9916 26988
rect 9864 26945 9873 26979
rect 9873 26945 9907 26979
rect 9907 26945 9916 26979
rect 9864 26936 9916 26945
rect 10968 27072 11020 27124
rect 11060 27072 11112 27124
rect 5908 26800 5960 26852
rect 3240 26732 3292 26784
rect 6184 26732 6236 26784
rect 6920 26732 6972 26784
rect 8208 26800 8260 26852
rect 12900 27115 12952 27124
rect 12900 27081 12909 27115
rect 12909 27081 12943 27115
rect 12943 27081 12952 27115
rect 12900 27072 12952 27081
rect 12992 27072 13044 27124
rect 13728 27072 13780 27124
rect 14648 27115 14700 27124
rect 14648 27081 14657 27115
rect 14657 27081 14691 27115
rect 14691 27081 14700 27115
rect 14648 27072 14700 27081
rect 16856 27072 16908 27124
rect 18328 27072 18380 27124
rect 18880 27072 18932 27124
rect 19524 27115 19576 27124
rect 19524 27081 19533 27115
rect 19533 27081 19567 27115
rect 19567 27081 19576 27115
rect 19524 27072 19576 27081
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 9864 26800 9916 26852
rect 10048 26800 10100 26852
rect 10784 26800 10836 26852
rect 12440 26843 12492 26852
rect 12440 26809 12449 26843
rect 12449 26809 12483 26843
rect 12483 26809 12492 26843
rect 12440 26800 12492 26809
rect 14280 26936 14332 26988
rect 13268 26911 13320 26920
rect 13268 26877 13277 26911
rect 13277 26877 13311 26911
rect 13311 26877 13320 26911
rect 13268 26868 13320 26877
rect 16304 26936 16356 26988
rect 17408 26936 17460 26988
rect 21364 27072 21416 27124
rect 22376 27072 22428 27124
rect 22744 27072 22796 27124
rect 26056 27072 26108 27124
rect 20812 27004 20864 27056
rect 15108 26800 15160 26852
rect 17776 26868 17828 26920
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 8392 26775 8444 26784
rect 8392 26741 8401 26775
rect 8401 26741 8435 26775
rect 8435 26741 8444 26775
rect 8392 26732 8444 26741
rect 9404 26775 9456 26784
rect 9404 26741 9413 26775
rect 9413 26741 9447 26775
rect 9447 26741 9456 26775
rect 9404 26732 9456 26741
rect 9680 26775 9732 26784
rect 9680 26741 9689 26775
rect 9689 26741 9723 26775
rect 9723 26741 9732 26775
rect 9680 26732 9732 26741
rect 10140 26732 10192 26784
rect 13176 26732 13228 26784
rect 15292 26732 15344 26784
rect 16580 26732 16632 26784
rect 19248 26732 19300 26784
rect 20628 26732 20680 26784
rect 21548 26775 21600 26784
rect 21548 26741 21557 26775
rect 21557 26741 21591 26775
rect 21591 26741 21600 26775
rect 21548 26732 21600 26741
rect 22744 26868 22796 26920
rect 27252 27004 27304 27056
rect 24216 26936 24268 26988
rect 25780 26936 25832 26988
rect 26516 26936 26568 26988
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 28264 26936 28316 26988
rect 24032 26868 24084 26920
rect 24860 26911 24912 26920
rect 24860 26877 24869 26911
rect 24869 26877 24903 26911
rect 24903 26877 24912 26911
rect 24860 26868 24912 26877
rect 25688 26868 25740 26920
rect 26148 26911 26200 26920
rect 26148 26877 26157 26911
rect 26157 26877 26191 26911
rect 26191 26877 26200 26911
rect 26148 26868 26200 26877
rect 26424 26868 26476 26920
rect 27620 26868 27672 26920
rect 24308 26775 24360 26784
rect 24308 26741 24317 26775
rect 24317 26741 24351 26775
rect 24351 26741 24360 26775
rect 24308 26732 24360 26741
rect 26332 26732 26384 26784
rect 26700 26732 26752 26784
rect 27712 26775 27764 26784
rect 27712 26741 27721 26775
rect 27721 26741 27755 26775
rect 27755 26741 27764 26775
rect 27712 26732 27764 26741
rect 28356 26775 28408 26784
rect 28356 26741 28365 26775
rect 28365 26741 28399 26775
rect 28399 26741 28408 26775
rect 28356 26732 28408 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 2228 26528 2280 26580
rect 2688 26528 2740 26580
rect 3516 26528 3568 26580
rect 5080 26528 5132 26580
rect 6828 26528 6880 26580
rect 8392 26528 8444 26580
rect 8484 26528 8536 26580
rect 9404 26571 9456 26580
rect 9404 26537 9413 26571
rect 9413 26537 9447 26571
rect 9447 26537 9456 26571
rect 9404 26528 9456 26537
rect 9772 26528 9824 26580
rect 12716 26528 12768 26580
rect 13176 26528 13228 26580
rect 5264 26392 5316 26444
rect 6184 26435 6236 26444
rect 6184 26401 6193 26435
rect 6193 26401 6227 26435
rect 6227 26401 6236 26435
rect 6184 26392 6236 26401
rect 4804 26367 4856 26376
rect 4804 26333 4813 26367
rect 4813 26333 4847 26367
rect 4847 26333 4856 26367
rect 6736 26460 6788 26512
rect 6920 26435 6972 26444
rect 6920 26401 6929 26435
rect 6929 26401 6963 26435
rect 6963 26401 6972 26435
rect 6920 26392 6972 26401
rect 7012 26392 7064 26444
rect 12440 26460 12492 26512
rect 13912 26571 13964 26580
rect 13912 26537 13921 26571
rect 13921 26537 13955 26571
rect 13955 26537 13964 26571
rect 13912 26528 13964 26537
rect 15844 26571 15896 26580
rect 15844 26537 15853 26571
rect 15853 26537 15887 26571
rect 15887 26537 15896 26571
rect 15844 26528 15896 26537
rect 15476 26460 15528 26512
rect 4804 26324 4856 26333
rect 7288 26324 7340 26376
rect 7656 26324 7708 26376
rect 7932 26324 7984 26376
rect 8208 26324 8260 26376
rect 8300 26324 8352 26376
rect 8852 26324 8904 26376
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 12348 26392 12400 26444
rect 8944 26324 8996 26333
rect 3240 26188 3292 26240
rect 4344 26231 4396 26240
rect 4344 26197 4353 26231
rect 4353 26197 4387 26231
rect 4387 26197 4396 26231
rect 4344 26188 4396 26197
rect 4896 26188 4948 26240
rect 5172 26188 5224 26240
rect 9588 26256 9640 26308
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 13268 26324 13320 26376
rect 16488 26392 16540 26444
rect 17500 26503 17552 26512
rect 17500 26469 17509 26503
rect 17509 26469 17543 26503
rect 17543 26469 17552 26503
rect 17500 26460 17552 26469
rect 18880 26528 18932 26580
rect 19248 26528 19300 26580
rect 19340 26528 19392 26580
rect 19616 26528 19668 26580
rect 21088 26528 21140 26580
rect 21272 26571 21324 26580
rect 21272 26537 21281 26571
rect 21281 26537 21315 26571
rect 21315 26537 21324 26571
rect 21272 26528 21324 26537
rect 21364 26528 21416 26580
rect 21548 26528 21600 26580
rect 23664 26528 23716 26580
rect 24860 26528 24912 26580
rect 17684 26392 17736 26444
rect 11704 26299 11756 26308
rect 11704 26265 11713 26299
rect 11713 26265 11747 26299
rect 11747 26265 11756 26299
rect 11704 26256 11756 26265
rect 12624 26256 12676 26308
rect 15200 26324 15252 26376
rect 16672 26324 16724 26376
rect 17040 26324 17092 26376
rect 14648 26256 14700 26308
rect 17592 26256 17644 26308
rect 8392 26188 8444 26240
rect 8576 26231 8628 26240
rect 8576 26197 8585 26231
rect 8585 26197 8619 26231
rect 8619 26197 8628 26231
rect 8576 26188 8628 26197
rect 10416 26231 10468 26240
rect 10416 26197 10425 26231
rect 10425 26197 10459 26231
rect 10459 26197 10468 26231
rect 10416 26188 10468 26197
rect 11152 26231 11204 26240
rect 11152 26197 11161 26231
rect 11161 26197 11195 26231
rect 11195 26197 11204 26231
rect 11152 26188 11204 26197
rect 14188 26188 14240 26240
rect 16948 26188 17000 26240
rect 19156 26324 19208 26376
rect 20168 26367 20220 26376
rect 20168 26333 20177 26367
rect 20177 26333 20211 26367
rect 20211 26333 20220 26367
rect 20168 26324 20220 26333
rect 22836 26392 22888 26444
rect 21272 26324 21324 26376
rect 23388 26324 23440 26376
rect 24952 26460 25004 26512
rect 25044 26392 25096 26444
rect 26976 26528 27028 26580
rect 27620 26528 27672 26580
rect 27712 26528 27764 26580
rect 27804 26528 27856 26580
rect 26148 26392 26200 26444
rect 26424 26392 26476 26444
rect 25136 26324 25188 26376
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 25780 26324 25832 26376
rect 18512 26299 18564 26308
rect 18512 26265 18521 26299
rect 18521 26265 18555 26299
rect 18555 26265 18564 26299
rect 18512 26256 18564 26265
rect 26700 26392 26752 26444
rect 28080 26460 28132 26512
rect 27068 26324 27120 26376
rect 28540 26367 28592 26376
rect 28540 26333 28549 26367
rect 28549 26333 28583 26367
rect 28583 26333 28592 26367
rect 28540 26324 28592 26333
rect 18880 26188 18932 26240
rect 27712 26256 27764 26308
rect 22284 26231 22336 26240
rect 22284 26197 22293 26231
rect 22293 26197 22327 26231
rect 22327 26197 22336 26231
rect 22284 26188 22336 26197
rect 23572 26231 23624 26240
rect 23572 26197 23581 26231
rect 23581 26197 23615 26231
rect 23615 26197 23624 26231
rect 23572 26188 23624 26197
rect 25136 26188 25188 26240
rect 25780 26188 25832 26240
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 26240 26188 26292 26240
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 2320 25984 2372 26036
rect 5908 25984 5960 26036
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 1400 25687 1452 25696
rect 1400 25653 1409 25687
rect 1409 25653 1443 25687
rect 1443 25653 1452 25687
rect 1400 25644 1452 25653
rect 2044 25687 2096 25696
rect 2044 25653 2053 25687
rect 2053 25653 2087 25687
rect 2087 25653 2096 25687
rect 2044 25644 2096 25653
rect 2504 25780 2556 25832
rect 3424 25823 3476 25832
rect 3424 25789 3433 25823
rect 3433 25789 3467 25823
rect 3467 25789 3476 25823
rect 3424 25780 3476 25789
rect 3608 25823 3660 25832
rect 3608 25789 3617 25823
rect 3617 25789 3651 25823
rect 3651 25789 3660 25823
rect 3608 25780 3660 25789
rect 3976 25712 4028 25764
rect 6368 25984 6420 26036
rect 7288 25984 7340 26036
rect 10416 26027 10468 26036
rect 10416 25993 10425 26027
rect 10425 25993 10459 26027
rect 10459 25993 10468 26027
rect 10416 25984 10468 25993
rect 12624 25984 12676 26036
rect 14372 25984 14424 26036
rect 14556 25984 14608 26036
rect 21548 25984 21600 26036
rect 22284 25984 22336 26036
rect 6184 25916 6236 25968
rect 6552 25959 6604 25968
rect 6552 25925 6561 25959
rect 6561 25925 6595 25959
rect 6595 25925 6604 25959
rect 6552 25916 6604 25925
rect 5172 25891 5224 25900
rect 8300 25916 8352 25968
rect 5172 25857 5189 25891
rect 5189 25857 5223 25891
rect 5223 25857 5224 25891
rect 5172 25848 5224 25857
rect 6460 25780 6512 25832
rect 8576 25848 8628 25900
rect 9588 25848 9640 25900
rect 9680 25848 9732 25900
rect 14188 25916 14240 25968
rect 14280 25916 14332 25968
rect 12348 25891 12400 25900
rect 12348 25857 12357 25891
rect 12357 25857 12391 25891
rect 12391 25857 12400 25891
rect 12348 25848 12400 25857
rect 3240 25644 3292 25696
rect 6092 25687 6144 25696
rect 6092 25653 6101 25687
rect 6101 25653 6135 25687
rect 6135 25653 6144 25687
rect 6092 25644 6144 25653
rect 7012 25755 7064 25764
rect 7012 25721 7021 25755
rect 7021 25721 7055 25755
rect 7055 25721 7064 25755
rect 7012 25712 7064 25721
rect 7840 25687 7892 25696
rect 7840 25653 7849 25687
rect 7849 25653 7883 25687
rect 7883 25653 7892 25687
rect 7840 25644 7892 25653
rect 9220 25823 9272 25832
rect 9220 25789 9229 25823
rect 9229 25789 9263 25823
rect 9263 25789 9272 25823
rect 9220 25780 9272 25789
rect 8484 25712 8536 25764
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 12440 25780 12492 25789
rect 12716 25780 12768 25832
rect 12808 25780 12860 25832
rect 15292 25848 15344 25900
rect 15384 25848 15436 25900
rect 17500 25848 17552 25900
rect 18512 25891 18564 25900
rect 18512 25857 18521 25891
rect 18521 25857 18555 25891
rect 18555 25857 18564 25891
rect 18512 25848 18564 25857
rect 20168 25916 20220 25968
rect 21456 25916 21508 25968
rect 24952 25984 25004 26036
rect 25596 25984 25648 26036
rect 26056 25984 26108 26036
rect 14740 25780 14792 25832
rect 15752 25823 15804 25832
rect 15752 25789 15761 25823
rect 15761 25789 15795 25823
rect 15795 25789 15804 25823
rect 15752 25780 15804 25789
rect 17408 25780 17460 25832
rect 17776 25823 17828 25832
rect 17776 25789 17785 25823
rect 17785 25789 17819 25823
rect 17819 25789 17828 25823
rect 17776 25780 17828 25789
rect 18696 25823 18748 25832
rect 18696 25789 18705 25823
rect 18705 25789 18739 25823
rect 18739 25789 18748 25823
rect 18696 25780 18748 25789
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 21916 25848 21968 25900
rect 22836 25848 22888 25900
rect 23572 25848 23624 25900
rect 24400 25891 24452 25900
rect 24400 25857 24409 25891
rect 24409 25857 24443 25891
rect 24443 25857 24452 25891
rect 24400 25848 24452 25857
rect 26332 25891 26384 25900
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 27712 25891 27764 25900
rect 27712 25857 27721 25891
rect 27721 25857 27755 25891
rect 27755 25857 27764 25891
rect 27712 25848 27764 25857
rect 28356 25848 28408 25900
rect 13912 25712 13964 25764
rect 20536 25823 20588 25832
rect 20536 25789 20545 25823
rect 20545 25789 20579 25823
rect 20579 25789 20588 25823
rect 20536 25780 20588 25789
rect 13176 25644 13228 25696
rect 15292 25644 15344 25696
rect 16120 25687 16172 25696
rect 16120 25653 16129 25687
rect 16129 25653 16163 25687
rect 16163 25653 16172 25687
rect 16120 25644 16172 25653
rect 16672 25687 16724 25696
rect 16672 25653 16681 25687
rect 16681 25653 16715 25687
rect 16715 25653 16724 25687
rect 16672 25644 16724 25653
rect 17224 25644 17276 25696
rect 17316 25687 17368 25696
rect 17316 25653 17325 25687
rect 17325 25653 17359 25687
rect 17359 25653 17368 25687
rect 17316 25644 17368 25653
rect 18788 25644 18840 25696
rect 21180 25823 21232 25832
rect 21180 25789 21189 25823
rect 21189 25789 21223 25823
rect 21223 25789 21232 25823
rect 21180 25780 21232 25789
rect 22008 25823 22060 25832
rect 22008 25789 22017 25823
rect 22017 25789 22051 25823
rect 22051 25789 22060 25823
rect 22008 25780 22060 25789
rect 23112 25823 23164 25832
rect 23112 25789 23121 25823
rect 23121 25789 23155 25823
rect 23155 25789 23164 25823
rect 23112 25780 23164 25789
rect 24308 25780 24360 25832
rect 26240 25780 26292 25832
rect 26516 25780 26568 25832
rect 20352 25644 20404 25696
rect 21364 25687 21416 25696
rect 21364 25653 21373 25687
rect 21373 25653 21407 25687
rect 21407 25653 21416 25687
rect 21364 25644 21416 25653
rect 21548 25644 21600 25696
rect 22560 25687 22612 25696
rect 22560 25653 22569 25687
rect 22569 25653 22603 25687
rect 22603 25653 22612 25687
rect 22560 25644 22612 25653
rect 24032 25687 24084 25696
rect 24032 25653 24041 25687
rect 24041 25653 24075 25687
rect 24075 25653 24084 25687
rect 24032 25644 24084 25653
rect 24584 25687 24636 25696
rect 24584 25653 24593 25687
rect 24593 25653 24627 25687
rect 24627 25653 24636 25687
rect 24584 25644 24636 25653
rect 27344 25687 27396 25696
rect 27344 25653 27353 25687
rect 27353 25653 27387 25687
rect 27387 25653 27396 25687
rect 27344 25644 27396 25653
rect 27988 25644 28040 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 1400 25440 1452 25492
rect 2044 25440 2096 25492
rect 3608 25440 3660 25492
rect 3976 25483 4028 25492
rect 3976 25449 3985 25483
rect 3985 25449 4019 25483
rect 4019 25449 4028 25483
rect 3976 25440 4028 25449
rect 6552 25440 6604 25492
rect 7840 25440 7892 25492
rect 9220 25440 9272 25492
rect 11704 25440 11756 25492
rect 13912 25483 13964 25492
rect 13912 25449 13921 25483
rect 13921 25449 13955 25483
rect 13955 25449 13964 25483
rect 13912 25440 13964 25449
rect 15476 25440 15528 25492
rect 16120 25440 16172 25492
rect 17040 25483 17092 25492
rect 17040 25449 17049 25483
rect 17049 25449 17083 25483
rect 17083 25449 17092 25483
rect 17040 25440 17092 25449
rect 17776 25440 17828 25492
rect 2504 25372 2556 25424
rect 1676 25236 1728 25288
rect 2596 25279 2648 25288
rect 2596 25245 2605 25279
rect 2605 25245 2639 25279
rect 2639 25245 2648 25279
rect 2596 25236 2648 25245
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 6460 25415 6512 25424
rect 6460 25381 6469 25415
rect 6469 25381 6503 25415
rect 6503 25381 6512 25415
rect 6460 25372 6512 25381
rect 3884 25304 3936 25356
rect 3056 25168 3108 25220
rect 4344 25236 4396 25288
rect 4804 25236 4856 25288
rect 4896 25236 4948 25288
rect 1952 25100 2004 25152
rect 2044 25100 2096 25152
rect 2780 25100 2832 25152
rect 2964 25143 3016 25152
rect 2964 25109 2973 25143
rect 2973 25109 3007 25143
rect 3007 25109 3016 25143
rect 2964 25100 3016 25109
rect 3240 25143 3292 25152
rect 3240 25109 3249 25143
rect 3249 25109 3283 25143
rect 3283 25109 3292 25143
rect 3240 25100 3292 25109
rect 3332 25100 3384 25152
rect 4252 25143 4304 25152
rect 4252 25109 4261 25143
rect 4261 25109 4295 25143
rect 4295 25109 4304 25143
rect 4252 25100 4304 25109
rect 4528 25143 4580 25152
rect 4528 25109 4537 25143
rect 4537 25109 4571 25143
rect 4571 25109 4580 25143
rect 4528 25100 4580 25109
rect 6736 25279 6788 25288
rect 6736 25245 6745 25279
rect 6745 25245 6779 25279
rect 6779 25245 6788 25279
rect 6736 25236 6788 25245
rect 9956 25372 10008 25424
rect 8392 25304 8444 25356
rect 12532 25347 12584 25356
rect 12532 25313 12541 25347
rect 12541 25313 12575 25347
rect 12575 25313 12584 25347
rect 12532 25304 12584 25313
rect 15384 25347 15436 25356
rect 15384 25313 15393 25347
rect 15393 25313 15427 25347
rect 15427 25313 15436 25347
rect 15384 25304 15436 25313
rect 16488 25372 16540 25424
rect 18696 25483 18748 25492
rect 18696 25449 18705 25483
rect 18705 25449 18739 25483
rect 18739 25449 18748 25483
rect 18696 25440 18748 25449
rect 18788 25440 18840 25492
rect 21180 25483 21232 25492
rect 21180 25449 21189 25483
rect 21189 25449 21223 25483
rect 21223 25449 21232 25483
rect 21180 25440 21232 25449
rect 21364 25440 21416 25492
rect 22560 25440 22612 25492
rect 23112 25483 23164 25492
rect 23112 25449 23121 25483
rect 23121 25449 23155 25483
rect 23155 25449 23164 25483
rect 23112 25440 23164 25449
rect 24032 25440 24084 25492
rect 27344 25440 27396 25492
rect 27896 25440 27948 25492
rect 28540 25440 28592 25492
rect 17316 25304 17368 25356
rect 8300 25279 8352 25288
rect 8300 25245 8309 25279
rect 8309 25245 8343 25279
rect 8343 25245 8352 25279
rect 8300 25236 8352 25245
rect 6092 25168 6144 25220
rect 8852 25168 8904 25220
rect 7196 25100 7248 25152
rect 8300 25100 8352 25152
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 11152 25236 11204 25288
rect 11060 25168 11112 25220
rect 12348 25236 12400 25288
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 15200 25236 15252 25288
rect 16948 25279 17000 25288
rect 16948 25245 16957 25279
rect 16957 25245 16991 25279
rect 16991 25245 17000 25279
rect 16948 25236 17000 25245
rect 17500 25275 17552 25288
rect 17500 25241 17509 25275
rect 17509 25241 17543 25275
rect 17543 25241 17552 25275
rect 17500 25236 17552 25241
rect 17684 25236 17736 25288
rect 17868 25279 17920 25288
rect 17868 25245 17877 25279
rect 17877 25245 17911 25279
rect 17911 25245 17920 25279
rect 17868 25236 17920 25245
rect 21456 25304 21508 25356
rect 21916 25347 21968 25356
rect 21916 25313 21925 25347
rect 21925 25313 21959 25347
rect 21959 25313 21968 25347
rect 21916 25304 21968 25313
rect 19064 25279 19116 25288
rect 19064 25245 19073 25279
rect 19073 25245 19107 25279
rect 19107 25245 19116 25279
rect 19064 25236 19116 25245
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 22008 25236 22060 25288
rect 25872 25347 25924 25356
rect 25872 25313 25881 25347
rect 25881 25313 25915 25347
rect 25915 25313 25924 25347
rect 25872 25304 25924 25313
rect 27988 25415 28040 25424
rect 27988 25381 27997 25415
rect 27997 25381 28031 25415
rect 28031 25381 28040 25415
rect 27988 25372 28040 25381
rect 28172 25304 28224 25356
rect 23112 25236 23164 25288
rect 23388 25279 23440 25288
rect 23388 25245 23397 25279
rect 23397 25245 23431 25279
rect 23431 25245 23440 25279
rect 23388 25236 23440 25245
rect 9588 25143 9640 25152
rect 9588 25109 9597 25143
rect 9597 25109 9631 25143
rect 9631 25109 9640 25143
rect 9588 25100 9640 25109
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 12440 25143 12492 25152
rect 12440 25109 12449 25143
rect 12449 25109 12483 25143
rect 12483 25109 12492 25143
rect 12440 25100 12492 25109
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 15200 25143 15252 25152
rect 15200 25109 15209 25143
rect 15209 25109 15243 25143
rect 15243 25109 15252 25143
rect 15200 25100 15252 25109
rect 16304 25168 16356 25220
rect 15660 25100 15712 25152
rect 16764 25143 16816 25152
rect 16764 25109 16773 25143
rect 16773 25109 16807 25143
rect 16807 25109 16816 25143
rect 16764 25100 16816 25109
rect 17684 25100 17736 25152
rect 19708 25100 19760 25152
rect 22192 25100 22244 25152
rect 24584 25211 24636 25220
rect 24584 25177 24593 25211
rect 24593 25177 24627 25211
rect 24627 25177 24636 25211
rect 24584 25168 24636 25177
rect 24860 25168 24912 25220
rect 25964 25236 26016 25288
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 25596 25143 25648 25152
rect 25596 25109 25605 25143
rect 25605 25109 25639 25143
rect 25639 25109 25648 25143
rect 25596 25100 25648 25109
rect 25780 25100 25832 25152
rect 26240 25100 26292 25152
rect 26792 25279 26844 25288
rect 26792 25245 26801 25279
rect 26801 25245 26835 25279
rect 26835 25245 26844 25279
rect 26792 25236 26844 25245
rect 27528 25279 27580 25288
rect 27528 25245 27537 25279
rect 27537 25245 27571 25279
rect 27571 25245 27580 25279
rect 27528 25236 27580 25245
rect 27160 25168 27212 25220
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 4528 24896 4580 24948
rect 7656 24896 7708 24948
rect 7748 24896 7800 24948
rect 10048 24896 10100 24948
rect 2780 24828 2832 24880
rect 1768 24556 1820 24608
rect 2504 24803 2556 24812
rect 2504 24769 2513 24803
rect 2513 24769 2547 24803
rect 2547 24769 2556 24803
rect 2504 24760 2556 24769
rect 3056 24803 3108 24812
rect 3056 24769 3065 24803
rect 3065 24769 3099 24803
rect 3099 24769 3108 24803
rect 3056 24760 3108 24769
rect 7288 24828 7340 24880
rect 3792 24803 3844 24812
rect 3792 24769 3801 24803
rect 3801 24769 3835 24803
rect 3835 24769 3844 24803
rect 3792 24760 3844 24769
rect 5816 24760 5868 24812
rect 3884 24692 3936 24744
rect 5540 24735 5592 24744
rect 5540 24701 5549 24735
rect 5549 24701 5583 24735
rect 5583 24701 5592 24735
rect 5540 24692 5592 24701
rect 5724 24735 5776 24744
rect 5724 24701 5733 24735
rect 5733 24701 5767 24735
rect 5767 24701 5776 24735
rect 5724 24692 5776 24701
rect 6552 24735 6604 24744
rect 6552 24701 6561 24735
rect 6561 24701 6595 24735
rect 6595 24701 6604 24735
rect 6552 24692 6604 24701
rect 7288 24692 7340 24744
rect 7564 24692 7616 24744
rect 8300 24803 8352 24812
rect 8300 24769 8309 24803
rect 8309 24769 8343 24803
rect 8343 24769 8352 24803
rect 8300 24760 8352 24769
rect 8760 24760 8812 24812
rect 10324 24828 10376 24880
rect 10692 24828 10744 24880
rect 9588 24760 9640 24812
rect 11060 24896 11112 24948
rect 14188 24896 14240 24948
rect 14740 24896 14792 24948
rect 15476 24896 15528 24948
rect 15660 24896 15712 24948
rect 11888 24760 11940 24812
rect 12716 24828 12768 24880
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 11704 24692 11756 24744
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 12256 24692 12308 24744
rect 12532 24692 12584 24744
rect 15200 24760 15252 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 17868 24896 17920 24948
rect 19064 24896 19116 24948
rect 20720 24896 20772 24948
rect 24216 24896 24268 24948
rect 16028 24760 16080 24812
rect 16764 24760 16816 24812
rect 17224 24828 17276 24880
rect 3056 24624 3108 24676
rect 7012 24624 7064 24676
rect 14924 24692 14976 24744
rect 2780 24599 2832 24608
rect 2780 24565 2789 24599
rect 2789 24565 2823 24599
rect 2823 24565 2832 24599
rect 2780 24556 2832 24565
rect 3700 24599 3752 24608
rect 3700 24565 3709 24599
rect 3709 24565 3743 24599
rect 3743 24565 3752 24599
rect 3700 24556 3752 24565
rect 3976 24556 4028 24608
rect 4804 24556 4856 24608
rect 5172 24556 5224 24608
rect 6092 24599 6144 24608
rect 6092 24565 6101 24599
rect 6101 24565 6135 24599
rect 6135 24565 6144 24599
rect 6092 24556 6144 24565
rect 7472 24599 7524 24608
rect 7472 24565 7481 24599
rect 7481 24565 7515 24599
rect 7515 24565 7524 24599
rect 7472 24556 7524 24565
rect 8300 24556 8352 24608
rect 10416 24599 10468 24608
rect 10416 24565 10425 24599
rect 10425 24565 10459 24599
rect 10459 24565 10468 24599
rect 10416 24556 10468 24565
rect 10876 24556 10928 24608
rect 11244 24556 11296 24608
rect 11796 24556 11848 24608
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 17592 24624 17644 24676
rect 21088 24828 21140 24880
rect 20628 24760 20680 24812
rect 22100 24803 22152 24812
rect 22100 24769 22134 24803
rect 22134 24769 22152 24803
rect 24032 24828 24084 24880
rect 26516 24896 26568 24948
rect 26792 24896 26844 24948
rect 28172 24896 28224 24948
rect 22100 24760 22152 24769
rect 19800 24692 19852 24744
rect 21456 24692 21508 24744
rect 13544 24556 13596 24608
rect 15384 24556 15436 24608
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 19524 24599 19576 24608
rect 19524 24565 19533 24599
rect 19533 24565 19567 24599
rect 19567 24565 19576 24599
rect 19524 24556 19576 24565
rect 19616 24556 19668 24608
rect 20076 24556 20128 24608
rect 22468 24556 22520 24608
rect 23112 24556 23164 24608
rect 23480 24556 23532 24608
rect 23572 24556 23624 24608
rect 24860 24760 24912 24812
rect 25136 24760 25188 24812
rect 26056 24760 26108 24812
rect 26516 24760 26568 24812
rect 27160 24828 27212 24880
rect 27068 24803 27120 24812
rect 27068 24769 27077 24803
rect 27077 24769 27111 24803
rect 27111 24769 27120 24803
rect 27068 24760 27120 24769
rect 28356 24760 28408 24812
rect 25688 24735 25740 24744
rect 25688 24701 25697 24735
rect 25697 24701 25731 24735
rect 25731 24701 25740 24735
rect 25688 24692 25740 24701
rect 27160 24692 27212 24744
rect 24676 24667 24728 24676
rect 24676 24633 24685 24667
rect 24685 24633 24719 24667
rect 24719 24633 24728 24667
rect 24676 24624 24728 24633
rect 26240 24624 26292 24676
rect 28264 24624 28316 24676
rect 24584 24556 24636 24608
rect 27988 24599 28040 24608
rect 27988 24565 27997 24599
rect 27997 24565 28031 24599
rect 28031 24565 28040 24599
rect 27988 24556 28040 24565
rect 28172 24599 28224 24608
rect 28172 24565 28181 24599
rect 28181 24565 28215 24599
rect 28215 24565 28224 24599
rect 28172 24556 28224 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 1768 24352 1820 24404
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 2136 24080 2188 24132
rect 2872 24352 2924 24404
rect 5724 24352 5776 24404
rect 5816 24352 5868 24404
rect 6552 24395 6604 24404
rect 6552 24361 6561 24395
rect 6561 24361 6595 24395
rect 6595 24361 6604 24395
rect 6552 24352 6604 24361
rect 6644 24352 6696 24404
rect 3700 24284 3752 24336
rect 2964 24216 3016 24268
rect 3240 24216 3292 24268
rect 4252 24148 4304 24200
rect 4896 24216 4948 24268
rect 7288 24284 7340 24336
rect 6828 24216 6880 24268
rect 5172 24191 5224 24200
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 5172 24148 5224 24157
rect 6920 24148 6972 24200
rect 10692 24352 10744 24404
rect 8852 24284 8904 24336
rect 9220 24284 9272 24336
rect 11520 24352 11572 24404
rect 11888 24352 11940 24404
rect 12164 24352 12216 24404
rect 14004 24352 14056 24404
rect 16948 24352 17000 24404
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 19524 24352 19576 24404
rect 19616 24352 19668 24404
rect 23572 24352 23624 24404
rect 24400 24352 24452 24404
rect 24676 24352 24728 24404
rect 25688 24352 25740 24404
rect 25964 24352 26016 24404
rect 27528 24395 27580 24404
rect 27528 24361 27537 24395
rect 27537 24361 27571 24395
rect 27571 24361 27580 24395
rect 27528 24352 27580 24361
rect 14740 24327 14792 24336
rect 14740 24293 14749 24327
rect 14749 24293 14783 24327
rect 14783 24293 14792 24327
rect 14740 24284 14792 24293
rect 15016 24284 15068 24336
rect 6276 24080 6328 24132
rect 3516 24055 3568 24064
rect 3516 24021 3525 24055
rect 3525 24021 3559 24055
rect 3559 24021 3568 24055
rect 3516 24012 3568 24021
rect 4804 24012 4856 24064
rect 4896 24055 4948 24064
rect 4896 24021 4905 24055
rect 4905 24021 4939 24055
rect 4939 24021 4948 24055
rect 4896 24012 4948 24021
rect 5080 24012 5132 24064
rect 7104 24055 7156 24064
rect 7104 24021 7113 24055
rect 7113 24021 7147 24055
rect 7147 24021 7156 24055
rect 7104 24012 7156 24021
rect 7656 24012 7708 24064
rect 7748 24055 7800 24064
rect 7748 24021 7757 24055
rect 7757 24021 7791 24055
rect 7791 24021 7800 24055
rect 7748 24012 7800 24021
rect 8576 24191 8628 24200
rect 8576 24157 8585 24191
rect 8585 24157 8619 24191
rect 8619 24157 8628 24191
rect 8576 24148 8628 24157
rect 8760 24148 8812 24200
rect 9588 24191 9640 24200
rect 9588 24157 9597 24191
rect 9597 24157 9631 24191
rect 9631 24157 9640 24191
rect 9588 24148 9640 24157
rect 10324 24080 10376 24132
rect 10508 24080 10560 24132
rect 11244 24148 11296 24200
rect 11980 24148 12032 24200
rect 8760 24012 8812 24064
rect 9312 24012 9364 24064
rect 10232 24055 10284 24064
rect 10232 24021 10241 24055
rect 10241 24021 10275 24055
rect 10275 24021 10284 24055
rect 10232 24012 10284 24021
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 11152 24080 11204 24132
rect 12440 24080 12492 24132
rect 13544 24167 13596 24200
rect 13544 24148 13553 24167
rect 13553 24148 13587 24167
rect 13587 24148 13596 24167
rect 13912 24191 13964 24200
rect 13912 24157 13921 24191
rect 13921 24157 13955 24191
rect 13955 24157 13964 24191
rect 13912 24148 13964 24157
rect 14004 24148 14056 24200
rect 14372 24191 14424 24200
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 14464 24080 14516 24132
rect 12900 24012 12952 24064
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 14004 24012 14056 24064
rect 14188 24055 14240 24064
rect 14188 24021 14197 24055
rect 14197 24021 14231 24055
rect 14231 24021 14240 24055
rect 14188 24012 14240 24021
rect 15016 24148 15068 24200
rect 15384 24191 15436 24200
rect 15384 24157 15393 24191
rect 15393 24157 15427 24191
rect 15427 24157 15436 24191
rect 15384 24148 15436 24157
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 16304 24148 16356 24157
rect 15476 24012 15528 24064
rect 15752 24012 15804 24064
rect 23664 24284 23716 24336
rect 20720 24148 20772 24200
rect 20628 24080 20680 24132
rect 20996 24191 21048 24200
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 21364 24080 21416 24132
rect 22284 24216 22336 24268
rect 22468 24191 22520 24200
rect 22468 24157 22477 24191
rect 22477 24157 22511 24191
rect 22511 24157 22520 24191
rect 22468 24148 22520 24157
rect 22376 24080 22428 24132
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23848 24080 23900 24132
rect 24676 24148 24728 24200
rect 24860 24080 24912 24132
rect 25504 24148 25556 24200
rect 25596 24148 25648 24200
rect 26056 24148 26108 24200
rect 17592 24055 17644 24064
rect 17592 24021 17601 24055
rect 17601 24021 17635 24055
rect 17635 24021 17644 24055
rect 17592 24012 17644 24021
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 19616 24055 19668 24064
rect 19616 24021 19625 24055
rect 19625 24021 19659 24055
rect 19659 24021 19668 24055
rect 19616 24012 19668 24021
rect 21456 24055 21508 24064
rect 21456 24021 21465 24055
rect 21465 24021 21499 24055
rect 21499 24021 21508 24055
rect 21456 24012 21508 24021
rect 21548 24012 21600 24064
rect 22192 24012 22244 24064
rect 22560 24055 22612 24064
rect 22560 24021 22569 24055
rect 22569 24021 22603 24055
rect 22603 24021 22612 24055
rect 22560 24012 22612 24021
rect 22836 24055 22888 24064
rect 22836 24021 22845 24055
rect 22845 24021 22879 24055
rect 22879 24021 22888 24055
rect 22836 24012 22888 24021
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 23756 24055 23808 24064
rect 23756 24021 23765 24055
rect 23765 24021 23799 24055
rect 23799 24021 23808 24055
rect 23756 24012 23808 24021
rect 24952 24012 25004 24064
rect 26516 24148 26568 24200
rect 26792 24080 26844 24132
rect 27160 24012 27212 24064
rect 27896 24123 27948 24132
rect 27896 24089 27905 24123
rect 27905 24089 27939 24123
rect 27939 24089 27948 24123
rect 27896 24080 27948 24089
rect 28080 24080 28132 24132
rect 28264 24080 28316 24132
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 2136 23851 2188 23860
rect 2136 23817 2145 23851
rect 2145 23817 2179 23851
rect 2179 23817 2188 23851
rect 2136 23808 2188 23817
rect 3792 23808 3844 23860
rect 3884 23740 3936 23792
rect 2228 23715 2280 23724
rect 2228 23681 2237 23715
rect 2237 23681 2271 23715
rect 2271 23681 2280 23715
rect 2228 23672 2280 23681
rect 3516 23672 3568 23724
rect 4896 23808 4948 23860
rect 6092 23851 6144 23860
rect 6092 23817 6101 23851
rect 6101 23817 6135 23851
rect 6135 23817 6144 23851
rect 6092 23808 6144 23817
rect 6276 23808 6328 23860
rect 6552 23808 6604 23860
rect 7564 23808 7616 23860
rect 7748 23808 7800 23860
rect 8668 23808 8720 23860
rect 4988 23672 5040 23724
rect 3240 23604 3292 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 8208 23740 8260 23792
rect 10232 23808 10284 23860
rect 10324 23808 10376 23860
rect 11704 23808 11756 23860
rect 12808 23808 12860 23860
rect 13360 23808 13412 23860
rect 14096 23808 14148 23860
rect 14188 23808 14240 23860
rect 14740 23808 14792 23860
rect 15384 23808 15436 23860
rect 18236 23808 18288 23860
rect 6000 23604 6052 23656
rect 7196 23672 7248 23724
rect 7656 23672 7708 23724
rect 8668 23672 8720 23724
rect 7380 23647 7432 23656
rect 7380 23613 7389 23647
rect 7389 23613 7423 23647
rect 7423 23613 7432 23647
rect 7380 23604 7432 23613
rect 4344 23536 4396 23588
rect 6920 23536 6972 23588
rect 8208 23604 8260 23656
rect 9864 23604 9916 23656
rect 10416 23604 10468 23656
rect 2596 23468 2648 23520
rect 4252 23468 4304 23520
rect 5172 23511 5224 23520
rect 5172 23477 5181 23511
rect 5181 23477 5215 23511
rect 5215 23477 5224 23511
rect 5172 23468 5224 23477
rect 7196 23511 7248 23520
rect 7196 23477 7205 23511
rect 7205 23477 7239 23511
rect 7239 23477 7248 23511
rect 7196 23468 7248 23477
rect 8576 23536 8628 23588
rect 7748 23511 7800 23520
rect 7748 23477 7757 23511
rect 7757 23477 7791 23511
rect 7791 23477 7800 23511
rect 7748 23468 7800 23477
rect 8668 23511 8720 23520
rect 8668 23477 8677 23511
rect 8677 23477 8711 23511
rect 8711 23477 8720 23511
rect 8668 23468 8720 23477
rect 9220 23536 9272 23588
rect 10968 23579 11020 23588
rect 10968 23545 10977 23579
rect 10977 23545 11011 23579
rect 11011 23545 11020 23579
rect 10968 23536 11020 23545
rect 11244 23536 11296 23588
rect 11520 23536 11572 23588
rect 12256 23604 12308 23656
rect 12072 23536 12124 23588
rect 9496 23468 9548 23520
rect 11704 23468 11756 23520
rect 12808 23468 12860 23520
rect 16028 23715 16080 23724
rect 16028 23681 16037 23715
rect 16037 23681 16071 23715
rect 16071 23681 16080 23715
rect 16028 23672 16080 23681
rect 17592 23672 17644 23724
rect 16304 23604 16356 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 20996 23808 21048 23860
rect 23572 23808 23624 23860
rect 23756 23808 23808 23860
rect 18880 23740 18932 23792
rect 19708 23740 19760 23792
rect 19984 23783 20036 23792
rect 19984 23749 19993 23783
rect 19993 23749 20027 23783
rect 20027 23749 20036 23783
rect 19984 23740 20036 23749
rect 20076 23740 20128 23792
rect 21456 23672 21508 23724
rect 22560 23672 22612 23724
rect 20260 23647 20312 23656
rect 20260 23613 20269 23647
rect 20269 23613 20303 23647
rect 20303 23613 20312 23647
rect 20260 23604 20312 23613
rect 20628 23604 20680 23656
rect 21272 23604 21324 23656
rect 22376 23604 22428 23656
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 23204 23740 23256 23792
rect 25044 23740 25096 23792
rect 26792 23851 26844 23860
rect 26792 23817 26801 23851
rect 26801 23817 26835 23851
rect 26835 23817 26844 23851
rect 26792 23808 26844 23817
rect 27988 23808 28040 23860
rect 28356 23851 28408 23860
rect 28356 23817 28365 23851
rect 28365 23817 28399 23851
rect 28399 23817 28408 23851
rect 28356 23808 28408 23817
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 24584 23672 24636 23724
rect 26056 23672 26108 23724
rect 19340 23536 19392 23588
rect 17040 23511 17092 23520
rect 17040 23477 17049 23511
rect 17049 23477 17083 23511
rect 17083 23477 17092 23511
rect 17040 23468 17092 23477
rect 19984 23468 20036 23520
rect 22192 23511 22244 23520
rect 22192 23477 22201 23511
rect 22201 23477 22235 23511
rect 22235 23477 22244 23511
rect 22192 23468 22244 23477
rect 23388 23468 23440 23520
rect 25136 23604 25188 23656
rect 24676 23536 24728 23588
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 25044 23468 25096 23520
rect 28264 23468 28316 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 2596 23264 2648 23316
rect 2780 23128 2832 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2228 23060 2280 23112
rect 3976 23264 4028 23316
rect 4988 23264 5040 23316
rect 4896 23196 4948 23248
rect 3884 23060 3936 23112
rect 7288 23264 7340 23316
rect 7748 23307 7800 23316
rect 7748 23273 7757 23307
rect 7757 23273 7791 23307
rect 7791 23273 7800 23307
rect 7748 23264 7800 23273
rect 8668 23307 8720 23316
rect 8668 23273 8677 23307
rect 8677 23273 8711 23307
rect 8711 23273 8720 23307
rect 8668 23264 8720 23273
rect 11152 23264 11204 23316
rect 10324 23196 10376 23248
rect 7472 23128 7524 23180
rect 8300 23171 8352 23180
rect 8300 23137 8309 23171
rect 8309 23137 8343 23171
rect 8343 23137 8352 23171
rect 8300 23128 8352 23137
rect 10232 23128 10284 23180
rect 11244 23128 11296 23180
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 12808 23171 12860 23180
rect 12808 23137 12817 23171
rect 12817 23137 12851 23171
rect 12851 23137 12860 23171
rect 12808 23128 12860 23137
rect 14004 23128 14056 23180
rect 3332 22992 3384 23044
rect 4252 22992 4304 23044
rect 5356 23035 5408 23044
rect 5356 23001 5365 23035
rect 5365 23001 5399 23035
rect 5399 23001 5408 23035
rect 5356 22992 5408 23001
rect 4160 22924 4212 22976
rect 6736 22992 6788 23044
rect 7104 22992 7156 23044
rect 7748 22992 7800 23044
rect 8576 23060 8628 23112
rect 9220 23060 9272 23112
rect 9312 23060 9364 23112
rect 9496 23103 9548 23112
rect 9496 23069 9505 23103
rect 9505 23069 9539 23103
rect 9539 23069 9548 23103
rect 9496 23060 9548 23069
rect 9588 23060 9640 23112
rect 9864 23060 9916 23112
rect 11888 23060 11940 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14280 23060 14332 23112
rect 16580 23060 16632 23112
rect 10140 23035 10192 23044
rect 10140 23001 10149 23035
rect 10149 23001 10183 23035
rect 10183 23001 10192 23035
rect 10140 22992 10192 23001
rect 7656 22924 7708 22976
rect 9772 22924 9824 22976
rect 10968 23035 11020 23044
rect 10968 23001 10977 23035
rect 10977 23001 11011 23035
rect 11011 23001 11020 23035
rect 10968 22992 11020 23001
rect 11060 23035 11112 23044
rect 11060 23001 11069 23035
rect 11069 23001 11103 23035
rect 11103 23001 11112 23035
rect 11060 22992 11112 23001
rect 11796 22992 11848 23044
rect 16488 22992 16540 23044
rect 17592 23307 17644 23316
rect 17592 23273 17601 23307
rect 17601 23273 17635 23307
rect 17635 23273 17644 23307
rect 17592 23264 17644 23273
rect 18052 23264 18104 23316
rect 21456 23264 21508 23316
rect 22192 23307 22244 23316
rect 22192 23273 22201 23307
rect 22201 23273 22235 23307
rect 22235 23273 22244 23307
rect 22192 23264 22244 23273
rect 17040 23128 17092 23180
rect 17224 23103 17276 23112
rect 17224 23069 17233 23103
rect 17233 23069 17267 23103
rect 17267 23069 17276 23103
rect 17224 23060 17276 23069
rect 17592 23060 17644 23112
rect 19708 23171 19760 23180
rect 19708 23137 19717 23171
rect 19717 23137 19751 23171
rect 19751 23137 19760 23171
rect 19708 23128 19760 23137
rect 20996 23196 21048 23248
rect 21548 23196 21600 23248
rect 22100 23128 22152 23180
rect 20628 23060 20680 23112
rect 20812 23060 20864 23112
rect 22468 23060 22520 23112
rect 14740 22967 14792 22976
rect 14740 22933 14749 22967
rect 14749 22933 14783 22967
rect 14783 22933 14792 22967
rect 14740 22924 14792 22933
rect 15200 22924 15252 22976
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 18512 22967 18564 22976
rect 18512 22933 18521 22967
rect 18521 22933 18555 22967
rect 18555 22933 18564 22967
rect 18512 22924 18564 22933
rect 18972 22992 19024 23044
rect 19340 23035 19392 23044
rect 19340 23001 19349 23035
rect 19349 23001 19383 23035
rect 19383 23001 19392 23035
rect 19340 22992 19392 23001
rect 19616 22992 19668 23044
rect 20720 22992 20772 23044
rect 21640 22992 21692 23044
rect 19892 22924 19944 22976
rect 20904 22924 20956 22976
rect 21548 22924 21600 22976
rect 23388 23264 23440 23316
rect 23572 23264 23624 23316
rect 23848 23264 23900 23316
rect 26056 23307 26108 23316
rect 26056 23273 26065 23307
rect 26065 23273 26099 23307
rect 26099 23273 26108 23307
rect 26056 23264 26108 23273
rect 23296 23196 23348 23248
rect 22836 23171 22888 23180
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 23480 23128 23532 23180
rect 24676 23171 24728 23180
rect 24676 23137 24685 23171
rect 24685 23137 24719 23171
rect 24719 23137 24728 23171
rect 24676 23128 24728 23137
rect 23572 23103 23624 23112
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23572 23060 23624 23069
rect 23664 23060 23716 23112
rect 24124 23103 24176 23112
rect 24124 23069 24133 23103
rect 24133 23069 24167 23103
rect 24167 23069 24176 23103
rect 24124 23060 24176 23069
rect 24952 23103 25004 23112
rect 24952 23069 24986 23103
rect 24986 23069 25004 23103
rect 23112 22992 23164 23044
rect 24952 23060 25004 23069
rect 27160 23264 27212 23316
rect 26976 23196 27028 23248
rect 28264 23196 28316 23248
rect 27988 23128 28040 23180
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 26792 22967 26844 22976
rect 26792 22933 26801 22967
rect 26801 22933 26835 22967
rect 26835 22933 26844 22967
rect 26792 22924 26844 22933
rect 27160 23060 27212 23112
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 27896 23035 27948 23044
rect 27896 23001 27905 23035
rect 27905 23001 27939 23035
rect 27939 23001 27948 23035
rect 27896 22992 27948 23001
rect 28172 22992 28224 23044
rect 27528 22967 27580 22976
rect 27528 22933 27537 22967
rect 27537 22933 27571 22967
rect 27571 22933 27580 22967
rect 27528 22924 27580 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 3332 22763 3384 22772
rect 3332 22729 3341 22763
rect 3341 22729 3375 22763
rect 3375 22729 3384 22763
rect 3332 22720 3384 22729
rect 4160 22720 4212 22772
rect 5448 22720 5500 22772
rect 6184 22720 6236 22772
rect 6644 22720 6696 22772
rect 7196 22720 7248 22772
rect 7380 22720 7432 22772
rect 3240 22652 3292 22704
rect 2504 22584 2556 22636
rect 2964 22584 3016 22636
rect 3608 22627 3660 22636
rect 3608 22593 3617 22627
rect 3617 22593 3651 22627
rect 3651 22593 3660 22627
rect 3608 22584 3660 22593
rect 4344 22584 4396 22636
rect 5172 22584 5224 22636
rect 6000 22584 6052 22636
rect 6828 22652 6880 22704
rect 11888 22720 11940 22772
rect 14372 22720 14424 22772
rect 14740 22720 14792 22772
rect 15476 22720 15528 22772
rect 17132 22720 17184 22772
rect 17224 22720 17276 22772
rect 18512 22720 18564 22772
rect 6368 22584 6420 22636
rect 2688 22559 2740 22568
rect 2688 22525 2697 22559
rect 2697 22525 2731 22559
rect 2731 22525 2740 22559
rect 2688 22516 2740 22525
rect 2412 22448 2464 22500
rect 4896 22516 4948 22568
rect 4988 22516 5040 22568
rect 5632 22448 5684 22500
rect 2780 22380 2832 22432
rect 5816 22380 5868 22432
rect 5908 22423 5960 22432
rect 5908 22389 5917 22423
rect 5917 22389 5951 22423
rect 5951 22389 5960 22423
rect 5908 22380 5960 22389
rect 7748 22584 7800 22636
rect 8116 22584 8168 22636
rect 8668 22652 8720 22704
rect 9588 22695 9640 22704
rect 9588 22661 9597 22695
rect 9597 22661 9631 22695
rect 9631 22661 9640 22695
rect 9588 22652 9640 22661
rect 10876 22652 10928 22704
rect 11704 22695 11756 22704
rect 11704 22661 11713 22695
rect 11713 22661 11747 22695
rect 11747 22661 11756 22695
rect 11704 22652 11756 22661
rect 14188 22584 14240 22636
rect 8300 22516 8352 22568
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 11060 22448 11112 22500
rect 8116 22380 8168 22432
rect 9128 22380 9180 22432
rect 11244 22380 11296 22432
rect 12256 22516 12308 22568
rect 15200 22516 15252 22568
rect 14464 22448 14516 22500
rect 15752 22559 15804 22568
rect 15752 22525 15761 22559
rect 15761 22525 15795 22559
rect 15795 22525 15804 22559
rect 15752 22516 15804 22525
rect 16028 22627 16080 22636
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 16304 22584 16356 22636
rect 19892 22695 19944 22704
rect 19892 22661 19901 22695
rect 19901 22661 19935 22695
rect 19935 22661 19944 22695
rect 19892 22652 19944 22661
rect 22560 22720 22612 22772
rect 23572 22720 23624 22772
rect 24124 22720 24176 22772
rect 24860 22720 24912 22772
rect 26056 22720 26108 22772
rect 26332 22720 26384 22772
rect 26792 22720 26844 22772
rect 20720 22584 20772 22636
rect 21088 22584 21140 22636
rect 17592 22516 17644 22568
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 18328 22559 18380 22568
rect 18328 22525 18337 22559
rect 18337 22525 18371 22559
rect 18371 22525 18380 22559
rect 18328 22516 18380 22525
rect 17684 22423 17736 22432
rect 17684 22389 17693 22423
rect 17693 22389 17727 22423
rect 17727 22389 17736 22423
rect 17684 22380 17736 22389
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 22008 22584 22060 22636
rect 22284 22627 22336 22636
rect 22284 22593 22293 22627
rect 22293 22593 22327 22627
rect 22327 22593 22336 22627
rect 22284 22584 22336 22593
rect 20444 22448 20496 22500
rect 20536 22448 20588 22500
rect 22376 22516 22428 22568
rect 21916 22491 21968 22500
rect 21916 22457 21925 22491
rect 21925 22457 21959 22491
rect 21959 22457 21968 22491
rect 21916 22448 21968 22457
rect 22008 22448 22060 22500
rect 22468 22448 22520 22500
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 25596 22584 25648 22636
rect 26608 22584 26660 22636
rect 27896 22720 27948 22772
rect 26240 22448 26292 22500
rect 27712 22516 27764 22568
rect 27896 22559 27948 22568
rect 27896 22525 27905 22559
rect 27905 22525 27939 22559
rect 27939 22525 27948 22559
rect 27896 22516 27948 22525
rect 19616 22380 19668 22432
rect 22192 22380 22244 22432
rect 23020 22423 23072 22432
rect 23020 22389 23029 22423
rect 23029 22389 23063 22423
rect 23063 22389 23072 22423
rect 23020 22380 23072 22389
rect 23480 22423 23532 22432
rect 23480 22389 23489 22423
rect 23489 22389 23523 22423
rect 23523 22389 23532 22423
rect 23480 22380 23532 22389
rect 24124 22423 24176 22432
rect 24124 22389 24133 22423
rect 24133 22389 24167 22423
rect 24167 22389 24176 22423
rect 24124 22380 24176 22389
rect 24768 22380 24820 22432
rect 25780 22423 25832 22432
rect 25780 22389 25789 22423
rect 25789 22389 25823 22423
rect 25823 22389 25832 22423
rect 25780 22380 25832 22389
rect 26332 22380 26384 22432
rect 26424 22423 26476 22432
rect 26424 22389 26433 22423
rect 26433 22389 26467 22423
rect 26467 22389 26476 22423
rect 26424 22380 26476 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 2688 22176 2740 22228
rect 3608 22176 3660 22228
rect 5356 22176 5408 22228
rect 2504 22108 2556 22160
rect 3332 22108 3384 22160
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 3700 22040 3752 22092
rect 6000 22108 6052 22160
rect 6184 22176 6236 22228
rect 7472 22176 7524 22228
rect 7564 22176 7616 22228
rect 9588 22176 9640 22228
rect 11704 22219 11756 22228
rect 11704 22185 11713 22219
rect 11713 22185 11747 22219
rect 11747 22185 11756 22219
rect 11704 22176 11756 22185
rect 14096 22176 14148 22228
rect 15108 22176 15160 22228
rect 16304 22176 16356 22228
rect 9864 22108 9916 22160
rect 10140 22108 10192 22160
rect 3148 22015 3200 22024
rect 3148 21981 3157 22015
rect 3157 21981 3191 22015
rect 3191 21981 3200 22015
rect 3148 21972 3200 21981
rect 3424 21972 3476 22024
rect 5264 22083 5316 22092
rect 5264 22049 5273 22083
rect 5273 22049 5307 22083
rect 5307 22049 5316 22083
rect 5264 22040 5316 22049
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 8392 22040 8444 22092
rect 8668 22040 8720 22092
rect 8852 22040 8904 22092
rect 10968 22040 11020 22092
rect 12256 22083 12308 22092
rect 12256 22049 12265 22083
rect 12265 22049 12299 22083
rect 12299 22049 12308 22083
rect 12256 22040 12308 22049
rect 4344 21972 4396 22024
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 2228 21904 2280 21956
rect 5540 21972 5592 22024
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 4068 21836 4120 21888
rect 4620 21879 4672 21888
rect 4620 21845 4629 21879
rect 4629 21845 4663 21879
rect 4663 21845 4672 21879
rect 4620 21836 4672 21845
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 5724 21836 5776 21888
rect 5816 21836 5868 21888
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 7656 22015 7708 22024
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12808 21972 12860 22024
rect 18144 22176 18196 22228
rect 19616 22219 19668 22228
rect 19616 22185 19625 22219
rect 19625 22185 19659 22219
rect 19659 22185 19668 22219
rect 19616 22176 19668 22185
rect 20536 22176 20588 22228
rect 20812 22176 20864 22228
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 16304 21972 16356 22024
rect 20444 22040 20496 22092
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 17684 21972 17736 22024
rect 6552 21836 6604 21888
rect 7748 21879 7800 21888
rect 7748 21845 7757 21879
rect 7757 21845 7791 21879
rect 7791 21845 7800 21879
rect 7748 21836 7800 21845
rect 8484 21836 8536 21888
rect 9680 21904 9732 21956
rect 9956 21947 10008 21956
rect 9956 21913 9965 21947
rect 9965 21913 9999 21947
rect 9999 21913 10008 21947
rect 9956 21904 10008 21913
rect 10140 21947 10192 21956
rect 10140 21913 10149 21947
rect 10149 21913 10183 21947
rect 10183 21913 10192 21947
rect 10140 21904 10192 21913
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 9772 21836 9824 21888
rect 10416 21904 10468 21956
rect 10324 21836 10376 21888
rect 13268 21904 13320 21956
rect 15568 21904 15620 21956
rect 13912 21836 13964 21888
rect 17500 21836 17552 21888
rect 19892 21972 19944 22024
rect 19984 22015 20036 22024
rect 19984 21981 19993 22015
rect 19993 21981 20027 22015
rect 20027 21981 20036 22015
rect 19984 21972 20036 21981
rect 25504 22151 25556 22160
rect 25504 22117 25513 22151
rect 25513 22117 25547 22151
rect 25547 22117 25556 22151
rect 25504 22108 25556 22117
rect 21548 22040 21600 22092
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 18788 21836 18840 21888
rect 20536 21836 20588 21888
rect 20628 21879 20680 21888
rect 20628 21845 20637 21879
rect 20637 21845 20671 21879
rect 20671 21845 20680 21879
rect 20628 21836 20680 21845
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 21364 21972 21416 22024
rect 22284 21972 22336 22024
rect 23296 22083 23348 22092
rect 23296 22049 23305 22083
rect 23305 22049 23339 22083
rect 23339 22049 23348 22083
rect 23296 22040 23348 22049
rect 24768 22040 24820 22092
rect 24952 22040 25004 22092
rect 26424 22040 26476 22092
rect 27528 22083 27580 22092
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 23480 21972 23532 22024
rect 24032 21972 24084 22024
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25320 22015 25372 22024
rect 25320 21981 25329 22015
rect 25329 21981 25363 22015
rect 25363 21981 25372 22015
rect 25320 21972 25372 21981
rect 25504 21904 25556 21956
rect 26792 22015 26844 22024
rect 26792 21981 26801 22015
rect 26801 21981 26835 22015
rect 26835 21981 26844 22015
rect 26792 21972 26844 21981
rect 27436 21972 27488 22024
rect 27896 21904 27948 21956
rect 22192 21836 22244 21888
rect 22652 21836 22704 21888
rect 23388 21836 23440 21888
rect 26240 21836 26292 21888
rect 28080 21879 28132 21888
rect 28080 21845 28089 21879
rect 28089 21845 28123 21879
rect 28123 21845 28132 21879
rect 28080 21836 28132 21845
rect 28356 21879 28408 21888
rect 28356 21845 28365 21879
rect 28365 21845 28399 21879
rect 28399 21845 28408 21879
rect 28356 21836 28408 21845
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 2228 21675 2280 21684
rect 2228 21641 2237 21675
rect 2237 21641 2271 21675
rect 2271 21641 2280 21675
rect 2228 21632 2280 21641
rect 2688 21632 2740 21684
rect 4620 21632 4672 21684
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 5540 21632 5592 21684
rect 7564 21632 7616 21684
rect 8484 21632 8536 21684
rect 9588 21632 9640 21684
rect 9956 21632 10008 21684
rect 11060 21632 11112 21684
rect 14280 21632 14332 21684
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 2044 21496 2096 21548
rect 4712 21564 4764 21616
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 2964 21496 3016 21548
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 4896 21496 4948 21548
rect 4988 21496 5040 21548
rect 5356 21496 5408 21548
rect 3884 21428 3936 21480
rect 5264 21428 5316 21480
rect 5540 21471 5592 21480
rect 5540 21437 5549 21471
rect 5549 21437 5583 21471
rect 5583 21437 5592 21471
rect 5540 21428 5592 21437
rect 7012 21564 7064 21616
rect 7656 21564 7708 21616
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 6828 21496 6880 21548
rect 8944 21564 8996 21616
rect 12900 21564 12952 21616
rect 8208 21471 8260 21480
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 10416 21496 10468 21548
rect 8944 21428 8996 21480
rect 9036 21471 9088 21480
rect 9036 21437 9045 21471
rect 9045 21437 9079 21471
rect 9079 21437 9088 21471
rect 9036 21428 9088 21437
rect 10692 21471 10744 21480
rect 6460 21360 6512 21412
rect 3700 21335 3752 21344
rect 3700 21301 3709 21335
rect 3709 21301 3743 21335
rect 3743 21301 3752 21335
rect 3700 21292 3752 21301
rect 7564 21292 7616 21344
rect 8116 21360 8168 21412
rect 8392 21292 8444 21344
rect 8852 21292 8904 21344
rect 9128 21292 9180 21344
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 12992 21496 13044 21548
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 15016 21496 15068 21548
rect 10600 21360 10652 21412
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 18236 21632 18288 21684
rect 19984 21632 20036 21684
rect 16580 21564 16632 21616
rect 15936 21496 15988 21548
rect 17500 21539 17552 21548
rect 17500 21505 17509 21539
rect 17509 21505 17543 21539
rect 17543 21505 17552 21539
rect 17500 21496 17552 21505
rect 19800 21564 19852 21616
rect 18696 21496 18748 21548
rect 23756 21632 23808 21684
rect 24952 21675 25004 21684
rect 24952 21641 24961 21675
rect 24961 21641 24995 21675
rect 24995 21641 25004 21675
rect 24952 21632 25004 21641
rect 25320 21675 25372 21684
rect 25320 21641 25329 21675
rect 25329 21641 25363 21675
rect 25363 21641 25372 21675
rect 25320 21632 25372 21641
rect 26240 21675 26292 21684
rect 26240 21641 26249 21675
rect 26249 21641 26283 21675
rect 26283 21641 26292 21675
rect 26240 21632 26292 21641
rect 26792 21632 26844 21684
rect 26976 21632 27028 21684
rect 11060 21360 11112 21412
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 16488 21428 16540 21480
rect 20628 21496 20680 21548
rect 20904 21496 20956 21548
rect 21640 21496 21692 21548
rect 22192 21496 22244 21548
rect 23388 21496 23440 21548
rect 24676 21564 24728 21616
rect 24860 21496 24912 21548
rect 20536 21428 20588 21480
rect 21088 21360 21140 21412
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 22928 21428 22980 21480
rect 23204 21428 23256 21480
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 23756 21428 23808 21480
rect 24492 21471 24544 21480
rect 24492 21437 24501 21471
rect 24501 21437 24535 21471
rect 24535 21437 24544 21471
rect 24492 21428 24544 21437
rect 26332 21496 26384 21548
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 9864 21292 9916 21344
rect 13636 21335 13688 21344
rect 13636 21301 13645 21335
rect 13645 21301 13679 21335
rect 13679 21301 13688 21335
rect 13636 21292 13688 21301
rect 14924 21335 14976 21344
rect 14924 21301 14933 21335
rect 14933 21301 14967 21335
rect 14967 21301 14976 21335
rect 14924 21292 14976 21301
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 21456 21292 21508 21344
rect 23940 21292 23992 21344
rect 28632 21292 28684 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 1676 21088 1728 21140
rect 3884 21088 3936 21140
rect 4344 21088 4396 21140
rect 5080 21088 5132 21140
rect 6460 21131 6512 21140
rect 6460 21097 6469 21131
rect 6469 21097 6503 21131
rect 6503 21097 6512 21131
rect 6460 21088 6512 21097
rect 6828 21088 6880 21140
rect 13268 21131 13320 21140
rect 13268 21097 13277 21131
rect 13277 21097 13311 21131
rect 13311 21097 13320 21131
rect 13268 21088 13320 21097
rect 13728 21088 13780 21140
rect 14924 21088 14976 21140
rect 15752 21088 15804 21140
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 16304 21088 16356 21140
rect 20904 21088 20956 21140
rect 22284 21131 22336 21140
rect 22284 21097 22293 21131
rect 22293 21097 22327 21131
rect 22327 21097 22336 21131
rect 22284 21088 22336 21097
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 3424 20927 3476 20936
rect 2596 20816 2648 20868
rect 3424 20893 3433 20927
rect 3433 20893 3467 20927
rect 3467 20893 3476 20927
rect 3424 20884 3476 20893
rect 3700 20884 3752 20936
rect 4068 20884 4120 20936
rect 3332 20816 3384 20868
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5908 20884 5960 20936
rect 9680 21020 9732 21072
rect 10324 21020 10376 21072
rect 10416 21020 10468 21072
rect 10968 20952 11020 21004
rect 8116 20816 8168 20868
rect 8208 20816 8260 20868
rect 9128 20859 9180 20868
rect 9128 20825 9137 20859
rect 9137 20825 9171 20859
rect 9171 20825 9180 20859
rect 9128 20816 9180 20825
rect 10048 20859 10100 20868
rect 10048 20825 10057 20859
rect 10057 20825 10091 20859
rect 10091 20825 10100 20859
rect 10048 20816 10100 20825
rect 10416 20816 10468 20868
rect 10692 20816 10744 20868
rect 18328 21063 18380 21072
rect 18328 21029 18337 21063
rect 18337 21029 18371 21063
rect 18371 21029 18380 21063
rect 18328 21020 18380 21029
rect 23480 21088 23532 21140
rect 23664 21088 23716 21140
rect 24492 21088 24544 21140
rect 11244 20884 11296 20936
rect 12992 20884 13044 20936
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 15292 20884 15344 20936
rect 16488 20927 16540 20936
rect 16488 20893 16497 20927
rect 16497 20893 16531 20927
rect 16531 20893 16540 20927
rect 16488 20884 16540 20893
rect 17224 20884 17276 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 20812 20952 20864 21004
rect 24308 21020 24360 21072
rect 26976 21063 27028 21072
rect 26976 21029 26985 21063
rect 26985 21029 27019 21063
rect 27019 21029 27028 21063
rect 26976 21020 27028 21029
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 19800 20884 19852 20936
rect 20076 20884 20128 20936
rect 3056 20748 3108 20800
rect 3884 20748 3936 20800
rect 4252 20748 4304 20800
rect 7288 20791 7340 20800
rect 7288 20757 7297 20791
rect 7297 20757 7331 20791
rect 7331 20757 7340 20791
rect 7288 20748 7340 20757
rect 9588 20748 9640 20800
rect 10876 20748 10928 20800
rect 15660 20816 15712 20868
rect 12900 20748 12952 20800
rect 13820 20748 13872 20800
rect 17040 20791 17092 20800
rect 17040 20757 17049 20791
rect 17049 20757 17083 20791
rect 17083 20757 17092 20791
rect 17040 20748 17092 20757
rect 17960 20791 18012 20800
rect 17960 20757 17969 20791
rect 17969 20757 18003 20791
rect 18003 20757 18012 20791
rect 17960 20748 18012 20757
rect 18236 20816 18288 20868
rect 20996 20748 21048 20800
rect 21364 20884 21416 20936
rect 23020 20952 23072 21004
rect 24124 20952 24176 21004
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 24032 20927 24084 20936
rect 24032 20893 24041 20927
rect 24041 20893 24075 20927
rect 24075 20893 24084 20927
rect 24032 20884 24084 20893
rect 25044 20952 25096 21004
rect 25780 20884 25832 20936
rect 26884 20884 26936 20936
rect 27528 20884 27580 20936
rect 27896 20927 27948 20936
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 27896 20884 27948 20893
rect 24032 20748 24084 20800
rect 27712 20816 27764 20868
rect 24860 20748 24912 20800
rect 27436 20791 27488 20800
rect 27436 20757 27445 20791
rect 27445 20757 27479 20791
rect 27479 20757 27488 20791
rect 27436 20748 27488 20757
rect 27620 20791 27672 20800
rect 27620 20757 27629 20791
rect 27629 20757 27663 20791
rect 27663 20757 27672 20791
rect 27620 20748 27672 20757
rect 28448 20748 28500 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 2596 20587 2648 20596
rect 2596 20553 2605 20587
rect 2605 20553 2639 20587
rect 2639 20553 2648 20587
rect 2596 20544 2648 20553
rect 3332 20544 3384 20596
rect 6920 20544 6972 20596
rect 7656 20544 7708 20596
rect 8392 20544 8444 20596
rect 3608 20476 3660 20528
rect 3240 20408 3292 20460
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 3884 20408 3936 20460
rect 5080 20476 5132 20528
rect 4344 20408 4396 20460
rect 2044 20383 2096 20392
rect 2044 20349 2053 20383
rect 2053 20349 2087 20383
rect 2087 20349 2096 20383
rect 2044 20340 2096 20349
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 4804 20408 4856 20460
rect 4988 20340 5040 20392
rect 6460 20408 6512 20460
rect 7288 20476 7340 20528
rect 8760 20408 8812 20460
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 11244 20476 11296 20528
rect 9588 20451 9640 20460
rect 9588 20417 9622 20451
rect 9622 20417 9640 20451
rect 9588 20408 9640 20417
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 10876 20408 10928 20460
rect 11796 20451 11848 20460
rect 11796 20417 11830 20451
rect 11830 20417 11848 20451
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 10324 20340 10376 20392
rect 2964 20204 3016 20256
rect 3332 20247 3384 20256
rect 3332 20213 3341 20247
rect 3341 20213 3375 20247
rect 3375 20213 3384 20247
rect 3332 20204 3384 20213
rect 3792 20247 3844 20256
rect 3792 20213 3801 20247
rect 3801 20213 3835 20247
rect 3835 20213 3844 20247
rect 3792 20204 3844 20213
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 4804 20204 4856 20256
rect 4896 20204 4948 20256
rect 5632 20247 5684 20256
rect 5632 20213 5641 20247
rect 5641 20213 5675 20247
rect 5675 20213 5684 20247
rect 5632 20204 5684 20213
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 6552 20204 6604 20256
rect 9128 20204 9180 20256
rect 10048 20204 10100 20256
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 10968 20247 11020 20256
rect 10968 20213 10977 20247
rect 10977 20213 11011 20247
rect 11011 20213 11020 20247
rect 10968 20204 11020 20213
rect 11796 20408 11848 20417
rect 13544 20544 13596 20596
rect 13544 20408 13596 20460
rect 14004 20408 14056 20460
rect 14648 20408 14700 20460
rect 15200 20544 15252 20596
rect 16488 20544 16540 20596
rect 17224 20544 17276 20596
rect 17500 20544 17552 20596
rect 18328 20544 18380 20596
rect 20260 20544 20312 20596
rect 19800 20476 19852 20528
rect 21180 20544 21232 20596
rect 21548 20544 21600 20596
rect 22284 20544 22336 20596
rect 24032 20587 24084 20596
rect 24032 20553 24041 20587
rect 24041 20553 24075 20587
rect 24075 20553 24084 20587
rect 24032 20544 24084 20553
rect 24308 20587 24360 20596
rect 24308 20553 24317 20587
rect 24317 20553 24351 20587
rect 24351 20553 24360 20587
rect 24308 20544 24360 20553
rect 24860 20544 24912 20596
rect 25044 20544 25096 20596
rect 27528 20544 27580 20596
rect 27712 20544 27764 20596
rect 21272 20476 21324 20528
rect 22836 20476 22888 20528
rect 23848 20519 23900 20528
rect 23848 20485 23857 20519
rect 23857 20485 23891 20519
rect 23891 20485 23900 20519
rect 23848 20476 23900 20485
rect 24676 20476 24728 20528
rect 16304 20408 16356 20460
rect 17040 20408 17092 20460
rect 17592 20451 17644 20460
rect 17592 20417 17601 20451
rect 17601 20417 17635 20451
rect 17635 20417 17644 20451
rect 17592 20408 17644 20417
rect 17960 20408 18012 20460
rect 12992 20272 13044 20324
rect 13360 20272 13412 20324
rect 14832 20315 14884 20324
rect 14832 20281 14841 20315
rect 14841 20281 14875 20315
rect 14875 20281 14884 20315
rect 15384 20383 15436 20392
rect 15384 20349 15393 20383
rect 15393 20349 15427 20383
rect 15427 20349 15436 20383
rect 15384 20340 15436 20349
rect 16856 20383 16908 20392
rect 16856 20349 16865 20383
rect 16865 20349 16899 20383
rect 16899 20349 16908 20383
rect 16856 20340 16908 20349
rect 18972 20383 19024 20392
rect 18972 20349 18981 20383
rect 18981 20349 19015 20383
rect 19015 20349 19024 20383
rect 18972 20340 19024 20349
rect 14832 20272 14884 20281
rect 12256 20204 12308 20256
rect 12716 20204 12768 20256
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 13728 20247 13780 20256
rect 13728 20213 13737 20247
rect 13737 20213 13771 20247
rect 13771 20213 13780 20247
rect 13728 20204 13780 20213
rect 13912 20204 13964 20256
rect 16580 20272 16632 20324
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 22284 20340 22336 20392
rect 20076 20272 20128 20324
rect 23112 20408 23164 20460
rect 23480 20408 23532 20460
rect 24768 20451 24820 20460
rect 24768 20417 24777 20451
rect 24777 20417 24811 20451
rect 24811 20417 24820 20451
rect 24768 20408 24820 20417
rect 26516 20451 26568 20460
rect 26516 20417 26525 20451
rect 26525 20417 26559 20451
rect 26559 20417 26568 20451
rect 26516 20408 26568 20417
rect 26884 20476 26936 20528
rect 27068 20408 27120 20460
rect 27436 20408 27488 20460
rect 27620 20408 27672 20460
rect 25596 20383 25648 20392
rect 25596 20349 25605 20383
rect 25605 20349 25639 20383
rect 25639 20349 25648 20383
rect 25596 20340 25648 20349
rect 25688 20340 25740 20392
rect 25780 20383 25832 20392
rect 25780 20349 25789 20383
rect 25789 20349 25823 20383
rect 25823 20349 25832 20383
rect 25780 20340 25832 20349
rect 26608 20340 26660 20392
rect 27712 20383 27764 20392
rect 27712 20349 27721 20383
rect 27721 20349 27755 20383
rect 27755 20349 27764 20383
rect 27712 20340 27764 20349
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 20536 20204 20588 20256
rect 21732 20204 21784 20256
rect 25964 20247 26016 20256
rect 25964 20213 25973 20247
rect 25973 20213 26007 20247
rect 26007 20213 26016 20247
rect 25964 20204 26016 20213
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 27528 20204 27580 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 2044 20000 2096 20052
rect 4252 20043 4304 20052
rect 4252 20009 4261 20043
rect 4261 20009 4295 20043
rect 4295 20009 4304 20043
rect 4252 20000 4304 20009
rect 4344 20000 4396 20052
rect 10784 20000 10836 20052
rect 13452 20000 13504 20052
rect 4712 19932 4764 19984
rect 4988 19932 5040 19984
rect 5448 19932 5500 19984
rect 8392 19932 8444 19984
rect 8760 19932 8812 19984
rect 9588 19932 9640 19984
rect 9956 19932 10008 19984
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 5080 19864 5132 19916
rect 6736 19864 6788 19916
rect 1400 19796 1452 19805
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 3056 19796 3108 19848
rect 3332 19796 3384 19848
rect 3516 19660 3568 19712
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 7288 19796 7340 19848
rect 10416 19864 10468 19916
rect 8208 19796 8260 19848
rect 4896 19771 4948 19780
rect 4896 19737 4905 19771
rect 4905 19737 4939 19771
rect 4939 19737 4948 19771
rect 4896 19728 4948 19737
rect 6000 19728 6052 19780
rect 6092 19728 6144 19780
rect 7196 19728 7248 19780
rect 9036 19796 9088 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 10508 19796 10560 19848
rect 10968 19771 11020 19780
rect 10968 19737 10977 19771
rect 10977 19737 11011 19771
rect 11011 19737 11020 19771
rect 10968 19728 11020 19737
rect 11336 19728 11388 19780
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 13912 19932 13964 19984
rect 14832 20043 14884 20052
rect 14832 20009 14841 20043
rect 14841 20009 14875 20043
rect 14875 20009 14884 20043
rect 14832 20000 14884 20009
rect 15384 20000 15436 20052
rect 16212 20000 16264 20052
rect 16856 20000 16908 20052
rect 17592 20000 17644 20052
rect 17960 20043 18012 20052
rect 17960 20009 17969 20043
rect 17969 20009 18003 20043
rect 18003 20009 18012 20043
rect 17960 20000 18012 20009
rect 20812 20000 20864 20052
rect 21640 20000 21692 20052
rect 15844 19975 15896 19984
rect 15844 19941 15853 19975
rect 15853 19941 15887 19975
rect 15887 19941 15896 19975
rect 15844 19932 15896 19941
rect 20904 19932 20956 19984
rect 21732 19932 21784 19984
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13820 19796 13872 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 16212 19796 16264 19848
rect 22376 19864 22428 19916
rect 23848 19864 23900 19916
rect 25780 20000 25832 20052
rect 25964 20000 26016 20052
rect 26332 20000 26384 20052
rect 26516 20000 26568 20052
rect 26976 20000 27028 20052
rect 27344 20000 27396 20052
rect 16304 19728 16356 19780
rect 17224 19796 17276 19848
rect 18052 19796 18104 19848
rect 8760 19660 8812 19669
rect 13084 19660 13136 19712
rect 15844 19660 15896 19712
rect 17224 19660 17276 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 21732 19796 21784 19848
rect 19616 19660 19668 19712
rect 21456 19728 21508 19780
rect 22560 19771 22612 19780
rect 22560 19737 22569 19771
rect 22569 19737 22603 19771
rect 22603 19737 22612 19771
rect 22560 19728 22612 19737
rect 25044 19864 25096 19916
rect 25320 19864 25372 19916
rect 23480 19728 23532 19780
rect 22468 19660 22520 19712
rect 22744 19660 22796 19712
rect 24860 19796 24912 19848
rect 27896 19932 27948 19984
rect 27160 19864 27212 19916
rect 26424 19728 26476 19780
rect 27528 19839 27580 19848
rect 27528 19805 27537 19839
rect 27537 19805 27571 19839
rect 27571 19805 27580 19839
rect 27528 19796 27580 19805
rect 27896 19839 27948 19848
rect 27896 19805 27905 19839
rect 27905 19805 27939 19839
rect 27939 19805 27948 19839
rect 27896 19796 27948 19805
rect 27252 19728 27304 19780
rect 27620 19728 27672 19780
rect 24308 19660 24360 19712
rect 24768 19703 24820 19712
rect 24768 19669 24777 19703
rect 24777 19669 24811 19703
rect 24811 19669 24820 19703
rect 24768 19660 24820 19669
rect 24952 19703 25004 19712
rect 24952 19669 24961 19703
rect 24961 19669 24995 19703
rect 24995 19669 25004 19703
rect 24952 19660 25004 19669
rect 25228 19703 25280 19712
rect 25228 19669 25237 19703
rect 25237 19669 25271 19703
rect 25271 19669 25280 19703
rect 25228 19660 25280 19669
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 27988 19703 28040 19712
rect 27988 19669 27997 19703
rect 27997 19669 28031 19703
rect 28031 19669 28040 19703
rect 27988 19660 28040 19669
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 1492 19456 1544 19508
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 3516 19499 3568 19508
rect 3516 19465 3525 19499
rect 3525 19465 3559 19499
rect 3559 19465 3568 19499
rect 3516 19456 3568 19465
rect 3792 19456 3844 19508
rect 3976 19456 4028 19508
rect 4896 19456 4948 19508
rect 5448 19456 5500 19508
rect 5632 19456 5684 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2228 19320 2280 19372
rect 3516 19320 3568 19372
rect 3700 19320 3752 19372
rect 4160 19320 4212 19372
rect 4252 19320 4304 19372
rect 4804 19320 4856 19372
rect 7748 19456 7800 19508
rect 9036 19456 9088 19508
rect 8300 19388 8352 19440
rect 9404 19388 9456 19440
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 7288 19320 7340 19372
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 10692 19456 10744 19508
rect 11336 19431 11388 19440
rect 11336 19397 11345 19431
rect 11345 19397 11379 19431
rect 11379 19397 11388 19431
rect 11336 19388 11388 19397
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 9864 19320 9916 19372
rect 7012 19227 7064 19236
rect 7012 19193 7021 19227
rect 7021 19193 7055 19227
rect 7055 19193 7064 19227
rect 7012 19184 7064 19193
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 12900 19456 12952 19508
rect 12992 19499 13044 19508
rect 12992 19465 13001 19499
rect 13001 19465 13035 19499
rect 13035 19465 13044 19499
rect 12992 19456 13044 19465
rect 15200 19456 15252 19508
rect 12440 19320 12492 19372
rect 13544 19320 13596 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14556 19388 14608 19440
rect 10324 19295 10376 19304
rect 10324 19261 10333 19295
rect 10333 19261 10367 19295
rect 10367 19261 10376 19295
rect 10324 19252 10376 19261
rect 11060 19184 11112 19236
rect 13176 19252 13228 19304
rect 13636 19295 13688 19304
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 13820 19252 13872 19304
rect 13728 19184 13780 19236
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 5448 19159 5500 19168
rect 5448 19125 5457 19159
rect 5457 19125 5491 19159
rect 5491 19125 5500 19159
rect 5448 19116 5500 19125
rect 6092 19159 6144 19168
rect 6092 19125 6101 19159
rect 6101 19125 6135 19159
rect 6135 19125 6144 19159
rect 6092 19116 6144 19125
rect 8300 19116 8352 19168
rect 8576 19116 8628 19168
rect 9036 19116 9088 19168
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 9864 19116 9916 19125
rect 14464 19295 14516 19304
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 14464 19252 14516 19261
rect 15384 19456 15436 19508
rect 18052 19499 18104 19508
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 19892 19456 19944 19508
rect 22468 19499 22520 19508
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 16304 19388 16356 19440
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 17316 19320 17368 19372
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18144 19320 18196 19329
rect 19616 19388 19668 19440
rect 23112 19388 23164 19440
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 20996 19320 21048 19372
rect 21364 19335 21365 19346
rect 21365 19335 21399 19346
rect 21399 19335 21416 19346
rect 15384 19116 15436 19168
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 21364 19294 21416 19335
rect 21456 19320 21508 19372
rect 25596 19388 25648 19440
rect 25780 19388 25832 19440
rect 18880 19184 18932 19236
rect 17592 19116 17644 19168
rect 20812 19116 20864 19168
rect 22836 19227 22888 19236
rect 22836 19193 22845 19227
rect 22845 19193 22879 19227
rect 22879 19193 22888 19227
rect 22836 19184 22888 19193
rect 25136 19320 25188 19372
rect 25228 19320 25280 19372
rect 27896 19388 27948 19440
rect 24400 19295 24452 19304
rect 24400 19261 24409 19295
rect 24409 19261 24443 19295
rect 24443 19261 24452 19295
rect 24400 19252 24452 19261
rect 24860 19252 24912 19304
rect 25044 19252 25096 19304
rect 26056 19184 26108 19236
rect 26700 19320 26752 19372
rect 27068 19320 27120 19372
rect 27528 19320 27580 19372
rect 27712 19295 27764 19304
rect 27712 19261 27721 19295
rect 27721 19261 27755 19295
rect 27755 19261 27764 19295
rect 27712 19252 27764 19261
rect 28080 19252 28132 19304
rect 28172 19252 28224 19304
rect 23940 19116 23992 19168
rect 24860 19159 24912 19168
rect 24860 19125 24869 19159
rect 24869 19125 24903 19159
rect 24903 19125 24912 19159
rect 24860 19116 24912 19125
rect 25596 19159 25648 19168
rect 25596 19125 25605 19159
rect 25605 19125 25639 19159
rect 25639 19125 25648 19159
rect 25596 19116 25648 19125
rect 26332 19159 26384 19168
rect 26332 19125 26341 19159
rect 26341 19125 26375 19159
rect 26375 19125 26384 19159
rect 26332 19116 26384 19125
rect 26516 19159 26568 19168
rect 26516 19125 26525 19159
rect 26525 19125 26559 19159
rect 26559 19125 26568 19159
rect 26516 19116 26568 19125
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 6460 18912 6512 18964
rect 10324 18912 10376 18964
rect 10508 18912 10560 18964
rect 11796 18912 11848 18964
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 12440 18912 12492 18921
rect 13084 18955 13136 18964
rect 13084 18921 13093 18955
rect 13093 18921 13127 18955
rect 13127 18921 13136 18955
rect 13084 18912 13136 18921
rect 14464 18912 14516 18964
rect 2872 18776 2924 18828
rect 2780 18708 2832 18760
rect 5172 18776 5224 18828
rect 6552 18776 6604 18828
rect 7012 18776 7064 18828
rect 7656 18776 7708 18828
rect 8944 18776 8996 18828
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 2320 18640 2372 18692
rect 4896 18708 4948 18760
rect 5448 18708 5500 18760
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 2504 18615 2556 18624
rect 2504 18581 2513 18615
rect 2513 18581 2547 18615
rect 2547 18581 2556 18615
rect 2504 18572 2556 18581
rect 4436 18615 4488 18624
rect 4436 18581 4445 18615
rect 4445 18581 4479 18615
rect 4479 18581 4488 18615
rect 4436 18572 4488 18581
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 8852 18708 8904 18760
rect 9864 18776 9916 18828
rect 7564 18640 7616 18692
rect 10140 18708 10192 18760
rect 11060 18708 11112 18760
rect 9864 18640 9916 18692
rect 11796 18640 11848 18692
rect 7472 18572 7524 18624
rect 8392 18615 8444 18624
rect 8392 18581 8401 18615
rect 8401 18581 8435 18615
rect 8435 18581 8444 18615
rect 8392 18572 8444 18581
rect 8484 18572 8536 18624
rect 10784 18572 10836 18624
rect 11060 18572 11112 18624
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13728 18708 13780 18760
rect 14648 18708 14700 18760
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 17868 18912 17920 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 23480 18955 23532 18964
rect 23480 18921 23489 18955
rect 23489 18921 23523 18955
rect 23523 18921 23532 18955
rect 23480 18912 23532 18921
rect 24768 18912 24820 18964
rect 24860 18912 24912 18964
rect 20444 18776 20496 18828
rect 20904 18819 20956 18828
rect 20904 18785 20913 18819
rect 20913 18785 20947 18819
rect 20947 18785 20956 18819
rect 20904 18776 20956 18785
rect 17592 18708 17644 18760
rect 18696 18708 18748 18760
rect 20996 18708 21048 18760
rect 25044 18887 25096 18896
rect 25044 18853 25053 18887
rect 25053 18853 25087 18887
rect 25087 18853 25096 18887
rect 25044 18844 25096 18853
rect 21456 18708 21508 18760
rect 24492 18776 24544 18828
rect 26332 18955 26384 18964
rect 26332 18921 26341 18955
rect 26341 18921 26375 18955
rect 26375 18921 26384 18955
rect 26332 18912 26384 18921
rect 26516 18776 26568 18828
rect 27528 18776 27580 18828
rect 27988 18776 28040 18828
rect 11980 18572 12032 18624
rect 13820 18572 13872 18624
rect 15292 18572 15344 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 22468 18640 22520 18692
rect 23756 18751 23808 18760
rect 23756 18717 23765 18751
rect 23765 18717 23799 18751
rect 23799 18717 23808 18751
rect 23756 18708 23808 18717
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 25320 18751 25372 18760
rect 25320 18717 25329 18751
rect 25329 18717 25363 18751
rect 25363 18717 25372 18751
rect 25320 18708 25372 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 21272 18572 21324 18624
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 22836 18572 22888 18624
rect 27252 18615 27304 18624
rect 27252 18581 27261 18615
rect 27261 18581 27295 18615
rect 27295 18581 27304 18615
rect 27252 18572 27304 18581
rect 28080 18615 28132 18624
rect 28080 18581 28089 18615
rect 28089 18581 28123 18615
rect 28123 18581 28132 18615
rect 28080 18572 28132 18581
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 2320 18368 2372 18420
rect 2504 18368 2556 18420
rect 2872 18368 2924 18420
rect 3976 18368 4028 18420
rect 4436 18368 4488 18420
rect 5724 18368 5776 18420
rect 6644 18368 6696 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 4804 18300 4856 18352
rect 5172 18300 5224 18352
rect 7472 18368 7524 18420
rect 8944 18368 8996 18420
rect 9312 18368 9364 18420
rect 10324 18368 10376 18420
rect 10784 18368 10836 18420
rect 12072 18368 12124 18420
rect 12440 18368 12492 18420
rect 13176 18411 13228 18420
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 15568 18368 15620 18420
rect 16028 18368 16080 18420
rect 17224 18368 17276 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 17868 18368 17920 18420
rect 3148 18207 3200 18216
rect 3148 18173 3157 18207
rect 3157 18173 3191 18207
rect 3191 18173 3200 18207
rect 3148 18164 3200 18173
rect 3976 18096 4028 18148
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 5448 18275 5500 18284
rect 5448 18241 5457 18275
rect 5457 18241 5491 18275
rect 5491 18241 5500 18275
rect 5448 18232 5500 18241
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 6092 18232 6144 18284
rect 7656 18232 7708 18284
rect 8668 18300 8720 18352
rect 7196 18164 7248 18216
rect 6736 18028 6788 18080
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 8944 18207 8996 18216
rect 8944 18173 8953 18207
rect 8953 18173 8987 18207
rect 8987 18173 8996 18207
rect 8944 18164 8996 18173
rect 9128 18164 9180 18216
rect 9956 18096 10008 18148
rect 10232 18232 10284 18284
rect 10600 18232 10652 18284
rect 11152 18232 11204 18284
rect 13728 18300 13780 18352
rect 13636 18232 13688 18284
rect 11888 18207 11940 18216
rect 11888 18173 11897 18207
rect 11897 18173 11931 18207
rect 11931 18173 11940 18207
rect 11888 18164 11940 18173
rect 12164 18164 12216 18216
rect 12440 18164 12492 18216
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 19892 18368 19944 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 19340 18300 19392 18352
rect 22192 18368 22244 18420
rect 22284 18368 22336 18420
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 23756 18368 23808 18420
rect 24400 18368 24452 18420
rect 24584 18368 24636 18420
rect 24952 18368 25004 18420
rect 25320 18368 25372 18420
rect 25596 18368 25648 18420
rect 20812 18232 20864 18284
rect 20904 18232 20956 18284
rect 21640 18232 21692 18284
rect 22100 18232 22152 18284
rect 22744 18232 22796 18284
rect 24308 18300 24360 18352
rect 28080 18368 28132 18420
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 24676 18232 24728 18241
rect 24952 18232 25004 18284
rect 11980 18096 12032 18148
rect 9036 18028 9088 18080
rect 13820 18096 13872 18148
rect 15844 18164 15896 18216
rect 17960 18207 18012 18216
rect 17960 18173 17969 18207
rect 17969 18173 18003 18207
rect 18003 18173 18012 18207
rect 17960 18164 18012 18173
rect 18052 18096 18104 18148
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 23756 18164 23808 18216
rect 23940 18164 23992 18216
rect 25136 18164 25188 18216
rect 27160 18232 27212 18284
rect 28356 18232 28408 18284
rect 27896 18207 27948 18216
rect 27896 18173 27905 18207
rect 27905 18173 27939 18207
rect 27939 18173 27948 18207
rect 27896 18164 27948 18173
rect 16488 18028 16540 18080
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 17776 18028 17828 18037
rect 23480 18028 23532 18080
rect 23848 18071 23900 18080
rect 23848 18037 23857 18071
rect 23857 18037 23891 18071
rect 23891 18037 23900 18071
rect 23848 18028 23900 18037
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 26884 18028 26936 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 3148 17824 3200 17876
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 6000 17824 6052 17876
rect 6644 17824 6696 17876
rect 6736 17824 6788 17876
rect 7288 17824 7340 17876
rect 8944 17824 8996 17876
rect 9128 17824 9180 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 3608 17620 3660 17672
rect 3976 17620 4028 17672
rect 4252 17620 4304 17672
rect 2320 17552 2372 17604
rect 6276 17620 6328 17672
rect 6736 17663 6788 17672
rect 6736 17629 6745 17663
rect 6745 17629 6779 17663
rect 6779 17629 6788 17663
rect 6736 17620 6788 17629
rect 7012 17552 7064 17604
rect 8484 17756 8536 17808
rect 8760 17799 8812 17808
rect 8760 17765 8769 17799
rect 8769 17765 8803 17799
rect 8803 17765 8812 17799
rect 8760 17756 8812 17765
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 8392 17688 8444 17740
rect 8208 17620 8260 17672
rect 10048 17824 10100 17876
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 15660 17824 15712 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 21548 17824 21600 17876
rect 23756 17824 23808 17876
rect 24860 17824 24912 17876
rect 27252 17824 27304 17876
rect 11336 17756 11388 17808
rect 14004 17756 14056 17808
rect 12716 17688 12768 17740
rect 16028 17688 16080 17740
rect 11612 17620 11664 17672
rect 12440 17663 12492 17672
rect 12440 17629 12449 17663
rect 12449 17629 12483 17663
rect 12483 17629 12492 17663
rect 12440 17620 12492 17629
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14004 17620 14056 17672
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14740 17620 14792 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 16488 17688 16540 17740
rect 18144 17756 18196 17808
rect 23572 17756 23624 17808
rect 23848 17756 23900 17808
rect 26332 17756 26384 17808
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 10232 17552 10284 17604
rect 11888 17552 11940 17604
rect 15476 17552 15528 17604
rect 17224 17552 17276 17604
rect 17776 17552 17828 17604
rect 7748 17484 7800 17536
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 11612 17484 11664 17536
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 13636 17484 13688 17536
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 18052 17484 18104 17536
rect 19616 17620 19668 17672
rect 20536 17620 20588 17672
rect 22008 17620 22060 17672
rect 26792 17688 26844 17740
rect 20720 17552 20772 17604
rect 19524 17484 19576 17536
rect 22192 17484 22244 17536
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 23480 17620 23532 17672
rect 23296 17552 23348 17604
rect 24768 17620 24820 17672
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 26240 17552 26292 17604
rect 26608 17595 26660 17604
rect 26608 17561 26617 17595
rect 26617 17561 26651 17595
rect 26651 17561 26660 17595
rect 26608 17552 26660 17561
rect 27436 17552 27488 17604
rect 23664 17527 23716 17536
rect 23664 17493 23673 17527
rect 23673 17493 23707 17527
rect 23707 17493 23716 17527
rect 23664 17484 23716 17493
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 28356 17527 28408 17536
rect 28356 17493 28365 17527
rect 28365 17493 28399 17527
rect 28399 17493 28408 17527
rect 28356 17484 28408 17493
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 3700 17280 3752 17332
rect 6828 17280 6880 17332
rect 1308 17144 1360 17196
rect 4344 17144 4396 17196
rect 2872 17076 2924 17128
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 4804 17076 4856 17128
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 7748 17212 7800 17264
rect 6460 17076 6512 17128
rect 7656 17144 7708 17196
rect 8392 17212 8444 17264
rect 9864 17280 9916 17332
rect 12164 17280 12216 17332
rect 12256 17280 12308 17332
rect 8300 17144 8352 17196
rect 4252 17008 4304 17060
rect 8576 17076 8628 17128
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 8852 17076 8904 17128
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 7472 17008 7524 17060
rect 6736 16940 6788 16992
rect 6920 16983 6972 16992
rect 6920 16949 6929 16983
rect 6929 16949 6963 16983
rect 6963 16949 6972 16983
rect 6920 16940 6972 16949
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 10600 17212 10652 17264
rect 11336 17212 11388 17264
rect 10140 17144 10192 17196
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 12624 17280 12676 17332
rect 13452 17280 13504 17332
rect 14280 17280 14332 17332
rect 15660 17280 15712 17332
rect 16120 17280 16172 17332
rect 17960 17280 18012 17332
rect 21088 17280 21140 17332
rect 23112 17280 23164 17332
rect 23664 17280 23716 17332
rect 23848 17323 23900 17332
rect 23848 17289 23857 17323
rect 23857 17289 23891 17323
rect 23891 17289 23900 17323
rect 23848 17280 23900 17289
rect 26424 17280 26476 17332
rect 13636 17144 13688 17196
rect 10600 17076 10652 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11796 17076 11848 17128
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 15476 17144 15528 17196
rect 15568 17119 15620 17128
rect 15568 17085 15577 17119
rect 15577 17085 15611 17119
rect 15611 17085 15620 17119
rect 15568 17076 15620 17085
rect 15660 17076 15712 17128
rect 16488 17144 16540 17196
rect 17776 17187 17828 17196
rect 17776 17153 17785 17187
rect 17785 17153 17819 17187
rect 17819 17153 17828 17187
rect 17776 17144 17828 17153
rect 20904 17212 20956 17264
rect 8208 16940 8260 16992
rect 8392 16940 8444 16992
rect 10600 16940 10652 16992
rect 19248 17144 19300 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 21364 17144 21416 17196
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 23296 17144 23348 17196
rect 26884 17212 26936 17264
rect 23756 17144 23808 17196
rect 25136 17144 25188 17196
rect 26056 17144 26108 17196
rect 26976 17187 27028 17196
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 27528 17144 27580 17196
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 20812 17008 20864 17060
rect 23480 17076 23532 17128
rect 28356 17280 28408 17332
rect 28080 17076 28132 17128
rect 15200 16940 15252 16992
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 19524 16940 19576 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 20904 16940 20956 16992
rect 23388 16940 23440 16992
rect 26516 16983 26568 16992
rect 26516 16949 26525 16983
rect 26525 16949 26559 16983
rect 26559 16949 26568 16983
rect 26516 16940 26568 16949
rect 27620 16940 27672 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 2872 16736 2924 16788
rect 1400 16600 1452 16652
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4344 16736 4396 16788
rect 7104 16736 7156 16788
rect 7564 16736 7616 16788
rect 6828 16668 6880 16720
rect 3332 16532 3384 16584
rect 3516 16532 3568 16584
rect 8944 16736 8996 16788
rect 9680 16736 9732 16788
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 6920 16532 6972 16584
rect 8392 16600 8444 16652
rect 8484 16600 8536 16652
rect 9864 16736 9916 16788
rect 10876 16736 10928 16788
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 11888 16736 11940 16788
rect 14464 16736 14516 16788
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11060 16668 11112 16720
rect 10048 16600 10100 16652
rect 10784 16600 10836 16652
rect 12716 16600 12768 16652
rect 15476 16779 15528 16788
rect 15476 16745 15485 16779
rect 15485 16745 15519 16779
rect 15519 16745 15528 16779
rect 15476 16736 15528 16745
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 16396 16736 16448 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 17316 16736 17368 16788
rect 17592 16736 17644 16788
rect 19616 16736 19668 16788
rect 19708 16736 19760 16788
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 10048 16464 10100 16516
rect 11244 16532 11296 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 13636 16532 13688 16584
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 14188 16532 14240 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 19340 16575 19392 16584
rect 19340 16541 19349 16575
rect 19349 16541 19383 16575
rect 19383 16541 19392 16575
rect 19340 16532 19392 16541
rect 19432 16532 19484 16584
rect 20628 16600 20680 16652
rect 22192 16736 22244 16788
rect 26240 16736 26292 16788
rect 27804 16736 27856 16788
rect 21456 16600 21508 16652
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20536 16532 20588 16584
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 21548 16532 21600 16541
rect 26332 16668 26384 16720
rect 27160 16600 27212 16652
rect 28632 16600 28684 16652
rect 11152 16464 11204 16516
rect 11428 16464 11480 16516
rect 11888 16464 11940 16516
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 7748 16396 7800 16448
rect 9772 16396 9824 16448
rect 11704 16396 11756 16448
rect 15292 16464 15344 16516
rect 16488 16464 16540 16516
rect 23388 16532 23440 16584
rect 14740 16396 14792 16448
rect 18972 16439 19024 16448
rect 18972 16405 18981 16439
rect 18981 16405 19015 16439
rect 19015 16405 19024 16439
rect 18972 16396 19024 16405
rect 20352 16396 20404 16448
rect 20904 16396 20956 16448
rect 21640 16439 21692 16448
rect 21640 16405 21649 16439
rect 21649 16405 21683 16439
rect 21683 16405 21692 16439
rect 21640 16396 21692 16405
rect 22376 16464 22428 16516
rect 22284 16396 22336 16448
rect 23020 16396 23072 16448
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 24584 16439 24636 16448
rect 24584 16405 24593 16439
rect 24593 16405 24627 16439
rect 24627 16405 24636 16439
rect 24584 16396 24636 16405
rect 24952 16396 25004 16448
rect 26884 16507 26936 16516
rect 26884 16473 26893 16507
rect 26893 16473 26927 16507
rect 26927 16473 26936 16507
rect 26884 16464 26936 16473
rect 28356 16464 28408 16516
rect 27804 16396 27856 16448
rect 28264 16396 28316 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 3332 16192 3384 16244
rect 3424 16192 3476 16244
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 2228 16056 2280 16108
rect 3700 16124 3752 16176
rect 7748 16192 7800 16244
rect 8484 16192 8536 16244
rect 9680 16192 9732 16244
rect 12624 16192 12676 16244
rect 3424 15988 3476 16040
rect 4160 15920 4212 15972
rect 7104 16124 7156 16176
rect 6920 16056 6972 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 10048 16124 10100 16176
rect 15200 16192 15252 16244
rect 15292 16192 15344 16244
rect 17224 16192 17276 16244
rect 19248 16192 19300 16244
rect 20260 16192 20312 16244
rect 20352 16192 20404 16244
rect 9772 16056 9824 16108
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 4804 15852 4856 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6736 15895 6788 15904
rect 6736 15861 6745 15895
rect 6745 15861 6779 15895
rect 6779 15861 6788 15895
rect 6736 15852 6788 15861
rect 7656 15852 7708 15904
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 10140 16031 10192 16040
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 12992 16056 13044 16108
rect 13268 16056 13320 16108
rect 9588 15852 9640 15904
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 11428 15852 11480 15904
rect 14096 16056 14148 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 13636 15988 13688 16040
rect 16212 16056 16264 16108
rect 17500 16056 17552 16108
rect 18144 16056 18196 16108
rect 15660 15988 15712 16040
rect 14556 15920 14608 15972
rect 14188 15852 14240 15904
rect 14924 15895 14976 15904
rect 14924 15861 14933 15895
rect 14933 15861 14967 15895
rect 14967 15861 14976 15895
rect 14924 15852 14976 15861
rect 19156 15988 19208 16040
rect 19432 15920 19484 15972
rect 20536 16192 20588 16244
rect 20812 16192 20864 16244
rect 21640 16192 21692 16244
rect 25044 16235 25096 16244
rect 25044 16201 25053 16235
rect 25053 16201 25087 16235
rect 25087 16201 25096 16235
rect 25044 16192 25096 16201
rect 26608 16192 26660 16244
rect 28540 16192 28592 16244
rect 22652 16124 22704 16176
rect 24952 16124 25004 16176
rect 21272 16056 21324 16108
rect 21456 16056 21508 16108
rect 21824 15988 21876 16040
rect 23388 16056 23440 16108
rect 24492 16056 24544 16108
rect 23020 15988 23072 16040
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 23572 15988 23624 16040
rect 25688 16056 25740 16108
rect 20628 15920 20680 15972
rect 20812 15920 20864 15972
rect 26332 16099 26384 16108
rect 26332 16065 26341 16099
rect 26341 16065 26375 16099
rect 26375 16065 26384 16099
rect 26332 16056 26384 16065
rect 26976 16056 27028 16108
rect 27160 16099 27212 16108
rect 27160 16065 27177 16099
rect 27177 16065 27211 16099
rect 27211 16065 27212 16099
rect 27160 16056 27212 16065
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 27436 16056 27488 16108
rect 15292 15852 15344 15904
rect 16672 15852 16724 15904
rect 17224 15852 17276 15904
rect 19340 15852 19392 15904
rect 24860 15920 24912 15972
rect 27068 15988 27120 16040
rect 27712 16031 27764 16040
rect 25964 15920 26016 15972
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 23572 15852 23624 15904
rect 24032 15895 24084 15904
rect 24032 15861 24041 15895
rect 24041 15861 24075 15895
rect 24075 15861 24084 15895
rect 24032 15852 24084 15861
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 26424 15895 26476 15904
rect 26424 15861 26433 15895
rect 26433 15861 26467 15895
rect 26467 15861 26476 15895
rect 26424 15852 26476 15861
rect 26792 15852 26844 15904
rect 27712 15997 27721 16031
rect 27721 15997 27755 16031
rect 27755 15997 27764 16031
rect 27712 15988 27764 15997
rect 28080 15895 28132 15904
rect 28080 15861 28089 15895
rect 28089 15861 28123 15895
rect 28123 15861 28132 15895
rect 28080 15852 28132 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6736 15648 6788 15700
rect 7748 15648 7800 15700
rect 8668 15648 8720 15700
rect 10140 15648 10192 15700
rect 10876 15648 10928 15700
rect 4160 15580 4212 15632
rect 3700 15512 3752 15564
rect 2228 15444 2280 15496
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 6368 15512 6420 15564
rect 8300 15512 8352 15564
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 5908 15444 5960 15496
rect 6184 15487 6236 15496
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 8484 15444 8536 15496
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 9588 15444 9640 15496
rect 12716 15648 12768 15700
rect 14924 15648 14976 15700
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 6920 15419 6972 15428
rect 6920 15385 6929 15419
rect 6929 15385 6963 15419
rect 6963 15385 6972 15419
rect 6920 15376 6972 15385
rect 7656 15419 7708 15428
rect 7656 15385 7665 15419
rect 7665 15385 7699 15419
rect 7699 15385 7708 15419
rect 7656 15376 7708 15385
rect 7748 15419 7800 15428
rect 7748 15385 7757 15419
rect 7757 15385 7791 15419
rect 7791 15385 7800 15419
rect 7748 15376 7800 15385
rect 11244 15444 11296 15496
rect 12164 15444 12216 15496
rect 15016 15580 15068 15632
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 3056 15308 3108 15360
rect 3976 15308 4028 15360
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 14832 15376 14884 15428
rect 17224 15444 17276 15496
rect 20536 15648 20588 15700
rect 21272 15691 21324 15700
rect 19156 15512 19208 15564
rect 19248 15512 19300 15564
rect 20628 15580 20680 15632
rect 21272 15657 21281 15691
rect 21281 15657 21315 15691
rect 21315 15657 21324 15691
rect 21272 15648 21324 15657
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 24032 15691 24084 15700
rect 24032 15657 24041 15691
rect 24041 15657 24075 15691
rect 24075 15657 24084 15691
rect 24032 15648 24084 15657
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 25780 15691 25832 15700
rect 25780 15657 25789 15691
rect 25789 15657 25823 15691
rect 25823 15657 25832 15691
rect 25780 15648 25832 15657
rect 25964 15648 26016 15700
rect 26424 15648 26476 15700
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 20812 15512 20864 15564
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 23204 15512 23256 15564
rect 24584 15512 24636 15564
rect 25596 15580 25648 15632
rect 19340 15376 19392 15428
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 22192 15444 22244 15496
rect 22468 15444 22520 15496
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 23020 15444 23072 15496
rect 11704 15308 11756 15360
rect 12072 15308 12124 15360
rect 14004 15308 14056 15360
rect 16120 15308 16172 15360
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 17592 15351 17644 15360
rect 17592 15317 17601 15351
rect 17601 15317 17635 15351
rect 17635 15317 17644 15351
rect 17592 15308 17644 15317
rect 18512 15308 18564 15360
rect 18972 15308 19024 15360
rect 21456 15376 21508 15428
rect 21824 15376 21876 15428
rect 23204 15376 23256 15428
rect 23940 15444 23992 15496
rect 26332 15512 26384 15564
rect 26700 15512 26752 15564
rect 28080 15648 28132 15700
rect 28356 15691 28408 15700
rect 28356 15657 28365 15691
rect 28365 15657 28399 15691
rect 28399 15657 28408 15691
rect 28356 15648 28408 15657
rect 27068 15580 27120 15632
rect 27620 15512 27672 15564
rect 27804 15555 27856 15564
rect 27804 15521 27813 15555
rect 27813 15521 27847 15555
rect 27847 15521 27856 15555
rect 27804 15512 27856 15521
rect 19984 15308 20036 15360
rect 20812 15351 20864 15360
rect 20812 15317 20821 15351
rect 20821 15317 20855 15351
rect 20855 15317 20864 15351
rect 20812 15308 20864 15317
rect 22928 15308 22980 15360
rect 23112 15351 23164 15360
rect 23112 15317 23121 15351
rect 23121 15317 23155 15351
rect 23155 15317 23164 15351
rect 23112 15308 23164 15317
rect 23480 15308 23532 15360
rect 24768 15308 24820 15360
rect 28356 15376 28408 15428
rect 26240 15308 26292 15360
rect 27344 15308 27396 15360
rect 27712 15308 27764 15360
rect 27804 15308 27856 15360
rect 28172 15308 28224 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 2228 15104 2280 15156
rect 4252 15104 4304 15156
rect 4712 15104 4764 15156
rect 5448 15104 5500 15156
rect 6184 15104 6236 15156
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 6552 15104 6604 15156
rect 2964 15036 3016 15088
rect 3976 15036 4028 15088
rect 7748 15104 7800 15156
rect 4068 14968 4120 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 3148 14764 3200 14816
rect 4804 14968 4856 15020
rect 5908 15011 5960 15020
rect 5908 14977 5917 15011
rect 5917 14977 5951 15011
rect 5951 14977 5960 15011
rect 5908 14968 5960 14977
rect 4344 14807 4396 14816
rect 4344 14773 4353 14807
rect 4353 14773 4387 14807
rect 4387 14773 4396 14807
rect 4344 14764 4396 14773
rect 4896 14764 4948 14816
rect 6368 14764 6420 14816
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 8300 15011 8352 15020
rect 8300 14977 8309 15011
rect 8309 14977 8343 15011
rect 8343 14977 8352 15011
rect 8300 14968 8352 14977
rect 12716 15036 12768 15088
rect 6736 14832 6788 14884
rect 6920 14832 6972 14884
rect 9496 14900 9548 14952
rect 13912 15104 13964 15156
rect 14556 15104 14608 15156
rect 15476 15104 15528 15156
rect 17224 15104 17276 15156
rect 10324 14900 10376 14952
rect 8484 14764 8536 14816
rect 10048 14764 10100 14816
rect 10692 14807 10744 14816
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 14464 15036 14516 15088
rect 18880 15104 18932 15156
rect 13728 15011 13780 15020
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 15384 14968 15436 15020
rect 15752 14968 15804 15020
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 15476 14900 15528 14952
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 17132 14875 17184 14884
rect 17132 14841 17141 14875
rect 17141 14841 17175 14875
rect 17175 14841 17184 14875
rect 17132 14832 17184 14841
rect 17592 14968 17644 15020
rect 18236 14900 18288 14952
rect 18512 14900 18564 14952
rect 19800 14968 19852 15020
rect 20812 15104 20864 15156
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 20720 15036 20772 15088
rect 21180 15036 21232 15088
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 19248 14900 19300 14952
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20168 14900 20220 14952
rect 21088 14968 21140 15020
rect 22376 15036 22428 15088
rect 25136 15036 25188 15088
rect 27712 15104 27764 15156
rect 27896 15104 27948 15156
rect 28448 15104 28500 15156
rect 26976 15036 27028 15088
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 21640 14900 21692 14952
rect 23388 14968 23440 15020
rect 24032 14968 24084 15020
rect 25780 14968 25832 15020
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 26608 14968 26660 15020
rect 27252 14968 27304 15020
rect 27528 14968 27580 15020
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 24400 14943 24452 14952
rect 24400 14909 24409 14943
rect 24409 14909 24443 14943
rect 24443 14909 24452 14943
rect 24400 14900 24452 14909
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 14096 14764 14148 14816
rect 17960 14807 18012 14816
rect 17960 14773 17969 14807
rect 17969 14773 18003 14807
rect 18003 14773 18012 14807
rect 17960 14764 18012 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 22928 14764 22980 14816
rect 24032 14764 24084 14816
rect 24952 14764 25004 14816
rect 26976 14807 27028 14816
rect 26976 14773 26985 14807
rect 26985 14773 27019 14807
rect 27019 14773 27028 14807
rect 26976 14764 27028 14773
rect 27620 14900 27672 14952
rect 28080 14807 28132 14816
rect 28080 14773 28089 14807
rect 28089 14773 28123 14807
rect 28123 14773 28132 14807
rect 28080 14764 28132 14773
rect 28540 14764 28592 14816
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 2872 14560 2924 14612
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 3332 14560 3384 14612
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 2964 14492 3016 14544
rect 3056 14424 3108 14476
rect 4160 14424 4212 14476
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 3240 14356 3292 14408
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 2320 14288 2372 14340
rect 4068 14288 4120 14340
rect 8024 14560 8076 14612
rect 10048 14560 10100 14612
rect 10692 14560 10744 14612
rect 12348 14560 12400 14612
rect 13728 14560 13780 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14004 14560 14056 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 18236 14560 18288 14612
rect 19156 14560 19208 14612
rect 20076 14560 20128 14612
rect 6368 14424 6420 14476
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 5356 14288 5408 14340
rect 5531 14331 5583 14340
rect 5531 14297 5563 14331
rect 5563 14297 5583 14331
rect 5531 14288 5583 14297
rect 7564 14288 7616 14340
rect 2044 14220 2096 14272
rect 5816 14220 5868 14272
rect 6736 14220 6788 14272
rect 8576 14220 8628 14272
rect 10232 14424 10284 14476
rect 10140 14356 10192 14408
rect 9956 14288 10008 14340
rect 10232 14220 10284 14272
rect 10324 14263 10376 14272
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 10876 14220 10928 14272
rect 12348 14424 12400 14476
rect 12164 14356 12216 14408
rect 13084 14356 13136 14408
rect 13452 14492 13504 14544
rect 16120 14492 16172 14544
rect 19432 14492 19484 14544
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 15292 14424 15344 14476
rect 17132 14424 17184 14476
rect 18144 14424 18196 14476
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 19156 14424 19208 14476
rect 20812 14560 20864 14612
rect 22008 14560 22060 14612
rect 22560 14560 22612 14612
rect 24400 14560 24452 14612
rect 22652 14492 22704 14544
rect 25872 14560 25924 14612
rect 26608 14603 26660 14612
rect 26608 14569 26617 14603
rect 26617 14569 26651 14603
rect 26651 14569 26660 14603
rect 26608 14560 26660 14569
rect 26976 14560 27028 14612
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 18788 14356 18840 14408
rect 18972 14356 19024 14408
rect 21272 14424 21324 14476
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 22284 14424 22336 14476
rect 25136 14424 25188 14476
rect 12256 14220 12308 14272
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 14188 14220 14240 14272
rect 15844 14220 15896 14272
rect 19432 14220 19484 14272
rect 21456 14288 21508 14340
rect 23020 14356 23072 14408
rect 23112 14356 23164 14408
rect 23204 14356 23256 14408
rect 24032 14356 24084 14408
rect 21640 14263 21692 14272
rect 21640 14229 21649 14263
rect 21649 14229 21683 14263
rect 21683 14229 21692 14263
rect 21640 14220 21692 14229
rect 25320 14356 25372 14408
rect 27344 14535 27396 14544
rect 27344 14501 27353 14535
rect 27353 14501 27387 14535
rect 27387 14501 27396 14535
rect 27344 14492 27396 14501
rect 27528 14424 27580 14476
rect 27804 14424 27856 14476
rect 24492 14331 24544 14340
rect 24492 14297 24501 14331
rect 24501 14297 24535 14331
rect 24535 14297 24544 14331
rect 24492 14288 24544 14297
rect 25228 14288 25280 14340
rect 26424 14288 26476 14340
rect 28172 14356 28224 14408
rect 28448 14288 28500 14340
rect 23296 14220 23348 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 2320 14016 2372 14068
rect 3700 14016 3752 14068
rect 4068 14016 4120 14068
rect 4804 14016 4856 14068
rect 7196 14016 7248 14068
rect 7564 14059 7616 14068
rect 7564 14025 7573 14059
rect 7573 14025 7607 14059
rect 7607 14025 7616 14059
rect 7564 14016 7616 14025
rect 8392 14016 8444 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12900 14016 12952 14068
rect 13360 14016 13412 14068
rect 14280 14016 14332 14068
rect 2780 13880 2832 13932
rect 4252 13948 4304 14000
rect 6920 13948 6972 14000
rect 7380 13948 7432 14000
rect 9496 13948 9548 14000
rect 4160 13880 4212 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 4988 13880 5040 13932
rect 5356 13880 5408 13932
rect 5908 13880 5960 13932
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 5632 13812 5684 13864
rect 6736 13812 6788 13864
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 10140 13948 10192 14000
rect 10968 13880 11020 13932
rect 14188 13948 14240 14000
rect 15844 14016 15896 14068
rect 15936 14016 15988 14068
rect 16028 14016 16080 14068
rect 7380 13744 7432 13796
rect 8116 13812 8168 13864
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10048 13812 10100 13821
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 13544 13923 13596 13932
rect 13544 13889 13578 13923
rect 13578 13889 13596 13923
rect 13544 13880 13596 13889
rect 16580 14016 16632 14068
rect 17408 14016 17460 14068
rect 17684 14016 17736 14068
rect 18972 13948 19024 14000
rect 9036 13744 9088 13796
rect 10508 13744 10560 13796
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 3608 13676 3660 13728
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 6092 13719 6144 13728
rect 6092 13685 6101 13719
rect 6101 13685 6135 13719
rect 6135 13685 6144 13719
rect 6092 13676 6144 13685
rect 7656 13719 7708 13728
rect 7656 13685 7665 13719
rect 7665 13685 7699 13719
rect 7699 13685 7708 13719
rect 7656 13676 7708 13685
rect 7840 13676 7892 13728
rect 7932 13676 7984 13728
rect 11060 13676 11112 13728
rect 11796 13812 11848 13864
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 18696 13880 18748 13932
rect 19984 13948 20036 14000
rect 20904 14016 20956 14068
rect 21456 14059 21508 14068
rect 21456 14025 21465 14059
rect 21465 14025 21499 14059
rect 21499 14025 21508 14059
rect 21456 14016 21508 14025
rect 27804 14016 27856 14068
rect 28356 14016 28408 14068
rect 18880 13812 18932 13864
rect 17960 13744 18012 13796
rect 19616 13923 19668 13932
rect 19616 13889 19625 13923
rect 19625 13889 19659 13923
rect 19659 13889 19668 13923
rect 19616 13880 19668 13889
rect 21456 13880 21508 13932
rect 22928 13880 22980 13932
rect 23020 13923 23072 13932
rect 23020 13889 23029 13923
rect 23029 13889 23063 13923
rect 23063 13889 23072 13923
rect 23020 13880 23072 13889
rect 21548 13812 21600 13864
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25780 13880 25832 13932
rect 26240 13880 26292 13932
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 27620 13948 27672 14000
rect 27068 13923 27120 13932
rect 27068 13889 27077 13923
rect 27077 13889 27111 13923
rect 27111 13889 27120 13923
rect 27068 13880 27120 13889
rect 28080 13880 28132 13932
rect 27344 13855 27396 13864
rect 27344 13821 27353 13855
rect 27353 13821 27387 13855
rect 27387 13821 27396 13855
rect 27344 13812 27396 13821
rect 27988 13855 28040 13864
rect 27988 13821 27997 13855
rect 27997 13821 28031 13855
rect 28031 13821 28040 13855
rect 27988 13812 28040 13821
rect 12440 13676 12492 13728
rect 16580 13676 16632 13728
rect 18972 13676 19024 13728
rect 19616 13676 19668 13728
rect 20536 13676 20588 13728
rect 22192 13744 22244 13796
rect 22836 13744 22888 13796
rect 28172 13812 28224 13864
rect 22560 13676 22612 13728
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 25320 13676 25372 13728
rect 25780 13719 25832 13728
rect 25780 13685 25789 13719
rect 25789 13685 25823 13719
rect 25823 13685 25832 13719
rect 25780 13676 25832 13685
rect 25964 13719 26016 13728
rect 25964 13685 25973 13719
rect 25973 13685 26007 13719
rect 26007 13685 26016 13719
rect 25964 13676 26016 13685
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 26608 13676 26660 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 2780 13472 2832 13524
rect 2872 13472 2924 13524
rect 4804 13515 4856 13524
rect 4804 13481 4813 13515
rect 4813 13481 4847 13515
rect 4847 13481 4856 13515
rect 4804 13472 4856 13481
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 5724 13472 5776 13524
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 8116 13472 8168 13524
rect 8484 13472 8536 13524
rect 9956 13515 10008 13524
rect 9956 13481 9965 13515
rect 9965 13481 9999 13515
rect 9999 13481 10008 13515
rect 9956 13472 10008 13481
rect 10416 13472 10468 13524
rect 10508 13472 10560 13524
rect 12532 13472 12584 13524
rect 13544 13472 13596 13524
rect 16028 13515 16080 13524
rect 16028 13481 16037 13515
rect 16037 13481 16071 13515
rect 16071 13481 16080 13515
rect 16028 13472 16080 13481
rect 19616 13515 19668 13524
rect 19616 13481 19625 13515
rect 19625 13481 19659 13515
rect 19659 13481 19668 13515
rect 19616 13472 19668 13481
rect 19892 13472 19944 13524
rect 20444 13472 20496 13524
rect 3240 13336 3292 13388
rect 5172 13336 5224 13388
rect 5356 13336 5408 13388
rect 6092 13336 6144 13388
rect 7656 13336 7708 13388
rect 940 13200 992 13252
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 2964 13268 3016 13320
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 3608 13200 3660 13252
rect 5540 13200 5592 13252
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 7840 13268 7892 13320
rect 8576 13268 8628 13320
rect 6276 13132 6328 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9220 13268 9272 13320
rect 10324 13336 10376 13388
rect 12348 13404 12400 13456
rect 12900 13336 12952 13388
rect 10508 13268 10560 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 10876 13268 10928 13320
rect 9680 13200 9732 13252
rect 9956 13200 10008 13252
rect 9220 13132 9272 13184
rect 10048 13132 10100 13184
rect 10784 13132 10836 13184
rect 11060 13132 11112 13184
rect 12164 13132 12216 13184
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 14648 13404 14700 13456
rect 13636 13268 13688 13320
rect 13452 13200 13504 13252
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 15292 13268 15344 13277
rect 15568 13200 15620 13252
rect 15752 13200 15804 13252
rect 17960 13268 18012 13320
rect 18236 13268 18288 13320
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 20996 13404 21048 13456
rect 24400 13472 24452 13524
rect 25044 13472 25096 13524
rect 25504 13515 25556 13524
rect 25504 13481 25513 13515
rect 25513 13481 25547 13515
rect 25547 13481 25556 13515
rect 25504 13472 25556 13481
rect 26424 13472 26476 13524
rect 27252 13472 27304 13524
rect 23848 13404 23900 13456
rect 23940 13404 23992 13456
rect 24676 13404 24728 13456
rect 28632 13404 28684 13456
rect 22284 13379 22336 13388
rect 22284 13345 22293 13379
rect 22293 13345 22327 13379
rect 22327 13345 22336 13379
rect 22284 13336 22336 13345
rect 24952 13336 25004 13388
rect 25964 13336 26016 13388
rect 26976 13336 27028 13388
rect 18788 13268 18840 13320
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 22744 13268 22796 13320
rect 23020 13311 23072 13320
rect 23020 13277 23029 13311
rect 23029 13277 23063 13311
rect 23063 13277 23072 13311
rect 23020 13268 23072 13277
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 23664 13268 23716 13320
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 21272 13200 21324 13252
rect 26240 13268 26292 13320
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 14280 13132 14332 13184
rect 17408 13132 17460 13184
rect 20260 13132 20312 13184
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 26516 13175 26568 13184
rect 26516 13141 26525 13175
rect 26525 13141 26559 13175
rect 26559 13141 26568 13175
rect 26516 13132 26568 13141
rect 27896 13200 27948 13252
rect 28080 13132 28132 13184
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 4160 12928 4212 12980
rect 4252 12928 4304 12980
rect 5632 12928 5684 12980
rect 6644 12928 6696 12980
rect 7564 12928 7616 12980
rect 9956 12928 10008 12980
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 5816 12860 5868 12912
rect 3884 12792 3936 12801
rect 6644 12792 6696 12844
rect 1400 12724 1452 12776
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 5080 12724 5132 12776
rect 5632 12724 5684 12776
rect 8024 12860 8076 12912
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7196 12792 7248 12844
rect 10508 12860 10560 12912
rect 10968 12928 11020 12980
rect 7380 12724 7432 12776
rect 5540 12588 5592 12640
rect 6276 12656 6328 12708
rect 7196 12656 7248 12708
rect 8392 12792 8444 12844
rect 8576 12792 8628 12844
rect 9680 12792 9732 12844
rect 9864 12724 9916 12776
rect 8576 12656 8628 12708
rect 10784 12792 10836 12844
rect 10876 12792 10928 12844
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 10968 12656 11020 12708
rect 11796 12724 11848 12776
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 12716 12928 12768 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13360 12928 13412 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 14096 12928 14148 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 14188 12860 14240 12912
rect 16580 12928 16632 12980
rect 16764 12928 16816 12980
rect 18328 12928 18380 12980
rect 20904 12928 20956 12980
rect 22192 12928 22244 12980
rect 22468 12928 22520 12980
rect 22652 12928 22704 12980
rect 23204 12928 23256 12980
rect 23756 12928 23808 12980
rect 23848 12928 23900 12980
rect 24400 12928 24452 12980
rect 26608 12928 26660 12980
rect 27252 12928 27304 12980
rect 28080 12928 28132 12980
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 12900 12724 12952 12776
rect 15752 12792 15804 12844
rect 17960 12835 18012 12844
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 17960 12792 18012 12801
rect 14280 12724 14332 12776
rect 13176 12656 13228 12708
rect 14096 12656 14148 12708
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 13912 12588 13964 12640
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 18880 12792 18932 12844
rect 21824 12860 21876 12912
rect 20260 12792 20312 12844
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 22928 12792 22980 12844
rect 23296 12792 23348 12844
rect 25780 12860 25832 12912
rect 24308 12792 24360 12844
rect 18144 12656 18196 12708
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 17960 12588 18012 12640
rect 18236 12588 18288 12640
rect 23664 12699 23716 12708
rect 23664 12665 23673 12699
rect 23673 12665 23707 12699
rect 23707 12665 23716 12699
rect 23664 12656 23716 12665
rect 23940 12656 23992 12708
rect 20812 12588 20864 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 22100 12631 22152 12640
rect 22100 12597 22109 12631
rect 22109 12597 22143 12631
rect 22143 12597 22152 12631
rect 22100 12588 22152 12597
rect 24952 12724 25004 12776
rect 27068 12767 27120 12776
rect 27068 12733 27077 12767
rect 27077 12733 27111 12767
rect 27111 12733 27120 12767
rect 27068 12724 27120 12733
rect 27712 12767 27764 12776
rect 27712 12733 27721 12767
rect 27721 12733 27755 12767
rect 27755 12733 27764 12767
rect 27712 12724 27764 12733
rect 26240 12656 26292 12708
rect 24768 12588 24820 12640
rect 26700 12631 26752 12640
rect 26700 12597 26709 12631
rect 26709 12597 26743 12631
rect 26743 12597 26752 12631
rect 26700 12588 26752 12597
rect 27436 12588 27488 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 3056 12384 3108 12436
rect 5356 12384 5408 12436
rect 2504 12248 2556 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3424 12180 3476 12232
rect 3700 12180 3752 12232
rect 4804 12180 4856 12232
rect 5264 12180 5316 12232
rect 6828 12384 6880 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 7748 12316 7800 12368
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 11704 12384 11756 12436
rect 12348 12384 12400 12436
rect 12808 12427 12860 12436
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 12992 12384 13044 12436
rect 4712 12112 4764 12164
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 6828 12180 6880 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 11244 12316 11296 12368
rect 9036 12248 9088 12300
rect 12808 12248 12860 12300
rect 6368 12112 6420 12164
rect 9772 12180 9824 12232
rect 9956 12223 10008 12232
rect 9956 12189 9990 12223
rect 9990 12189 10008 12223
rect 9956 12180 10008 12189
rect 10692 12180 10744 12232
rect 11980 12180 12032 12232
rect 14096 12316 14148 12368
rect 6920 12044 6972 12096
rect 8116 12044 8168 12096
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 12164 12044 12216 12096
rect 12440 12044 12492 12096
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 13544 12180 13596 12232
rect 14280 12180 14332 12232
rect 16764 12384 16816 12436
rect 18144 12384 18196 12436
rect 19248 12384 19300 12436
rect 19984 12384 20036 12436
rect 20720 12384 20772 12436
rect 16672 12316 16724 12368
rect 18788 12248 18840 12300
rect 14464 12112 14516 12164
rect 15292 12180 15344 12232
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 16212 12180 16264 12232
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 18052 12180 18104 12232
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 22100 12384 22152 12436
rect 24308 12384 24360 12436
rect 26332 12384 26384 12436
rect 21364 12359 21416 12368
rect 21364 12325 21373 12359
rect 21373 12325 21407 12359
rect 21407 12325 21416 12359
rect 21364 12316 21416 12325
rect 21456 12316 21508 12368
rect 23296 12223 23348 12232
rect 23296 12189 23305 12223
rect 23305 12189 23339 12223
rect 23339 12189 23348 12223
rect 23296 12180 23348 12189
rect 24124 12248 24176 12300
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 25596 12291 25648 12300
rect 25596 12257 25605 12291
rect 25605 12257 25639 12291
rect 25639 12257 25648 12291
rect 25596 12248 25648 12257
rect 26700 12248 26752 12300
rect 26792 12291 26844 12300
rect 26792 12257 26801 12291
rect 26801 12257 26835 12291
rect 26835 12257 26844 12291
rect 26792 12248 26844 12257
rect 27712 12291 27764 12300
rect 27712 12257 27721 12291
rect 27721 12257 27755 12291
rect 27755 12257 27764 12291
rect 27712 12248 27764 12257
rect 27988 12316 28040 12368
rect 14096 12044 14148 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 22744 12155 22796 12164
rect 22744 12121 22753 12155
rect 22753 12121 22787 12155
rect 22787 12121 22796 12155
rect 22744 12112 22796 12121
rect 25136 12112 25188 12164
rect 25504 12223 25556 12232
rect 25504 12189 25513 12223
rect 25513 12189 25547 12223
rect 25547 12189 25556 12223
rect 25504 12180 25556 12189
rect 26240 12112 26292 12164
rect 23572 12044 23624 12096
rect 24308 12044 24360 12096
rect 24492 12044 24544 12096
rect 25964 12044 26016 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 4712 11883 4764 11892
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 4988 11840 5040 11892
rect 5172 11840 5224 11892
rect 7012 11840 7064 11892
rect 7748 11840 7800 11892
rect 9680 11840 9732 11892
rect 10048 11840 10100 11892
rect 10692 11883 10744 11892
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 12808 11883 12860 11892
rect 12808 11849 12817 11883
rect 12817 11849 12851 11883
rect 12851 11849 12860 11883
rect 12808 11840 12860 11849
rect 2044 11815 2096 11824
rect 2044 11781 2053 11815
rect 2053 11781 2087 11815
rect 2087 11781 2096 11815
rect 2044 11772 2096 11781
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 4620 11772 4672 11824
rect 13452 11840 13504 11892
rect 14188 11840 14240 11892
rect 14280 11840 14332 11892
rect 14464 11840 14516 11892
rect 15568 11840 15620 11892
rect 16212 11840 16264 11892
rect 3424 11704 3476 11756
rect 2596 11568 2648 11620
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 4804 11679 4856 11688
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 7380 11636 7432 11688
rect 8484 11704 8536 11756
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11244 11704 11296 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 5448 11500 5500 11552
rect 6276 11500 6328 11552
rect 8300 11568 8352 11620
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 9864 11500 9916 11552
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 11060 11636 11112 11688
rect 12072 11636 12124 11688
rect 12808 11704 12860 11756
rect 13084 11704 13136 11756
rect 13544 11704 13596 11756
rect 17040 11840 17092 11892
rect 14464 11636 14516 11688
rect 19524 11772 19576 11824
rect 21272 11772 21324 11824
rect 21640 11772 21692 11824
rect 22008 11815 22060 11824
rect 22008 11781 22017 11815
rect 22017 11781 22051 11815
rect 22051 11781 22060 11815
rect 22008 11772 22060 11781
rect 23296 11772 23348 11824
rect 24032 11704 24084 11756
rect 27068 11840 27120 11892
rect 26424 11772 26476 11824
rect 19064 11636 19116 11688
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 22744 11679 22796 11688
rect 22744 11645 22753 11679
rect 22753 11645 22787 11679
rect 22787 11645 22796 11679
rect 22744 11636 22796 11645
rect 23664 11679 23716 11688
rect 23664 11645 23673 11679
rect 23673 11645 23707 11679
rect 23707 11645 23716 11679
rect 23664 11636 23716 11645
rect 23756 11636 23808 11688
rect 26976 11704 27028 11756
rect 28172 11883 28224 11892
rect 28172 11849 28181 11883
rect 28181 11849 28215 11883
rect 28215 11849 28224 11883
rect 28172 11840 28224 11849
rect 28448 11840 28500 11892
rect 27436 11747 27488 11756
rect 27436 11713 27445 11747
rect 27445 11713 27479 11747
rect 27479 11713 27488 11747
rect 27436 11704 27488 11713
rect 27988 11704 28040 11756
rect 28540 11704 28592 11756
rect 18696 11500 18748 11552
rect 23480 11568 23532 11620
rect 21640 11543 21692 11552
rect 21640 11509 21649 11543
rect 21649 11509 21683 11543
rect 21683 11509 21692 11543
rect 21640 11500 21692 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 27344 11636 27396 11688
rect 24860 11500 24912 11552
rect 26608 11500 26660 11552
rect 26792 11543 26844 11552
rect 26792 11509 26801 11543
rect 26801 11509 26835 11543
rect 26835 11509 26844 11543
rect 26792 11500 26844 11509
rect 27252 11543 27304 11552
rect 27252 11509 27261 11543
rect 27261 11509 27295 11543
rect 27295 11509 27304 11543
rect 27252 11500 27304 11509
rect 28080 11500 28132 11552
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 2596 11296 2648 11348
rect 2504 11160 2556 11212
rect 6644 11296 6696 11348
rect 6736 11296 6788 11348
rect 4712 11271 4764 11280
rect 4712 11237 4721 11271
rect 4721 11237 4755 11271
rect 4755 11237 4764 11271
rect 4712 11228 4764 11237
rect 5540 11228 5592 11280
rect 10140 11296 10192 11348
rect 11888 11296 11940 11348
rect 3424 11160 3476 11212
rect 3792 11160 3844 11212
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 2688 11092 2740 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 4252 11092 4304 11144
rect 6736 11160 6788 11212
rect 7840 11160 7892 11212
rect 5448 11092 5500 11144
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6184 11092 6236 11144
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 9588 11092 9640 11144
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 11152 11160 11204 11212
rect 10784 11092 10836 11144
rect 2596 10956 2648 11008
rect 8392 11024 8444 11076
rect 10968 11092 11020 11144
rect 14464 11228 14516 11280
rect 14648 11228 14700 11280
rect 12624 11092 12676 11144
rect 13176 11092 13228 11144
rect 14096 11092 14148 11144
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 17316 11160 17368 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17776 11092 17828 11144
rect 20904 11296 20956 11348
rect 22008 11296 22060 11348
rect 23664 11296 23716 11348
rect 24124 11339 24176 11348
rect 24124 11305 24133 11339
rect 24133 11305 24167 11339
rect 24167 11305 24176 11339
rect 24124 11296 24176 11305
rect 25596 11296 25648 11348
rect 24400 11228 24452 11280
rect 26608 11271 26660 11280
rect 26608 11237 26617 11271
rect 26617 11237 26651 11271
rect 26651 11237 26660 11271
rect 26608 11228 26660 11237
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 24860 11160 24912 11212
rect 4252 10956 4304 11008
rect 7104 10956 7156 11008
rect 7564 10956 7616 11008
rect 15660 11024 15712 11076
rect 20904 11092 20956 11144
rect 21640 11092 21692 11144
rect 23020 11092 23072 11144
rect 23572 11092 23624 11144
rect 24124 11092 24176 11144
rect 24492 11092 24544 11144
rect 24768 11092 24820 11144
rect 28264 11160 28316 11212
rect 26884 11092 26936 11144
rect 28172 11092 28224 11144
rect 26148 11024 26200 11076
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 17132 10956 17184 11008
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 18236 10956 18288 11008
rect 18788 10956 18840 11008
rect 21088 10956 21140 11008
rect 22284 10956 22336 11008
rect 24216 10956 24268 11008
rect 25044 10999 25096 11008
rect 25044 10965 25053 10999
rect 25053 10965 25087 10999
rect 25087 10965 25096 10999
rect 25044 10956 25096 10965
rect 27528 10956 27580 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 2964 10752 3016 10804
rect 3332 10752 3384 10804
rect 5356 10752 5408 10804
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 6092 10752 6144 10804
rect 6920 10752 6972 10804
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 10048 10752 10100 10804
rect 10140 10752 10192 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 12808 10752 12860 10804
rect 2412 10684 2464 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 3516 10616 3568 10668
rect 4804 10684 4856 10736
rect 6368 10684 6420 10736
rect 4252 10616 4304 10668
rect 4896 10616 4948 10668
rect 4988 10616 5040 10668
rect 5264 10616 5316 10668
rect 5540 10616 5592 10668
rect 7196 10616 7248 10668
rect 9864 10616 9916 10668
rect 5264 10480 5316 10532
rect 6092 10480 6144 10532
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 10784 10548 10836 10600
rect 14556 10752 14608 10804
rect 14648 10752 14700 10804
rect 16028 10752 16080 10804
rect 18144 10752 18196 10804
rect 19524 10752 19576 10804
rect 19708 10752 19760 10804
rect 11520 10548 11572 10600
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 12992 10616 13044 10668
rect 12624 10548 12676 10600
rect 12808 10548 12860 10600
rect 13728 10548 13780 10600
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 17132 10684 17184 10736
rect 18696 10684 18748 10736
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 4344 10412 4396 10464
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 7104 10412 7156 10464
rect 12348 10412 12400 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16764 10455 16816 10464
rect 16764 10421 16773 10455
rect 16773 10421 16807 10455
rect 16807 10421 16816 10455
rect 16764 10412 16816 10421
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 18236 10616 18288 10668
rect 21088 10684 21140 10736
rect 21640 10684 21692 10736
rect 22284 10684 22336 10736
rect 18052 10548 18104 10600
rect 18696 10548 18748 10600
rect 19156 10480 19208 10532
rect 19984 10548 20036 10600
rect 21456 10548 21508 10600
rect 23112 10727 23164 10736
rect 23112 10693 23121 10727
rect 23121 10693 23155 10727
rect 23155 10693 23164 10727
rect 23112 10684 23164 10693
rect 23296 10684 23348 10736
rect 24492 10752 24544 10804
rect 25044 10752 25096 10804
rect 26148 10752 26200 10804
rect 23940 10684 23992 10736
rect 23388 10616 23440 10668
rect 24952 10684 25004 10736
rect 26792 10684 26844 10736
rect 27344 10752 27396 10804
rect 25228 10616 25280 10668
rect 26424 10616 26476 10668
rect 26884 10616 26936 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 27252 10616 27304 10668
rect 28264 10659 28316 10668
rect 28264 10625 28273 10659
rect 28273 10625 28307 10659
rect 28307 10625 28316 10659
rect 28264 10616 28316 10625
rect 24492 10591 24544 10600
rect 24492 10557 24501 10591
rect 24501 10557 24535 10591
rect 24535 10557 24544 10591
rect 24492 10548 24544 10557
rect 24860 10548 24912 10600
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 19708 10412 19760 10464
rect 19800 10455 19852 10464
rect 19800 10421 19809 10455
rect 19809 10421 19843 10455
rect 19843 10421 19852 10455
rect 19800 10412 19852 10421
rect 21456 10412 21508 10464
rect 22100 10412 22152 10464
rect 24768 10480 24820 10532
rect 23572 10412 23624 10464
rect 27436 10480 27488 10532
rect 26700 10455 26752 10464
rect 26700 10421 26709 10455
rect 26709 10421 26743 10455
rect 26743 10421 26752 10455
rect 26700 10412 26752 10421
rect 27712 10412 27764 10464
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 2872 10208 2924 10260
rect 3332 10208 3384 10260
rect 2596 10072 2648 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 4344 10208 4396 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 5724 10208 5776 10260
rect 5908 10208 5960 10260
rect 7840 10251 7892 10260
rect 7840 10217 7849 10251
rect 7849 10217 7883 10251
rect 7883 10217 7892 10251
rect 7840 10208 7892 10217
rect 8024 10208 8076 10260
rect 11796 10208 11848 10260
rect 15292 10208 15344 10260
rect 7656 10140 7708 10192
rect 8392 10140 8444 10192
rect 5540 10072 5592 10124
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 5264 10004 5316 10056
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 5448 10004 5500 10056
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 2964 9936 3016 9988
rect 4436 9936 4488 9988
rect 7012 10004 7064 10056
rect 7564 10004 7616 10056
rect 7748 10004 7800 10056
rect 8484 10004 8536 10056
rect 13912 10140 13964 10192
rect 11888 10072 11940 10124
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 9772 9936 9824 9988
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 13728 10047 13780 10056
rect 13728 10013 13745 10047
rect 13745 10013 13779 10047
rect 13779 10013 13780 10047
rect 15384 10140 15436 10192
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 17224 10208 17276 10260
rect 17960 10208 18012 10260
rect 13728 10004 13780 10013
rect 16764 10072 16816 10124
rect 17224 10072 17276 10124
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 19432 10140 19484 10192
rect 19156 10072 19208 10124
rect 19708 10072 19760 10124
rect 16304 9936 16356 9988
rect 18236 9936 18288 9988
rect 18788 10004 18840 10056
rect 18972 10004 19024 10056
rect 19892 10004 19944 10056
rect 20904 10004 20956 10056
rect 18880 9936 18932 9988
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 5724 9868 5776 9920
rect 6920 9868 6972 9920
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7012 9868 7064 9877
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 11796 9868 11848 9920
rect 11888 9868 11940 9920
rect 14096 9868 14148 9920
rect 14556 9868 14608 9920
rect 17040 9868 17092 9920
rect 17684 9868 17736 9920
rect 18972 9868 19024 9920
rect 20720 9979 20772 9988
rect 20720 9945 20729 9979
rect 20729 9945 20763 9979
rect 20763 9945 20772 9979
rect 20720 9936 20772 9945
rect 22100 10208 22152 10260
rect 21364 10183 21416 10192
rect 21364 10149 21373 10183
rect 21373 10149 21407 10183
rect 21407 10149 21416 10183
rect 21364 10140 21416 10149
rect 21088 10047 21140 10056
rect 21088 10013 21097 10047
rect 21097 10013 21131 10047
rect 21131 10013 21140 10047
rect 21088 10004 21140 10013
rect 21640 10140 21692 10192
rect 21732 10072 21784 10124
rect 23204 10208 23256 10260
rect 24124 10208 24176 10260
rect 24492 10208 24544 10260
rect 27068 10208 27120 10260
rect 22192 10047 22244 10056
rect 22192 10013 22201 10047
rect 22201 10013 22235 10047
rect 22235 10013 22244 10047
rect 22192 10004 22244 10013
rect 23020 10072 23072 10124
rect 23112 10072 23164 10124
rect 25044 10072 25096 10124
rect 26148 10115 26200 10124
rect 26148 10081 26157 10115
rect 26157 10081 26191 10115
rect 26191 10081 26200 10115
rect 26148 10072 26200 10081
rect 26240 10072 26292 10124
rect 26700 10072 26752 10124
rect 28264 10072 28316 10124
rect 23296 10004 23348 10056
rect 23848 10047 23900 10056
rect 23848 10013 23857 10047
rect 23857 10013 23891 10047
rect 23891 10013 23900 10047
rect 23848 10004 23900 10013
rect 23940 10004 23992 10056
rect 24216 10004 24268 10056
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 23572 9936 23624 9988
rect 23480 9868 23532 9920
rect 24952 9868 25004 9920
rect 25136 9868 25188 9920
rect 25412 9868 25464 9920
rect 28540 9936 28592 9988
rect 27620 9868 27672 9920
rect 27804 9868 27856 9920
rect 28448 9911 28500 9920
rect 28448 9877 28457 9911
rect 28457 9877 28491 9911
rect 28491 9877 28500 9911
rect 28448 9868 28500 9877
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 2872 9664 2924 9716
rect 3056 9639 3108 9648
rect 3056 9605 3065 9639
rect 3065 9605 3099 9639
rect 3099 9605 3108 9639
rect 3056 9596 3108 9605
rect 5540 9664 5592 9716
rect 5632 9596 5684 9648
rect 6092 9639 6144 9648
rect 6092 9605 6101 9639
rect 6101 9605 6135 9639
rect 6135 9605 6144 9639
rect 6092 9596 6144 9605
rect 9588 9664 9640 9716
rect 11704 9664 11756 9716
rect 12532 9664 12584 9716
rect 8392 9596 8444 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 4436 9528 4488 9580
rect 4804 9528 4856 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 8668 9528 8720 9580
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 11796 9528 11848 9580
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 1768 9392 1820 9444
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 5356 9460 5408 9512
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 5264 9392 5316 9444
rect 6920 9392 6972 9444
rect 10048 9460 10100 9512
rect 10876 9460 10928 9512
rect 12716 9528 12768 9580
rect 13544 9528 13596 9580
rect 13912 9664 13964 9716
rect 14096 9664 14148 9716
rect 14648 9664 14700 9716
rect 16028 9528 16080 9580
rect 18880 9596 18932 9648
rect 20720 9664 20772 9716
rect 21180 9664 21232 9716
rect 21640 9664 21692 9716
rect 23756 9664 23808 9716
rect 23848 9664 23900 9716
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 17408 9528 17460 9580
rect 18144 9528 18196 9580
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 17684 9392 17736 9444
rect 19156 9528 19208 9580
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21272 9528 21324 9580
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 22744 9528 22796 9580
rect 22836 9571 22888 9580
rect 22836 9537 22845 9571
rect 22845 9537 22879 9571
rect 22879 9537 22888 9571
rect 22836 9528 22888 9537
rect 23204 9528 23256 9580
rect 23296 9528 23348 9580
rect 24952 9664 25004 9716
rect 24860 9596 24912 9648
rect 26700 9664 26752 9716
rect 27712 9664 27764 9716
rect 27988 9664 28040 9716
rect 28448 9664 28500 9716
rect 25964 9596 26016 9648
rect 19432 9460 19484 9512
rect 19524 9503 19576 9512
rect 19524 9469 19533 9503
rect 19533 9469 19567 9503
rect 19567 9469 19576 9503
rect 19524 9460 19576 9469
rect 20076 9460 20128 9512
rect 21732 9460 21784 9512
rect 22100 9503 22152 9512
rect 22100 9469 22109 9503
rect 22109 9469 22143 9503
rect 22143 9469 22152 9503
rect 22100 9460 22152 9469
rect 22284 9503 22336 9512
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 24952 9460 25004 9512
rect 2228 9324 2280 9376
rect 3608 9324 3660 9376
rect 3884 9324 3936 9376
rect 8484 9324 8536 9376
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 17224 9324 17276 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 19708 9324 19760 9376
rect 20352 9324 20404 9376
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 23112 9392 23164 9444
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 22744 9367 22796 9376
rect 22744 9333 22753 9367
rect 22753 9333 22787 9367
rect 22787 9333 22796 9367
rect 22744 9324 22796 9333
rect 25044 9324 25096 9376
rect 26332 9367 26384 9376
rect 26332 9333 26341 9367
rect 26341 9333 26375 9367
rect 26375 9333 26384 9367
rect 26332 9324 26384 9333
rect 26792 9571 26844 9580
rect 26792 9537 26801 9571
rect 26801 9537 26835 9571
rect 26835 9537 26844 9571
rect 26792 9528 26844 9537
rect 27068 9528 27120 9580
rect 27896 9596 27948 9648
rect 27344 9460 27396 9512
rect 27988 9392 28040 9444
rect 26700 9324 26752 9376
rect 26884 9324 26936 9376
rect 27068 9367 27120 9376
rect 27068 9333 27077 9367
rect 27077 9333 27111 9367
rect 27111 9333 27120 9367
rect 27068 9324 27120 9333
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 2136 9120 2188 9172
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 5356 9163 5408 9172
rect 5356 9129 5365 9163
rect 5365 9129 5399 9163
rect 5399 9129 5408 9163
rect 5356 9120 5408 9129
rect 7380 9120 7432 9172
rect 8300 9120 8352 9172
rect 9036 9120 9088 9172
rect 9220 9120 9272 9172
rect 10048 9120 10100 9172
rect 10600 9120 10652 9172
rect 13176 9120 13228 9172
rect 14096 9120 14148 9172
rect 15108 9120 15160 9172
rect 15844 9120 15896 9172
rect 17316 9120 17368 9172
rect 18052 9120 18104 9172
rect 18788 9120 18840 9172
rect 19524 9120 19576 9172
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 2228 8916 2280 8968
rect 3884 8984 3936 9036
rect 4252 8984 4304 9036
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 2780 8780 2832 8832
rect 6368 9052 6420 9104
rect 7196 9095 7248 9104
rect 7196 9061 7205 9095
rect 7205 9061 7239 9095
rect 7239 9061 7248 9095
rect 7196 9052 7248 9061
rect 5264 8984 5316 9036
rect 6920 8984 6972 9036
rect 8484 9052 8536 9104
rect 7564 8984 7616 9036
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5356 8916 5408 8968
rect 6828 8916 6880 8968
rect 8668 8916 8720 8968
rect 5724 8848 5776 8900
rect 7472 8891 7524 8900
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 10416 8916 10468 8968
rect 12716 9052 12768 9104
rect 11888 8984 11940 9036
rect 21640 9120 21692 9172
rect 22100 9120 22152 9172
rect 22744 9120 22796 9172
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 25136 9120 25188 9172
rect 14188 9052 14240 9104
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 11704 8916 11756 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 15936 8916 15988 8968
rect 16304 8916 16356 8968
rect 16488 8916 16540 8968
rect 16580 8916 16632 8968
rect 16856 8984 16908 9036
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 19616 8984 19668 9036
rect 19708 8984 19760 9036
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 16028 8848 16080 8900
rect 8392 8780 8444 8832
rect 8576 8780 8628 8832
rect 9036 8780 9088 8832
rect 10508 8780 10560 8832
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 16856 8780 16908 8832
rect 17500 8780 17552 8832
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 17868 8780 17920 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19616 8823 19668 8832
rect 19616 8789 19625 8823
rect 19625 8789 19659 8823
rect 19659 8789 19668 8823
rect 19616 8780 19668 8789
rect 19708 8823 19760 8832
rect 19708 8789 19717 8823
rect 19717 8789 19751 8823
rect 19751 8789 19760 8823
rect 19708 8780 19760 8789
rect 20628 9052 20680 9104
rect 20168 8984 20220 9036
rect 20720 8984 20772 9036
rect 23112 8984 23164 9036
rect 23480 9052 23532 9104
rect 26608 9120 26660 9172
rect 27068 9120 27120 9172
rect 27620 9163 27672 9172
rect 27620 9129 27629 9163
rect 27629 9129 27663 9163
rect 27663 9129 27672 9163
rect 27620 9120 27672 9129
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 20076 8959 20128 8968
rect 20076 8925 20085 8959
rect 20085 8925 20119 8959
rect 20119 8925 20128 8959
rect 20076 8916 20128 8925
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 21548 8916 21600 8968
rect 21640 8916 21692 8968
rect 20720 8848 20772 8900
rect 20996 8848 21048 8900
rect 22468 8916 22520 8968
rect 24860 8984 24912 9036
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 24768 8916 24820 8968
rect 27620 8916 27672 8968
rect 27804 8916 27856 8968
rect 24400 8848 24452 8900
rect 24860 8848 24912 8900
rect 22008 8780 22060 8832
rect 22560 8780 22612 8832
rect 23020 8780 23072 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 26884 8780 26936 8832
rect 28356 8823 28408 8832
rect 28356 8789 28365 8823
rect 28365 8789 28399 8823
rect 28399 8789 28408 8823
rect 28356 8780 28408 8789
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1584 8576 1636 8628
rect 1768 8576 1820 8628
rect 1860 8576 1912 8628
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 4160 8576 4212 8628
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 4252 8508 4304 8560
rect 7472 8576 7524 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11060 8576 11112 8628
rect 11704 8576 11756 8628
rect 2780 8372 2832 8424
rect 4344 8440 4396 8492
rect 7012 8508 7064 8560
rect 7656 8508 7708 8560
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 3608 8304 3660 8356
rect 5816 8304 5868 8356
rect 8944 8440 8996 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 6368 8304 6420 8356
rect 7472 8372 7524 8424
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8576 8304 8628 8356
rect 9312 8347 9364 8356
rect 9312 8313 9321 8347
rect 9321 8313 9355 8347
rect 9355 8313 9364 8347
rect 9312 8304 9364 8313
rect 9680 8508 9732 8560
rect 10324 8508 10376 8560
rect 14280 8576 14332 8628
rect 16488 8576 16540 8628
rect 18696 8576 18748 8628
rect 19708 8576 19760 8628
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 10968 8440 11020 8492
rect 10508 8372 10560 8424
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11152 8372 11204 8424
rect 12164 8440 12216 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14096 8440 14148 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17776 8440 17828 8492
rect 17868 8440 17920 8492
rect 18236 8508 18288 8560
rect 19340 8508 19392 8560
rect 19432 8508 19484 8560
rect 19984 8551 20036 8560
rect 19984 8517 19993 8551
rect 19993 8517 20027 8551
rect 20027 8517 20036 8551
rect 19984 8508 20036 8517
rect 20076 8508 20128 8560
rect 20536 8576 20588 8628
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 20720 8508 20772 8560
rect 22192 8576 22244 8628
rect 22560 8576 22612 8628
rect 23480 8576 23532 8628
rect 24584 8576 24636 8628
rect 26332 8576 26384 8628
rect 28356 8576 28408 8628
rect 20996 8440 21048 8492
rect 17408 8372 17460 8424
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22468 8440 22520 8492
rect 22744 8440 22796 8492
rect 23940 8508 23992 8560
rect 24768 8508 24820 8560
rect 24860 8508 24912 8560
rect 25044 8551 25096 8560
rect 25044 8517 25053 8551
rect 25053 8517 25087 8551
rect 25087 8517 25096 8551
rect 25044 8508 25096 8517
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 15660 8304 15712 8356
rect 22928 8372 22980 8424
rect 23204 8415 23256 8424
rect 23204 8381 23213 8415
rect 23213 8381 23247 8415
rect 23247 8381 23256 8415
rect 23204 8372 23256 8381
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 26976 8440 27028 8492
rect 25780 8372 25832 8424
rect 3056 8236 3108 8288
rect 5080 8236 5132 8288
rect 7288 8236 7340 8288
rect 10232 8236 10284 8288
rect 12716 8279 12768 8288
rect 12716 8245 12725 8279
rect 12725 8245 12759 8279
rect 12759 8245 12768 8279
rect 12716 8236 12768 8245
rect 14648 8236 14700 8288
rect 15844 8279 15896 8288
rect 15844 8245 15853 8279
rect 15853 8245 15887 8279
rect 15887 8245 15896 8279
rect 15844 8236 15896 8245
rect 17868 8236 17920 8288
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 23388 8304 23440 8356
rect 23572 8347 23624 8356
rect 23572 8313 23581 8347
rect 23581 8313 23615 8347
rect 23615 8313 23624 8347
rect 23572 8304 23624 8313
rect 21456 8236 21508 8288
rect 22468 8236 22520 8288
rect 22652 8236 22704 8288
rect 26884 8372 26936 8424
rect 27896 8372 27948 8424
rect 27988 8415 28040 8424
rect 27988 8381 27997 8415
rect 27997 8381 28031 8415
rect 28031 8381 28040 8415
rect 27988 8372 28040 8381
rect 25964 8279 26016 8288
rect 25964 8245 25973 8279
rect 25973 8245 26007 8279
rect 26007 8245 26016 8279
rect 25964 8236 26016 8245
rect 26148 8236 26200 8288
rect 27528 8279 27580 8288
rect 27528 8245 27537 8279
rect 27537 8245 27571 8279
rect 27571 8245 27580 8279
rect 27528 8236 27580 8245
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 3608 8032 3660 8084
rect 4252 8032 4304 8084
rect 4896 7964 4948 8016
rect 10048 8032 10100 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 14556 8032 14608 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16764 8032 16816 8084
rect 18788 8032 18840 8084
rect 19064 8032 19116 8084
rect 20076 8032 20128 8084
rect 7012 8007 7064 8016
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 3240 7803 3292 7812
rect 3240 7769 3249 7803
rect 3249 7769 3283 7803
rect 3283 7769 3292 7803
rect 3240 7760 3292 7769
rect 3792 7828 3844 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 5080 7896 5132 7948
rect 7012 7973 7021 8007
rect 7021 7973 7055 8007
rect 7055 7973 7064 8007
rect 7012 7964 7064 7973
rect 7380 7964 7432 8016
rect 6000 7896 6052 7948
rect 9588 7964 9640 8016
rect 9312 7896 9364 7948
rect 10968 7896 11020 7948
rect 11888 7896 11940 7948
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6368 7828 6420 7880
rect 6736 7828 6788 7880
rect 7104 7760 7156 7812
rect 8576 7828 8628 7880
rect 9588 7760 9640 7812
rect 9772 7871 9824 7882
rect 9772 7837 9788 7871
rect 9788 7837 9822 7871
rect 9822 7837 9824 7871
rect 9772 7830 9824 7837
rect 11152 7828 11204 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 13728 7896 13780 7948
rect 4344 7692 4396 7744
rect 5172 7692 5224 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 5908 7692 5960 7744
rect 7288 7692 7340 7744
rect 7472 7692 7524 7744
rect 9036 7692 9088 7744
rect 12440 7760 12492 7812
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14004 7828 14056 7880
rect 14280 7828 14332 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14556 7828 14608 7880
rect 16212 7828 16264 7880
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17868 7964 17920 8016
rect 17776 7828 17828 7880
rect 19064 7896 19116 7948
rect 20076 7896 20128 7948
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 19708 7828 19760 7880
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 13176 7692 13228 7744
rect 15200 7692 15252 7744
rect 16120 7692 16172 7744
rect 18236 7760 18288 7812
rect 20628 8032 20680 8084
rect 20720 8032 20772 8084
rect 22008 8032 22060 8084
rect 22836 8032 22888 8084
rect 23112 8032 23164 8084
rect 23204 8032 23256 8084
rect 24584 8032 24636 8084
rect 24768 8075 24820 8084
rect 24768 8041 24777 8075
rect 24777 8041 24811 8075
rect 24811 8041 24820 8075
rect 24768 8032 24820 8041
rect 25320 8032 25372 8084
rect 26148 8032 26200 8084
rect 28080 8032 28132 8084
rect 17224 7692 17276 7744
rect 18420 7692 18472 7744
rect 18512 7692 18564 7744
rect 19524 7692 19576 7744
rect 20812 7828 20864 7880
rect 21272 7896 21324 7948
rect 21456 7964 21508 8016
rect 23204 7896 23256 7948
rect 22192 7828 22244 7880
rect 24032 7896 24084 7948
rect 24216 7896 24268 7948
rect 20904 7692 20956 7744
rect 20996 7735 21048 7744
rect 20996 7701 21005 7735
rect 21005 7701 21039 7735
rect 21039 7701 21048 7735
rect 20996 7692 21048 7701
rect 21180 7692 21232 7744
rect 22744 7735 22796 7744
rect 22744 7701 22753 7735
rect 22753 7701 22787 7735
rect 22787 7701 22796 7735
rect 22744 7692 22796 7701
rect 22928 7735 22980 7744
rect 22928 7701 22937 7735
rect 22937 7701 22971 7735
rect 22971 7701 22980 7735
rect 22928 7692 22980 7701
rect 23848 7828 23900 7880
rect 24492 7828 24544 7880
rect 24124 7692 24176 7744
rect 27436 7964 27488 8016
rect 28172 7964 28224 8016
rect 24952 7939 25004 7948
rect 24952 7905 24961 7939
rect 24961 7905 24995 7939
rect 24995 7905 25004 7939
rect 24952 7896 25004 7905
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 25964 7828 26016 7880
rect 26700 7871 26752 7880
rect 26700 7837 26709 7871
rect 26709 7837 26743 7871
rect 26743 7837 26752 7871
rect 26700 7828 26752 7837
rect 26792 7828 26844 7880
rect 28632 7828 28684 7880
rect 26148 7692 26200 7744
rect 28356 7735 28408 7744
rect 28356 7701 28365 7735
rect 28365 7701 28399 7735
rect 28399 7701 28408 7735
rect 28356 7692 28408 7701
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1584 7488 1636 7540
rect 3516 7488 3568 7540
rect 4620 7488 4672 7540
rect 6092 7488 6144 7540
rect 3792 7420 3844 7472
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 4160 7352 4212 7404
rect 4988 7352 5040 7404
rect 5908 7352 5960 7404
rect 4344 7284 4396 7336
rect 5264 7284 5316 7336
rect 6368 7352 6420 7404
rect 10600 7488 10652 7540
rect 11244 7488 11296 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 14648 7488 14700 7540
rect 15200 7488 15252 7540
rect 7472 7420 7524 7472
rect 9772 7420 9824 7472
rect 9864 7463 9916 7472
rect 9864 7429 9873 7463
rect 9873 7429 9907 7463
rect 9907 7429 9916 7463
rect 9864 7420 9916 7429
rect 10692 7420 10744 7472
rect 8300 7352 8352 7404
rect 9036 7352 9088 7404
rect 9588 7352 9640 7404
rect 13176 7420 13228 7472
rect 13452 7352 13504 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15752 7488 15804 7540
rect 16212 7488 16264 7540
rect 17684 7488 17736 7540
rect 18604 7488 18656 7540
rect 19708 7531 19760 7540
rect 19708 7497 19717 7531
rect 19717 7497 19751 7531
rect 19751 7497 19760 7531
rect 19708 7488 19760 7497
rect 20260 7488 20312 7540
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 17316 7420 17368 7472
rect 3884 7216 3936 7268
rect 4896 7216 4948 7268
rect 6736 7216 6788 7268
rect 6920 7148 6972 7200
rect 7104 7148 7156 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 12072 7284 12124 7336
rect 11152 7148 11204 7200
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 17132 7284 17184 7336
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 17684 7284 17736 7336
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 17316 7216 17368 7268
rect 19156 7420 19208 7472
rect 19340 7420 19392 7472
rect 21180 7488 21232 7540
rect 21272 7488 21324 7540
rect 21364 7488 21416 7540
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 18420 7352 18472 7404
rect 18512 7284 18564 7336
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 20076 7352 20128 7404
rect 22192 7488 22244 7540
rect 21640 7420 21692 7472
rect 22652 7488 22704 7540
rect 22744 7488 22796 7540
rect 23480 7488 23532 7540
rect 23848 7488 23900 7540
rect 24492 7488 24544 7540
rect 25780 7488 25832 7540
rect 19524 7216 19576 7268
rect 19708 7216 19760 7268
rect 22284 7284 22336 7336
rect 21088 7148 21140 7200
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 21548 7148 21600 7200
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 25688 7395 25740 7404
rect 23388 7284 23440 7336
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 25412 7284 25464 7336
rect 25688 7361 25697 7395
rect 25697 7361 25731 7395
rect 25731 7361 25740 7395
rect 25688 7352 25740 7361
rect 25780 7352 25832 7404
rect 26148 7395 26200 7404
rect 26148 7361 26157 7395
rect 26157 7361 26191 7395
rect 26191 7361 26200 7395
rect 26148 7352 26200 7361
rect 27436 7395 27488 7404
rect 27436 7361 27445 7395
rect 27445 7361 27479 7395
rect 27479 7361 27488 7395
rect 27436 7352 27488 7361
rect 25320 7148 25372 7200
rect 25872 7148 25924 7200
rect 26056 7148 26108 7200
rect 27896 7191 27948 7200
rect 27896 7157 27905 7191
rect 27905 7157 27939 7191
rect 27939 7157 27948 7191
rect 27896 7148 27948 7157
rect 28264 7191 28316 7200
rect 28264 7157 28273 7191
rect 28273 7157 28307 7191
rect 28307 7157 28316 7191
rect 28264 7148 28316 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 3792 6944 3844 6996
rect 4160 6987 4212 6996
rect 4160 6953 4169 6987
rect 4169 6953 4203 6987
rect 4203 6953 4212 6987
rect 4160 6944 4212 6953
rect 5264 6944 5316 6996
rect 4344 6876 4396 6928
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 7012 6944 7064 6996
rect 8300 6944 8352 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 12256 6944 12308 6996
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 12440 6944 12492 6953
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 14556 6944 14608 6996
rect 15568 6987 15620 6996
rect 15568 6953 15577 6987
rect 15577 6953 15611 6987
rect 15611 6953 15620 6987
rect 15568 6944 15620 6953
rect 15936 6944 15988 6996
rect 16028 6944 16080 6996
rect 18144 6944 18196 6996
rect 19892 6944 19944 6996
rect 3240 6808 3292 6860
rect 3884 6808 3936 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 6920 6808 6972 6860
rect 2780 6740 2832 6792
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 3516 6740 3568 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 8116 6740 8168 6792
rect 8760 6740 8812 6792
rect 6368 6672 6420 6724
rect 6736 6672 6788 6724
rect 9036 6672 9088 6724
rect 9588 6740 9640 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11060 6808 11112 6860
rect 12348 6876 12400 6928
rect 13452 6876 13504 6928
rect 11980 6808 12032 6860
rect 17960 6876 18012 6928
rect 18052 6876 18104 6928
rect 21548 6944 21600 6996
rect 22192 6944 22244 6996
rect 23848 6944 23900 6996
rect 26240 6944 26292 6996
rect 26608 6944 26660 6996
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 2872 6604 2924 6656
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 4160 6604 4212 6656
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 9496 6604 9548 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 11980 6672 12032 6724
rect 12072 6672 12124 6724
rect 13636 6740 13688 6792
rect 14004 6740 14056 6792
rect 14280 6740 14332 6792
rect 14464 6740 14516 6792
rect 14096 6604 14148 6656
rect 15108 6672 15160 6724
rect 15844 6740 15896 6792
rect 16580 6808 16632 6860
rect 16580 6715 16632 6724
rect 16580 6681 16589 6715
rect 16589 6681 16623 6715
rect 16623 6681 16632 6715
rect 16580 6672 16632 6681
rect 16764 6672 16816 6724
rect 17040 6783 17092 6792
rect 17040 6749 17073 6783
rect 17073 6749 17092 6783
rect 17592 6808 17644 6860
rect 18604 6808 18656 6860
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 21456 6808 21508 6860
rect 22284 6919 22336 6928
rect 22284 6885 22293 6919
rect 22293 6885 22327 6919
rect 22327 6885 22336 6919
rect 22284 6876 22336 6885
rect 23388 6876 23440 6928
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 22928 6808 22980 6860
rect 23572 6851 23624 6860
rect 23572 6817 23581 6851
rect 23581 6817 23615 6851
rect 23615 6817 23624 6851
rect 23572 6808 23624 6817
rect 17040 6740 17092 6749
rect 17316 6740 17368 6792
rect 14648 6604 14700 6656
rect 15292 6604 15344 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 15752 6604 15804 6656
rect 15936 6604 15988 6656
rect 16212 6604 16264 6656
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 17408 6604 17460 6656
rect 17868 6740 17920 6792
rect 18512 6740 18564 6792
rect 19340 6740 19392 6792
rect 19984 6783 20036 6792
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 21548 6740 21600 6792
rect 19156 6672 19208 6724
rect 17776 6604 17828 6656
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 19064 6604 19116 6656
rect 19248 6604 19300 6656
rect 21364 6672 21416 6724
rect 24216 6783 24268 6792
rect 24216 6749 24225 6783
rect 24225 6749 24259 6783
rect 24259 6749 24268 6783
rect 24216 6740 24268 6749
rect 24768 6808 24820 6860
rect 24860 6740 24912 6792
rect 23388 6672 23440 6724
rect 27528 6876 27580 6928
rect 25136 6808 25188 6860
rect 26608 6808 26660 6860
rect 22008 6604 22060 6656
rect 24676 6604 24728 6656
rect 25228 6715 25280 6724
rect 25228 6681 25237 6715
rect 25237 6681 25271 6715
rect 25271 6681 25280 6715
rect 25228 6672 25280 6681
rect 25412 6672 25464 6724
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 27896 6740 27948 6792
rect 27988 6783 28040 6792
rect 27988 6749 27997 6783
rect 27997 6749 28031 6783
rect 28031 6749 28040 6783
rect 27988 6740 28040 6749
rect 26332 6604 26384 6656
rect 27804 6604 27856 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1400 6332 1452 6384
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 6368 6400 6420 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 9220 6400 9272 6452
rect 3792 6264 3844 6316
rect 4988 6264 5040 6316
rect 5448 6264 5500 6316
rect 5264 6196 5316 6248
rect 3884 6128 3936 6180
rect 7104 6264 7156 6316
rect 8208 6196 8260 6248
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 12072 6443 12124 6452
rect 12072 6409 12081 6443
rect 12081 6409 12115 6443
rect 12115 6409 12124 6443
rect 12072 6400 12124 6409
rect 12348 6400 12400 6452
rect 12532 6400 12584 6452
rect 13636 6400 13688 6452
rect 14188 6400 14240 6452
rect 15200 6400 15252 6452
rect 15292 6400 15344 6452
rect 11796 6264 11848 6316
rect 12072 6264 12124 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 14188 6264 14240 6316
rect 8668 6196 8720 6248
rect 9496 6196 9548 6248
rect 9588 6196 9640 6248
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 13084 6196 13136 6248
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13544 6196 13596 6248
rect 18604 6400 18656 6452
rect 19340 6400 19392 6452
rect 22284 6400 22336 6452
rect 2320 6060 2372 6112
rect 2780 6060 2832 6112
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 10784 6128 10836 6180
rect 11060 6128 11112 6180
rect 12440 6128 12492 6180
rect 12808 6128 12860 6180
rect 16764 6332 16816 6384
rect 20260 6332 20312 6384
rect 25228 6400 25280 6452
rect 26608 6400 26660 6452
rect 23020 6332 23072 6384
rect 24400 6332 24452 6384
rect 24492 6332 24544 6384
rect 24952 6332 25004 6384
rect 14648 6060 14700 6112
rect 16028 6128 16080 6180
rect 16212 6103 16264 6112
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 18420 6196 18472 6248
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 19156 6264 19208 6316
rect 19248 6264 19300 6316
rect 19432 6264 19484 6316
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 22652 6307 22704 6316
rect 22652 6273 22661 6307
rect 22661 6273 22695 6307
rect 22695 6273 22704 6307
rect 22652 6264 22704 6273
rect 23940 6264 23992 6316
rect 24032 6264 24084 6316
rect 25780 6332 25832 6384
rect 26056 6332 26108 6384
rect 26240 6332 26292 6384
rect 27896 6400 27948 6452
rect 25136 6196 25188 6248
rect 27804 6196 27856 6248
rect 17684 6060 17736 6112
rect 17960 6060 18012 6112
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 19156 6060 19208 6112
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 24216 6103 24268 6112
rect 24216 6069 24225 6103
rect 24225 6069 24259 6103
rect 24259 6069 24268 6103
rect 24216 6060 24268 6069
rect 25044 6128 25096 6180
rect 25412 6128 25464 6180
rect 27620 6103 27672 6112
rect 27620 6069 27629 6103
rect 27629 6069 27663 6103
rect 27663 6069 27672 6103
rect 27620 6060 27672 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 3792 5856 3844 5908
rect 5816 5856 5868 5908
rect 7472 5856 7524 5908
rect 7564 5856 7616 5908
rect 8576 5856 8628 5908
rect 9588 5899 9640 5908
rect 9588 5865 9597 5899
rect 9597 5865 9631 5899
rect 9631 5865 9640 5899
rect 9588 5856 9640 5865
rect 9956 5856 10008 5908
rect 11060 5856 11112 5908
rect 11704 5856 11756 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13176 5856 13228 5908
rect 13360 5856 13412 5908
rect 15752 5856 15804 5908
rect 16028 5856 16080 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 17224 5856 17276 5908
rect 17868 5856 17920 5908
rect 19248 5856 19300 5908
rect 20904 5899 20956 5908
rect 20904 5865 20913 5899
rect 20913 5865 20947 5899
rect 20947 5865 20956 5899
rect 20904 5856 20956 5865
rect 21364 5856 21416 5908
rect 1400 5652 1452 5704
rect 1860 5652 1912 5704
rect 2320 5695 2372 5704
rect 2320 5661 2354 5695
rect 2354 5661 2372 5695
rect 2320 5652 2372 5661
rect 4160 5652 4212 5704
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 7748 5720 7800 5772
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 6736 5695 6788 5704
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 3056 5516 3108 5568
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 7104 5516 7156 5568
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 7564 5652 7616 5704
rect 8300 5652 8352 5704
rect 11244 5788 11296 5840
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10600 5720 10652 5772
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11980 5652 12032 5704
rect 11520 5584 11572 5636
rect 11796 5584 11848 5636
rect 14372 5720 14424 5772
rect 15292 5720 15344 5772
rect 16580 5788 16632 5840
rect 14372 5584 14424 5636
rect 15200 5584 15252 5636
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 16764 5652 16816 5704
rect 18604 5831 18656 5840
rect 18604 5797 18613 5831
rect 18613 5797 18647 5831
rect 18647 5797 18656 5831
rect 18604 5788 18656 5797
rect 17776 5652 17828 5704
rect 18328 5652 18380 5704
rect 19800 5720 19852 5772
rect 19892 5720 19944 5772
rect 23572 5899 23624 5908
rect 23572 5865 23581 5899
rect 23581 5865 23615 5899
rect 23615 5865 23624 5899
rect 23572 5856 23624 5865
rect 24216 5856 24268 5908
rect 25136 5856 25188 5908
rect 25504 5899 25556 5908
rect 25504 5865 25513 5899
rect 25513 5865 25547 5899
rect 25547 5865 25556 5899
rect 25504 5856 25556 5865
rect 26792 5856 26844 5908
rect 27620 5856 27672 5908
rect 19616 5652 19668 5704
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 10600 5516 10652 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 17684 5516 17736 5568
rect 19984 5584 20036 5636
rect 18236 5516 18288 5568
rect 19156 5516 19208 5568
rect 19340 5516 19392 5568
rect 19800 5516 19852 5568
rect 22836 5720 22888 5772
rect 24308 5788 24360 5840
rect 25780 5720 25832 5772
rect 26424 5763 26476 5772
rect 26424 5729 26433 5763
rect 26433 5729 26467 5763
rect 26467 5729 26476 5763
rect 26424 5720 26476 5729
rect 22928 5652 22980 5704
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 24124 5652 24176 5704
rect 24676 5652 24728 5704
rect 24860 5584 24912 5636
rect 25136 5695 25188 5704
rect 25136 5661 25145 5695
rect 25145 5661 25179 5695
rect 25179 5661 25188 5695
rect 25136 5652 25188 5661
rect 25596 5652 25648 5704
rect 25688 5652 25740 5704
rect 26148 5695 26200 5704
rect 26148 5661 26157 5695
rect 26157 5661 26191 5695
rect 26191 5661 26200 5695
rect 26148 5652 26200 5661
rect 28540 5856 28592 5908
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 27528 5584 27580 5636
rect 28172 5516 28224 5568
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 5080 5312 5132 5364
rect 6736 5312 6788 5364
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 7472 5355 7524 5364
rect 7472 5321 7481 5355
rect 7481 5321 7515 5355
rect 7515 5321 7524 5355
rect 7472 5312 7524 5321
rect 8944 5312 8996 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2136 5176 2188 5228
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3516 5176 3568 5228
rect 3148 5108 3200 5160
rect 5264 5176 5316 5228
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 5908 5219 5960 5228
rect 5908 5185 5925 5219
rect 5925 5185 5959 5219
rect 5959 5185 5960 5219
rect 5908 5176 5960 5185
rect 6276 5176 6328 5228
rect 8300 5244 8352 5296
rect 9496 5312 9548 5364
rect 10232 5312 10284 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 11520 5312 11572 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 16488 5312 16540 5364
rect 16580 5312 16632 5364
rect 12072 5287 12124 5296
rect 7656 5176 7708 5228
rect 5080 5108 5132 5160
rect 6644 5151 6696 5160
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 7748 5108 7800 5160
rect 6552 5040 6604 5092
rect 12072 5253 12081 5287
rect 12081 5253 12115 5287
rect 12115 5253 12124 5287
rect 12072 5244 12124 5253
rect 13084 5244 13136 5296
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 8300 4972 8352 5024
rect 8392 4972 8444 5024
rect 8668 4972 8720 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 11796 5176 11848 5228
rect 14556 5244 14608 5296
rect 10048 5108 10100 5160
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 12532 5108 12584 5160
rect 10692 5040 10744 5092
rect 13544 5108 13596 5160
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 14280 5108 14332 5160
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 17316 5312 17368 5364
rect 18236 5312 18288 5364
rect 18604 5312 18656 5364
rect 20628 5312 20680 5364
rect 20812 5312 20864 5364
rect 23204 5312 23256 5364
rect 23848 5312 23900 5364
rect 23940 5312 23992 5364
rect 25136 5312 25188 5364
rect 25504 5312 25556 5364
rect 16948 5108 17000 5160
rect 17316 5176 17368 5228
rect 17592 5108 17644 5160
rect 17868 5108 17920 5160
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18788 5244 18840 5296
rect 19340 5244 19392 5296
rect 19524 5244 19576 5296
rect 19892 5287 19944 5296
rect 19892 5253 19901 5287
rect 19901 5253 19935 5287
rect 19935 5253 19944 5287
rect 19892 5244 19944 5253
rect 20444 5244 20496 5296
rect 25044 5244 25096 5296
rect 19248 5176 19300 5228
rect 20720 5176 20772 5228
rect 15384 4972 15436 5024
rect 21088 5108 21140 5160
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 21640 5176 21692 5228
rect 21916 5176 21968 5228
rect 22652 5176 22704 5228
rect 17684 5015 17736 5024
rect 17684 4981 17693 5015
rect 17693 4981 17727 5015
rect 17727 4981 17736 5015
rect 17684 4972 17736 4981
rect 18052 4972 18104 5024
rect 20352 5083 20404 5092
rect 20352 5049 20361 5083
rect 20361 5049 20395 5083
rect 20395 5049 20404 5083
rect 20352 5040 20404 5049
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 22100 5040 22152 5092
rect 22192 5083 22244 5092
rect 22192 5049 22201 5083
rect 22201 5049 22235 5083
rect 22235 5049 22244 5083
rect 22192 5040 22244 5049
rect 22376 5040 22428 5092
rect 23664 4972 23716 5024
rect 23756 4972 23808 5024
rect 24216 4972 24268 5024
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 24768 5176 24820 5228
rect 26700 5312 26752 5364
rect 28540 5355 28592 5364
rect 28540 5321 28549 5355
rect 28549 5321 28583 5355
rect 28583 5321 28592 5355
rect 28540 5312 28592 5321
rect 26884 5244 26936 5296
rect 27528 5244 27580 5296
rect 26240 5176 26292 5228
rect 26424 5176 26476 5228
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 25320 5151 25372 5160
rect 25320 5117 25329 5151
rect 25329 5117 25363 5151
rect 25363 5117 25372 5151
rect 25320 5108 25372 5117
rect 25780 5040 25832 5092
rect 24952 4972 25004 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 5264 4768 5316 4820
rect 6644 4768 6696 4820
rect 7564 4768 7616 4820
rect 8392 4768 8444 4820
rect 8484 4811 8536 4820
rect 8484 4777 8493 4811
rect 8493 4777 8527 4811
rect 8527 4777 8536 4811
rect 8484 4768 8536 4777
rect 1400 4632 1452 4684
rect 2136 4632 2188 4684
rect 1952 4564 2004 4616
rect 2320 4564 2372 4616
rect 4712 4564 4764 4616
rect 5080 4564 5132 4616
rect 5908 4700 5960 4752
rect 6920 4700 6972 4752
rect 4252 4496 4304 4548
rect 7012 4632 7064 4684
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 5816 4428 5868 4480
rect 12808 4768 12860 4820
rect 13452 4768 13504 4820
rect 13636 4768 13688 4820
rect 14372 4768 14424 4820
rect 15752 4768 15804 4820
rect 16028 4768 16080 4820
rect 16948 4768 17000 4820
rect 17132 4768 17184 4820
rect 17960 4768 18012 4820
rect 19340 4768 19392 4820
rect 20720 4768 20772 4820
rect 22100 4768 22152 4820
rect 22376 4768 22428 4820
rect 8760 4632 8812 4684
rect 8576 4564 8628 4616
rect 10232 4632 10284 4684
rect 11244 4632 11296 4684
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 13084 4700 13136 4752
rect 13728 4700 13780 4752
rect 8668 4428 8720 4480
rect 11336 4496 11388 4548
rect 12808 4496 12860 4548
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 11796 4428 11848 4480
rect 13452 4496 13504 4548
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 16212 4632 16264 4684
rect 18144 4632 18196 4684
rect 16580 4564 16632 4616
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 14096 4428 14148 4480
rect 18052 4496 18104 4548
rect 18144 4496 18196 4548
rect 18420 4539 18472 4548
rect 18420 4505 18429 4539
rect 18429 4505 18463 4539
rect 18463 4505 18472 4539
rect 18420 4496 18472 4505
rect 18788 4496 18840 4548
rect 21088 4700 21140 4752
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 20628 4564 20680 4616
rect 20260 4496 20312 4548
rect 24308 4768 24360 4820
rect 25136 4768 25188 4820
rect 25780 4811 25832 4820
rect 25780 4777 25789 4811
rect 25789 4777 25823 4811
rect 25823 4777 25832 4811
rect 25780 4768 25832 4777
rect 27804 4768 27856 4820
rect 23664 4743 23716 4752
rect 23664 4709 23673 4743
rect 23673 4709 23707 4743
rect 23707 4709 23716 4743
rect 23664 4700 23716 4709
rect 23848 4700 23900 4752
rect 24584 4700 24636 4752
rect 23756 4632 23808 4684
rect 23204 4564 23256 4616
rect 27068 4632 27120 4684
rect 27252 4632 27304 4684
rect 27620 4632 27672 4684
rect 23572 4496 23624 4548
rect 24400 4607 24452 4616
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 23296 4428 23348 4480
rect 24308 4496 24360 4548
rect 24860 4564 24912 4616
rect 24952 4564 25004 4616
rect 25504 4564 25556 4616
rect 26148 4607 26200 4616
rect 26148 4573 26157 4607
rect 26157 4573 26191 4607
rect 26191 4573 26200 4607
rect 26148 4564 26200 4573
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 26792 4564 26844 4616
rect 27620 4496 27672 4548
rect 25412 4428 25464 4480
rect 26240 4428 26292 4480
rect 26792 4428 26844 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 4712 4224 4764 4276
rect 5448 4267 5500 4276
rect 5448 4233 5457 4267
rect 5457 4233 5491 4267
rect 5491 4233 5500 4267
rect 5448 4224 5500 4233
rect 5816 4224 5868 4276
rect 6920 4224 6972 4276
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 3240 4088 3292 4140
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 4344 4020 4396 4029
rect 4988 4088 5040 4140
rect 5448 4088 5500 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6736 4156 6788 4208
rect 13084 4224 13136 4276
rect 13360 4224 13412 4276
rect 16212 4267 16264 4276
rect 16212 4233 16221 4267
rect 16221 4233 16255 4267
rect 16255 4233 16264 4267
rect 16212 4224 16264 4233
rect 19708 4224 19760 4276
rect 8116 4135 8168 4140
rect 8116 4101 8125 4135
rect 8125 4101 8159 4135
rect 8159 4101 8168 4135
rect 8116 4088 8168 4101
rect 8300 4088 8352 4140
rect 5356 4020 5408 4072
rect 4804 3995 4856 4004
rect 4804 3961 4813 3995
rect 4813 3961 4847 3995
rect 4847 3961 4856 3995
rect 4804 3952 4856 3961
rect 6644 4020 6696 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 7012 3952 7064 4004
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 10140 4088 10192 4140
rect 11244 4088 11296 4140
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 13544 4156 13596 4208
rect 10508 4020 10560 4072
rect 13728 4020 13780 4072
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 15292 4088 15344 4140
rect 17960 4199 18012 4208
rect 17960 4165 17969 4199
rect 17969 4165 18003 4199
rect 18003 4165 18012 4199
rect 17960 4156 18012 4165
rect 19156 4156 19208 4208
rect 16120 4131 16172 4140
rect 13820 4020 13872 4029
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 18052 4020 18104 4072
rect 19524 4088 19576 4140
rect 20260 4156 20312 4208
rect 21180 4156 21232 4208
rect 21456 4224 21508 4276
rect 24308 4224 24360 4276
rect 24400 4224 24452 4276
rect 24768 4267 24820 4276
rect 24768 4233 24777 4267
rect 24777 4233 24811 4267
rect 24811 4233 24820 4267
rect 24768 4224 24820 4233
rect 27620 4224 27672 4276
rect 25504 4156 25556 4208
rect 4252 3884 4304 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6460 3884 6512 3936
rect 19248 4063 19300 4072
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 19984 4088 20036 4140
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 9864 3884 9916 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 12532 3884 12584 3936
rect 15660 3884 15712 3936
rect 19340 3952 19392 4004
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 17408 3884 17460 3936
rect 18512 3884 18564 3936
rect 20628 3884 20680 3936
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 21456 3884 21508 3936
rect 23388 4088 23440 4140
rect 25136 4088 25188 4140
rect 25412 4088 25464 4140
rect 25688 4088 25740 4140
rect 26792 4088 26844 4140
rect 26976 4088 27028 4140
rect 27712 4088 27764 4140
rect 23664 4020 23716 4072
rect 24032 4063 24084 4072
rect 24032 4029 24041 4063
rect 24041 4029 24075 4063
rect 24075 4029 24084 4063
rect 24032 4020 24084 4029
rect 24216 4063 24268 4072
rect 24216 4029 24225 4063
rect 24225 4029 24259 4063
rect 24259 4029 24268 4063
rect 24216 4020 24268 4029
rect 24860 4020 24912 4072
rect 25780 4020 25832 4072
rect 26148 4020 26200 4072
rect 26332 4020 26384 4072
rect 26516 4020 26568 4072
rect 22744 3884 22796 3936
rect 23204 3927 23256 3936
rect 23204 3893 23213 3927
rect 23213 3893 23247 3927
rect 23247 3893 23256 3927
rect 23204 3884 23256 3893
rect 23388 3884 23440 3936
rect 25136 3884 25188 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 3148 3680 3200 3732
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 4344 3680 4396 3732
rect 5356 3680 5408 3732
rect 7288 3680 7340 3732
rect 8208 3680 8260 3732
rect 9312 3680 9364 3732
rect 9680 3680 9732 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 4712 3612 4764 3664
rect 5172 3612 5224 3664
rect 5632 3612 5684 3664
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 1676 3476 1728 3528
rect 1860 3476 1912 3528
rect 1952 3476 2004 3528
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 6644 3544 6696 3596
rect 6736 3544 6788 3596
rect 12440 3680 12492 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 13820 3680 13872 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 11704 3544 11756 3596
rect 14004 3612 14056 3664
rect 16764 3680 16816 3732
rect 17224 3680 17276 3732
rect 19616 3680 19668 3732
rect 21364 3680 21416 3732
rect 21456 3680 21508 3732
rect 3240 3476 3292 3528
rect 3424 3521 3476 3528
rect 3424 3487 3433 3521
rect 3433 3487 3467 3521
rect 3467 3487 3476 3521
rect 3424 3476 3476 3487
rect 3608 3476 3660 3528
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4252 3476 4304 3528
rect 3148 3408 3200 3460
rect 5172 3451 5224 3460
rect 5172 3417 5181 3451
rect 5181 3417 5215 3451
rect 5215 3417 5224 3451
rect 5172 3408 5224 3417
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5724 3476 5776 3528
rect 6276 3476 6328 3528
rect 6000 3408 6052 3460
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 6644 3451 6696 3460
rect 6644 3417 6653 3451
rect 6653 3417 6687 3451
rect 6687 3417 6696 3451
rect 6644 3408 6696 3417
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 3424 3340 3476 3392
rect 8668 3476 8720 3528
rect 9680 3408 9732 3460
rect 10048 3476 10100 3528
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 10324 3408 10376 3460
rect 11152 3408 11204 3460
rect 13084 3476 13136 3528
rect 14188 3476 14240 3528
rect 16672 3612 16724 3664
rect 18696 3612 18748 3664
rect 20628 3612 20680 3664
rect 13544 3408 13596 3460
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 16856 3476 16908 3528
rect 19432 3544 19484 3596
rect 19524 3544 19576 3596
rect 20260 3544 20312 3596
rect 24308 3680 24360 3732
rect 24400 3680 24452 3732
rect 25872 3680 25924 3732
rect 26148 3680 26200 3732
rect 26608 3723 26660 3732
rect 26608 3689 26617 3723
rect 26617 3689 26651 3723
rect 26651 3689 26660 3723
rect 26608 3680 26660 3689
rect 26792 3680 26844 3732
rect 23664 3612 23716 3664
rect 16764 3408 16816 3460
rect 17868 3408 17920 3460
rect 18972 3476 19024 3528
rect 23388 3587 23440 3596
rect 23388 3553 23397 3587
rect 23397 3553 23431 3587
rect 23431 3553 23440 3587
rect 23388 3544 23440 3553
rect 23940 3612 23992 3664
rect 25688 3612 25740 3664
rect 23848 3544 23900 3596
rect 25872 3587 25924 3596
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 26056 3587 26108 3596
rect 26056 3553 26065 3587
rect 26065 3553 26099 3587
rect 26099 3553 26108 3587
rect 26056 3544 26108 3553
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 16580 3383 16632 3392
rect 16580 3349 16589 3383
rect 16589 3349 16623 3383
rect 16623 3349 16632 3383
rect 16580 3340 16632 3349
rect 18236 3340 18288 3392
rect 19156 3408 19208 3460
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 24492 3476 24544 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 27344 3680 27396 3732
rect 27160 3587 27212 3596
rect 27160 3553 27169 3587
rect 27169 3553 27203 3587
rect 27203 3553 27212 3587
rect 27160 3544 27212 3553
rect 20444 3408 20496 3460
rect 24676 3408 24728 3460
rect 27988 3408 28040 3460
rect 19340 3340 19392 3392
rect 20352 3340 20404 3392
rect 21272 3340 21324 3392
rect 25688 3340 25740 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 3240 3136 3292 3188
rect 3332 3136 3384 3188
rect 5264 3136 5316 3188
rect 6460 3179 6512 3188
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 7748 3136 7800 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 2136 3068 2188 3120
rect 4068 3000 4120 3052
rect 4528 3000 4580 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 8576 3136 8628 3188
rect 8668 3136 8720 3188
rect 11428 3136 11480 3188
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8208 3068 8260 3120
rect 6828 2932 6880 2984
rect 2504 2796 2556 2848
rect 4344 2907 4396 2916
rect 4344 2873 4353 2907
rect 4353 2873 4387 2907
rect 4387 2873 4396 2907
rect 4344 2864 4396 2873
rect 4160 2796 4212 2848
rect 5448 2796 5500 2848
rect 10600 3000 10652 3052
rect 11244 3000 11296 3052
rect 14004 3136 14056 3188
rect 14188 3136 14240 3188
rect 14924 3136 14976 3188
rect 16120 3136 16172 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 17776 3136 17828 3188
rect 18052 3136 18104 3188
rect 18696 3136 18748 3188
rect 18788 3136 18840 3188
rect 12348 3068 12400 3120
rect 16764 3068 16816 3120
rect 16580 3000 16632 3052
rect 19156 3068 19208 3120
rect 19432 3068 19484 3120
rect 20168 3068 20220 3120
rect 20444 3136 20496 3188
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 17592 2932 17644 2984
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 21272 3000 21324 3052
rect 22652 3136 22704 3188
rect 23756 3179 23808 3188
rect 23756 3145 23765 3179
rect 23765 3145 23799 3179
rect 23799 3145 23808 3179
rect 23756 3136 23808 3145
rect 23848 3136 23900 3188
rect 24860 3136 24912 3188
rect 27160 3136 27212 3188
rect 19800 2932 19852 2984
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 19984 2864 20036 2916
rect 20996 2864 21048 2916
rect 15292 2796 15344 2848
rect 18144 2796 18196 2848
rect 18696 2796 18748 2848
rect 20904 2796 20956 2848
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 25136 3000 25188 3052
rect 23296 2907 23348 2916
rect 23296 2873 23305 2907
rect 23305 2873 23339 2907
rect 23339 2873 23348 2907
rect 23296 2864 23348 2873
rect 23388 2839 23440 2848
rect 23388 2805 23397 2839
rect 23397 2805 23431 2839
rect 23431 2805 23440 2839
rect 23388 2796 23440 2805
rect 24676 2796 24728 2848
rect 26700 3000 26752 3052
rect 27252 3043 27304 3052
rect 27252 3009 27286 3043
rect 27286 3009 27304 3043
rect 27252 3000 27304 3009
rect 27160 2796 27212 2848
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 2136 2592 2188 2644
rect 2504 2592 2556 2644
rect 2044 2524 2096 2576
rect 3240 2592 3292 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 10048 2592 10100 2644
rect 10324 2592 10376 2644
rect 10876 2592 10928 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 3516 2456 3568 2508
rect 1400 2388 1452 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 3240 2388 3292 2440
rect 3424 2388 3476 2440
rect 4160 2456 4212 2508
rect 5816 2456 5868 2508
rect 10416 2524 10468 2576
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 14464 2592 14516 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 15292 2592 15344 2644
rect 16948 2592 17000 2644
rect 19892 2592 19944 2644
rect 19984 2592 20036 2644
rect 24584 2592 24636 2644
rect 13084 2524 13136 2533
rect 8208 2456 8260 2508
rect 11244 2456 11296 2508
rect 6276 2388 6328 2440
rect 3148 2252 3200 2304
rect 8024 2320 8076 2372
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 10508 2388 10560 2440
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 13176 2252 13228 2304
rect 13636 2252 13688 2304
rect 14924 2388 14976 2440
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 17868 2524 17920 2576
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 17960 2456 18012 2508
rect 16764 2388 16816 2440
rect 17684 2388 17736 2440
rect 17776 2388 17828 2440
rect 18236 2320 18288 2372
rect 19524 2388 19576 2440
rect 21548 2524 21600 2576
rect 20352 2456 20404 2508
rect 20628 2499 20680 2508
rect 20628 2465 20637 2499
rect 20637 2465 20671 2499
rect 20671 2465 20680 2499
rect 20628 2456 20680 2465
rect 21088 2499 21140 2508
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 20812 2431 20864 2440
rect 20812 2397 20821 2431
rect 20821 2397 20855 2431
rect 20855 2397 20864 2431
rect 20812 2388 20864 2397
rect 21916 2499 21968 2508
rect 21916 2465 21925 2499
rect 21925 2465 21959 2499
rect 21959 2465 21968 2499
rect 21916 2456 21968 2465
rect 23572 2524 23624 2576
rect 24768 2567 24820 2576
rect 24768 2533 24777 2567
rect 24777 2533 24811 2567
rect 24811 2533 24820 2567
rect 24768 2524 24820 2533
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 23112 2456 23164 2508
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 23848 2431 23900 2440
rect 23848 2397 23857 2431
rect 23857 2397 23891 2431
rect 23891 2397 23900 2431
rect 23848 2388 23900 2397
rect 24952 2431 25004 2440
rect 24952 2397 24961 2431
rect 24961 2397 24995 2431
rect 24995 2397 25004 2431
rect 24952 2388 25004 2397
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 21548 2320 21600 2372
rect 23388 2320 23440 2372
rect 24768 2320 24820 2372
rect 25596 2592 25648 2644
rect 26056 2592 26108 2644
rect 26700 2592 26752 2644
rect 27252 2592 27304 2644
rect 27988 2592 28040 2644
rect 25688 2456 25740 2508
rect 27068 2499 27120 2508
rect 27068 2465 27077 2499
rect 27077 2465 27111 2499
rect 27111 2465 27120 2499
rect 27068 2456 27120 2465
rect 28540 2456 28592 2508
rect 28356 2388 28408 2440
rect 23480 2295 23532 2304
rect 23480 2261 23489 2295
rect 23489 2261 23523 2295
rect 23523 2261 23532 2295
rect 23480 2252 23532 2261
rect 23572 2295 23624 2304
rect 23572 2261 23581 2295
rect 23581 2261 23615 2295
rect 23615 2261 23624 2295
rect 23572 2252 23624 2261
rect 23664 2252 23716 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 2044 2048 2096 2100
rect 2136 2048 2188 2100
rect 23388 2048 23440 2100
rect 23480 2048 23532 2100
rect 23572 2048 23624 2100
rect 4804 1980 4856 2032
rect 10416 1980 10468 2032
rect 11336 1980 11388 2032
rect 11612 1980 11664 2032
rect 13636 1980 13688 2032
rect 15476 1980 15528 2032
rect 19800 1980 19852 2032
rect 17500 1912 17552 1964
rect 21548 1912 21600 1964
rect 9864 1776 9916 1828
rect 13084 1776 13136 1828
rect 16764 1776 16816 1828
rect 23204 1912 23256 1964
rect 18788 1708 18840 1760
rect 24216 1640 24268 1692
<< metal2 >>
rect 3790 29200 3846 30000
rect 11242 29200 11298 30000
rect 18694 29200 18750 30000
rect 26146 29200 26202 30000
rect 3804 27606 3832 29200
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 9692 27606 9720 27814
rect 3792 27600 3844 27606
rect 3792 27542 3844 27548
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 11256 27554 11284 29200
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 1492 27396 1544 27402
rect 1492 27338 1544 27344
rect 940 27328 992 27334
rect 938 27296 940 27305
rect 992 27296 994 27305
rect 938 27231 994 27240
rect 1504 27130 1532 27338
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4632 27130 4660 27270
rect 1492 27124 1544 27130
rect 1492 27066 1544 27072
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 2596 27056 2648 27062
rect 2594 27024 2596 27033
rect 2688 27056 2740 27062
rect 2648 27024 2650 27033
rect 2320 26988 2372 26994
rect 2688 26998 2740 27004
rect 2594 26959 2650 26968
rect 2320 26930 2372 26936
rect 2228 26784 2280 26790
rect 2228 26726 2280 26732
rect 2240 26586 2268 26726
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2332 26042 2360 26930
rect 2700 26586 2728 26998
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3516 26920 3568 26926
rect 3804 26897 3832 26930
rect 3516 26862 3568 26868
rect 3790 26888 3846 26897
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 2688 26580 2740 26586
rect 2688 26522 2740 26528
rect 3252 26246 3280 26726
rect 3528 26586 3556 26862
rect 3790 26823 3846 26832
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 4816 26382 4844 27270
rect 4908 27130 4936 27270
rect 4896 27124 4948 27130
rect 4896 27066 4948 27072
rect 5092 26586 5120 27406
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 5080 26580 5132 26586
rect 5080 26522 5132 26528
rect 5276 26450 5304 26794
rect 5264 26444 5316 26450
rect 5264 26386 5316 26392
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 3240 26240 3292 26246
rect 3240 26182 3292 26188
rect 4344 26240 4396 26246
rect 4344 26182 4396 26188
rect 4896 26240 4948 26246
rect 4896 26182 4948 26188
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1400 25696 1452 25702
rect 1400 25638 1452 25644
rect 1412 25498 1440 25638
rect 1400 25492 1452 25498
rect 1400 25434 1452 25440
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23118 1440 24142
rect 1596 23769 1624 25842
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2044 25696 2096 25702
rect 2044 25638 2096 25644
rect 2056 25498 2084 25638
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 2516 25430 2544 25774
rect 3252 25702 3280 26182
rect 3424 25832 3476 25838
rect 3422 25800 3424 25809
rect 3608 25832 3660 25838
rect 3476 25800 3478 25809
rect 3608 25774 3660 25780
rect 3422 25735 3478 25744
rect 3240 25696 3292 25702
rect 3292 25644 3372 25650
rect 3240 25638 3372 25644
rect 3252 25622 3372 25638
rect 2504 25424 2556 25430
rect 2504 25366 2556 25372
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1582 23760 1638 23769
rect 1582 23695 1638 23704
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22098 1440 23054
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1412 21010 1440 22034
rect 1688 21554 1716 25230
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1964 24993 1992 25094
rect 1950 24984 2006 24993
rect 1950 24919 2006 24928
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 1780 24410 1808 24550
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 2056 21554 2084 25094
rect 2516 24818 2544 25366
rect 2596 25288 2648 25294
rect 2596 25230 2648 25236
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2136 24132 2188 24138
rect 2136 24074 2188 24080
rect 2148 23866 2176 24074
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2240 23118 2268 23666
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2516 22642 2544 24754
rect 2608 23526 2636 25230
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2792 24886 2820 25094
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2608 23322 2636 23462
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2792 23186 2820 24550
rect 2884 24410 2912 25230
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2976 24274 3004 25094
rect 3068 24818 3096 25162
rect 3344 25158 3372 25622
rect 3620 25498 3648 25774
rect 3976 25764 4028 25770
rect 3976 25706 4028 25712
rect 3988 25498 4016 25706
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3884 25356 3936 25362
rect 3884 25298 3936 25304
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 3056 24676 3108 24682
rect 3056 24618 3108 24624
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2516 22522 2544 22578
rect 2424 22506 2544 22522
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2412 22500 2544 22506
rect 2464 22494 2544 22500
rect 2412 22442 2464 22448
rect 2516 22166 2544 22494
rect 2700 22234 2728 22510
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2504 22160 2556 22166
rect 2504 22102 2556 22108
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 2240 21690 2268 21898
rect 2700 21690 2728 22170
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2792 21554 2820 22374
rect 2976 21554 3004 22578
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 1688 21146 1716 21490
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 3068 20890 3096 24618
rect 3252 24274 3280 25094
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3344 24154 3372 25094
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3712 24342 3740 24550
rect 3700 24336 3752 24342
rect 3700 24278 3752 24284
rect 3252 24126 3372 24154
rect 3252 23662 3280 24126
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3528 23730 3556 24006
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3252 23474 3280 23598
rect 3160 23446 3280 23474
rect 3160 22030 3188 23446
rect 3332 23044 3384 23050
rect 3332 22986 3384 22992
rect 3344 22778 3372 22986
rect 3332 22772 3384 22778
rect 3332 22714 3384 22720
rect 3240 22704 3292 22710
rect 3240 22646 3292 22652
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2976 20862 3096 20890
rect 2608 20602 2636 20810
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2780 20392 2832 20398
rect 2976 20369 3004 20862
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2780 20334 2832 20340
rect 2962 20360 3018 20369
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19378 1440 19790
rect 1504 19514 1532 20198
rect 2056 20058 2084 20334
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2792 19514 2820 20334
rect 2962 20295 3018 20304
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2976 19854 3004 20198
rect 3068 19854 3096 20742
rect 3252 20466 3280 22646
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 3620 22234 3648 22578
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3332 22160 3384 22166
rect 3384 22120 3556 22148
rect 3332 22102 3384 22108
rect 3528 22094 3556 22120
rect 3712 22098 3740 24278
rect 3804 23866 3832 24754
rect 3896 24750 3924 25298
rect 4356 25294 4384 26182
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4908 25294 4936 26182
rect 5184 25906 5212 26182
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 4896 25288 4948 25294
rect 4896 25230 4948 25236
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 3896 23798 3924 24686
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3884 23792 3936 23798
rect 3884 23734 3936 23740
rect 3896 23118 3924 23734
rect 3988 23322 4016 24550
rect 4264 24206 4292 25094
rect 4540 24954 4568 25094
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 4816 24614 4844 25230
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4908 24274 4936 25230
rect 5184 24614 5212 25842
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 4896 24268 4948 24274
rect 4896 24210 4948 24216
rect 5184 24206 5212 24550
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4252 23520 4304 23526
rect 4252 23462 4304 23468
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 4264 23050 4292 23462
rect 4252 23044 4304 23050
rect 4252 22986 4304 22992
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4172 22778 4200 22918
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 3528 22066 3648 22094
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3436 20942 3464 21966
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3344 20602 3372 20810
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3620 20534 3648 22066
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3712 20942 3740 21286
rect 3896 21146 3924 21422
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 4080 20942 4108 21830
rect 4172 21554 4200 22714
rect 4356 22642 4384 23530
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4816 22094 4844 24006
rect 4908 23866 4936 24006
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 5000 23322 5028 23666
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4896 23248 4948 23254
rect 4896 23190 4948 23196
rect 4908 22574 4936 23190
rect 5000 22574 5028 23258
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4816 22066 5028 22094
rect 4344 22024 4396 22030
rect 4344 21966 4396 21972
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4356 21146 4384 21966
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4632 21690 4660 21830
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4724 21622 4752 21830
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 19854 3372 20198
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 19514 3556 19654
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 1412 18290 1440 19314
rect 2240 18970 2268 19314
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2332 18426 2360 18634
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2516 18426 2544 18566
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17746 1440 18226
rect 2792 17882 2820 18702
rect 2884 18426 2912 18770
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3160 17882 3188 18158
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 1320 16697 1348 17138
rect 1306 16688 1362 16697
rect 1412 16658 1440 17682
rect 2320 17604 2372 17610
rect 2320 17546 2372 17552
rect 2332 17338 2360 17546
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 2884 16794 2912 17070
rect 3252 16794 3280 17070
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 1306 16623 1362 16632
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16114 1440 16594
rect 3528 16590 3556 19314
rect 3620 19258 3648 20470
rect 3896 20466 3924 20742
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3712 19378 3740 20402
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19514 3832 20198
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3620 19230 3740 19258
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 17678 3648 19110
rect 3712 18290 3740 19230
rect 3896 18306 3924 20402
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3988 19514 4016 19790
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4172 19378 4200 20198
rect 4264 20058 4292 20742
rect 4816 20466 4844 21626
rect 4908 21554 4936 21966
rect 5000 21554 5028 22066
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 5092 21146 5120 24006
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5184 22642 5212 23462
rect 5368 23050 5396 27474
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6826 27432 6882 27441
rect 6276 27396 6328 27402
rect 6276 27338 6328 27344
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 5460 27130 5488 27270
rect 5736 27130 5764 27270
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 6012 26994 6040 27270
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 5908 26852 5960 26858
rect 5908 26794 5960 26800
rect 5920 26042 5948 26794
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5368 22234 5396 22986
rect 5460 22778 5488 23598
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5262 22128 5318 22137
rect 5262 22063 5264 22072
rect 5316 22063 5318 22072
rect 5264 22034 5316 22040
rect 5552 22030 5580 24686
rect 5736 24410 5764 24686
rect 5828 24410 5856 24754
rect 5724 24404 5776 24410
rect 5724 24346 5776 24352
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 6012 23662 6040 26930
rect 6288 26926 6316 27338
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6656 27062 6684 27270
rect 6748 27130 6776 27406
rect 6826 27367 6882 27376
rect 6840 27334 6868 27367
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6644 27056 6696 27062
rect 6644 26998 6696 27004
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6196 26450 6224 26726
rect 6184 26444 6236 26450
rect 6184 26386 6236 26392
rect 6196 25974 6224 26386
rect 6380 26353 6408 26862
rect 6932 26790 6960 27270
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 8312 27130 8340 27270
rect 8404 27130 8432 27270
rect 8300 27124 8352 27130
rect 8300 27066 8352 27072
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 7012 27056 7064 27062
rect 7012 26998 7064 27004
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6736 26512 6788 26518
rect 6736 26454 6788 26460
rect 6366 26344 6422 26353
rect 6366 26279 6422 26288
rect 6380 26042 6408 26279
rect 6368 26036 6420 26042
rect 6368 25978 6420 25984
rect 6184 25968 6236 25974
rect 6184 25910 6236 25916
rect 6552 25968 6604 25974
rect 6552 25910 6604 25916
rect 6460 25832 6512 25838
rect 6460 25774 6512 25780
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6104 25226 6132 25638
rect 6472 25430 6500 25774
rect 6564 25498 6592 25910
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6460 25424 6512 25430
rect 6460 25366 6512 25372
rect 6748 25294 6776 26454
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6092 25220 6144 25226
rect 6092 25162 6144 25168
rect 6366 24984 6422 24993
rect 6366 24919 6422 24928
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6104 23866 6132 24550
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 6288 23866 6316 24074
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5184 21672 5212 21966
rect 5552 21690 5580 21966
rect 5540 21684 5592 21690
rect 5184 21644 5488 21672
rect 5460 21570 5488 21644
rect 5540 21626 5592 21632
rect 5644 21570 5672 22442
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5828 21894 5856 22374
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5356 21548 5408 21554
rect 5460 21542 5672 21570
rect 5736 21554 5764 21830
rect 5724 21548 5776 21554
rect 5356 21490 5408 21496
rect 5724 21490 5776 21496
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5092 20534 5120 20878
rect 5080 20528 5132 20534
rect 5080 20470 5132 20476
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4356 20058 4384 20402
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4264 19378 4292 19994
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4724 19854 4752 19926
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4816 19378 4844 20198
rect 4908 19786 4936 20198
rect 5000 19990 5028 20334
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4908 19514 4936 19722
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 3988 18426 4016 18702
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4448 18426 4476 18566
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4436 18420 4488 18426
rect 4436 18362 4488 18368
rect 4804 18352 4856 18358
rect 3700 18284 3752 18290
rect 3896 18278 4016 18306
rect 4804 18294 4856 18300
rect 3700 18226 3752 18232
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3712 17338 3740 18226
rect 3988 18154 4016 18278
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3988 17678 4016 18090
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4816 17882 4844 18294
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3344 16250 3372 16526
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16250 3464 16390
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3528 16130 3556 16526
rect 3712 16182 3740 17274
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 3436 16102 3556 16130
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 2240 15706 2268 16050
rect 3436 16046 3464 16102
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 2240 15162 2268 15438
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 13870 1440 14894
rect 2240 14414 2268 15098
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2332 14346 2360 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2976 15094 3004 15302
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14618 2912 14894
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 952 13161 980 13194
rect 938 13152 994 13161
rect 938 13087 994 13096
rect 1412 12782 1440 13806
rect 2056 13326 2084 14214
rect 2332 14074 2360 14282
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13530 2820 13874
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2884 13530 2912 13806
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 13410 3004 14486
rect 3068 14482 3096 15302
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3160 14618 3188 14758
rect 3344 14618 3372 15438
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3436 14414 3464 15982
rect 3712 15570 3740 16118
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3252 13734 3280 14350
rect 3712 14074 3740 15506
rect 3988 15366 4016 17614
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 15978 4200 17070
rect 4264 17066 4292 17614
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4356 16794 4384 17138
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4816 15910 4844 17070
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3988 15094 4016 15302
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 4080 15026 4108 15302
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4172 14482 4200 15574
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4252 15360 4304 15366
rect 4540 15337 4568 15438
rect 4252 15302 4304 15308
rect 4526 15328 4582 15337
rect 4264 15162 4292 15302
rect 4526 15263 4582 15272
rect 4724 15162 4752 15438
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4816 15026 4844 15846
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4356 14618 4384 14758
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 14074 4108 14282
rect 4816 14074 4844 14962
rect 4908 14822 4936 18702
rect 5000 18290 5028 19926
rect 5092 19922 5120 20470
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5184 18358 5212 18770
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15706 5212 15846
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 5276 14498 5304 21422
rect 5368 17218 5396 21490
rect 5540 21480 5592 21486
rect 5538 21448 5540 21457
rect 5592 21448 5594 21457
rect 5538 21383 5594 21392
rect 5920 20942 5948 22374
rect 6012 22166 6040 22578
rect 6196 22234 6224 22714
rect 6380 22642 6408 24919
rect 6552 24744 6604 24750
rect 6552 24686 6604 24692
rect 6564 24410 6592 24686
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6564 23866 6592 24346
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6656 22778 6684 24346
rect 6840 24274 6868 26522
rect 6932 26450 6960 26726
rect 7024 26450 7052 26998
rect 8208 26988 8260 26994
rect 8260 26948 8340 26976
rect 8208 26930 8260 26936
rect 8208 26852 8260 26858
rect 8208 26794 8260 26800
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 8220 26382 8248 26794
rect 8312 26466 8340 26948
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8404 26586 8432 26726
rect 8496 26586 8524 27542
rect 11256 27538 11468 27554
rect 8944 27532 8996 27538
rect 11256 27532 11480 27538
rect 11256 27526 11428 27532
rect 8944 27474 8996 27480
rect 11428 27474 11480 27480
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8588 26466 8616 27270
rect 8312 26438 8708 26466
rect 7288 26376 7340 26382
rect 7286 26344 7288 26353
rect 7656 26376 7708 26382
rect 7340 26344 7342 26353
rect 7932 26376 7984 26382
rect 7656 26318 7708 26324
rect 7760 26336 7932 26364
rect 7286 26279 7342 26288
rect 7288 26036 7340 26042
rect 7288 25978 7340 25984
rect 7012 25764 7064 25770
rect 7012 25706 7064 25712
rect 7024 24682 7052 25706
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7012 24676 7064 24682
rect 7012 24618 7064 24624
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6932 23594 6960 24142
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 6000 22024 6052 22030
rect 5998 21992 6000 22001
rect 6052 21992 6054 22001
rect 5998 21927 6054 21936
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21554 6592 21830
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6472 21146 6500 21354
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 6472 20466 6500 21082
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5460 19514 5488 19926
rect 5644 19514 5672 20198
rect 6104 19786 6132 20198
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 6012 19378 6040 19722
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 5460 18766 5488 19110
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5736 18426 5764 18702
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 6104 18290 6132 19110
rect 6472 18970 6500 19246
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6564 18834 6592 20198
rect 6748 19922 6776 22986
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6840 22030 6868 22646
rect 7024 22216 7052 24618
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7116 23050 7144 24006
rect 7208 23730 7236 25094
rect 7300 24886 7328 25978
rect 7668 24954 7696 26318
rect 7760 24954 7788 26336
rect 7932 26318 7984 26324
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 8312 25974 8340 26318
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7852 25498 7880 25638
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 8404 25362 8432 26182
rect 8588 25906 8616 26182
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8482 25800 8538 25809
rect 8482 25735 8484 25744
rect 8536 25735 8538 25744
rect 8484 25706 8536 25712
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8300 25288 8352 25294
rect 8680 25242 8708 26438
rect 8956 26382 8984 27474
rect 11992 27470 12020 27814
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15752 27600 15804 27606
rect 15752 27542 15804 27548
rect 10140 27464 10192 27470
rect 10416 27464 10468 27470
rect 10140 27406 10192 27412
rect 10230 27432 10286 27441
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9048 27062 9076 27270
rect 9036 27056 9088 27062
rect 9036 26998 9088 27004
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 9416 26586 9444 26726
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8352 25236 8708 25242
rect 8300 25230 8708 25236
rect 8312 25214 8708 25230
rect 8864 25226 8892 26318
rect 9600 26314 9628 27270
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9692 25906 9720 26726
rect 9784 26586 9812 27270
rect 10046 27024 10102 27033
rect 9864 26988 9916 26994
rect 9916 26948 9996 26976
rect 10152 27010 10180 27406
rect 10286 27412 10416 27418
rect 10286 27406 10468 27412
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 10286 27390 10456 27406
rect 10230 27367 10286 27376
rect 10508 27328 10560 27334
rect 10508 27270 10560 27276
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 10102 26982 10180 27010
rect 10046 26959 10102 26968
rect 9864 26930 9916 26936
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9876 26081 9904 26794
rect 9862 26072 9918 26081
rect 9862 26007 9918 26016
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9232 25498 9260 25774
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 9600 25242 9628 25842
rect 9968 25430 9996 26948
rect 10046 26888 10102 26897
rect 10046 26823 10048 26832
rect 10100 26823 10102 26832
rect 10048 26794 10100 26800
rect 10152 26790 10180 26982
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10428 26042 10456 26182
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 9956 25424 10008 25430
rect 9956 25366 10008 25372
rect 10324 25288 10376 25294
rect 8852 25220 8904 25226
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7288 24880 7340 24886
rect 7288 24822 7340 24828
rect 8312 24818 8340 25094
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8588 24750 8616 25214
rect 9600 25214 9720 25242
rect 10324 25230 10376 25236
rect 8852 25162 8904 25168
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 7300 24342 7328 24686
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7288 24336 7340 24342
rect 7288 24278 7340 24284
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7208 22778 7236 23462
rect 7300 23322 7328 24278
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7392 22778 7420 23598
rect 7484 23186 7512 24550
rect 7576 23866 7604 24686
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7564 23860 7616 23866
rect 7564 23802 7616 23808
rect 7472 23180 7524 23186
rect 7472 23122 7524 23128
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7576 22658 7604 23802
rect 7668 23730 7696 24006
rect 7760 23866 7788 24006
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 8220 23662 8248 23734
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7760 23322 7788 23462
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 8220 23066 8248 23598
rect 8312 23186 8340 24550
rect 8588 24206 8616 24686
rect 8772 24206 8800 24754
rect 8864 24342 8892 25162
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24818 9628 25094
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 8588 23594 8616 24142
rect 8772 24070 8800 24142
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8680 23730 8708 23802
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8680 23322 8708 23462
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8576 23112 8628 23118
rect 7748 23044 7800 23050
rect 8220 23038 8340 23066
rect 8576 23054 8628 23060
rect 7748 22986 7800 22992
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 6932 22188 7052 22216
rect 7300 22630 7604 22658
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6840 21554 6868 21966
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6840 21146 6868 21490
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6932 20602 6960 22188
rect 7300 22094 7328 22630
rect 7668 22386 7696 22918
rect 7760 22642 7788 22986
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 8312 22658 8340 23038
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 8116 22636 8168 22642
rect 8312 22630 8432 22658
rect 8116 22578 8168 22584
rect 8128 22438 8156 22578
rect 8300 22568 8352 22574
rect 8298 22536 8300 22545
rect 8352 22536 8354 22545
rect 8298 22471 8354 22480
rect 7484 22358 7696 22386
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 7484 22234 7512 22358
rect 8114 22264 8170 22273
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7564 22228 7616 22234
rect 8114 22199 8170 22208
rect 7564 22170 7616 22176
rect 7024 22066 7328 22094
rect 7024 21622 7052 22066
rect 7576 21690 7604 22170
rect 8128 22098 8156 22199
rect 8206 22128 8262 22137
rect 8116 22092 8168 22098
rect 8262 22086 8340 22114
rect 8404 22098 8432 22630
rect 8206 22063 8262 22072
rect 8116 22034 8168 22040
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7668 21622 7696 21966
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7012 21616 7064 21622
rect 7012 21558 7064 21564
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 7300 20534 7328 20742
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7286 19952 7342 19961
rect 6736 19916 6788 19922
rect 7286 19887 7342 19896
rect 6736 19858 6788 19864
rect 7300 19854 7328 19887
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7196 19780 7248 19786
rect 7196 19722 7248 19728
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 7024 18834 7052 19178
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 5460 18057 5488 18226
rect 5446 18048 5502 18057
rect 5446 17983 5502 17992
rect 6012 17882 6040 18226
rect 6366 17912 6422 17921
rect 6000 17876 6052 17882
rect 6656 17882 6684 18362
rect 7208 18222 7236 19722
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6748 17882 6776 18022
rect 7300 17882 7328 19314
rect 7576 18698 7604 21286
rect 7668 20602 7696 21558
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7760 19514 7788 21830
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8128 20874 8156 21354
rect 8220 20874 8248 21422
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 8208 19848 8260 19854
rect 8312 19836 8340 22086
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 21690 8524 21830
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 20602 8432 21286
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8260 19808 8340 19836
rect 8404 19825 8432 19926
rect 8208 19790 8260 19796
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 8312 19446 8340 19808
rect 8390 19816 8446 19825
rect 8390 19751 8446 19760
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18834 7696 19314
rect 8588 19174 8616 23054
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8680 22273 8708 22646
rect 8666 22264 8722 22273
rect 8666 22199 8722 22208
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7484 18426 7512 18566
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 6366 17847 6422 17856
rect 6644 17876 6696 17882
rect 6000 17818 6052 17824
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 5446 17232 5502 17241
rect 5368 17190 5446 17218
rect 5446 17167 5502 17176
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5460 15162 5488 15438
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5920 15026 5948 15438
rect 6196 15162 6224 15438
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5184 14470 5304 14498
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 2976 13382 3096 13410
rect 3252 13394 3280 13670
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2976 12986 3004 13262
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3068 12782 3096 13382
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3620 13258 3648 13670
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 4172 12986 4200 13874
rect 4264 12986 4292 13942
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4816 13530 4844 13670
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 1412 12238 1440 12718
rect 3068 12442 3096 12718
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 2056 11354 2084 11766
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2516 11218 2544 12242
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3700 12232 3752 12238
rect 3896 12186 3924 12786
rect 3752 12180 3924 12186
rect 3700 12174 3924 12180
rect 3436 11762 3464 12174
rect 3712 12158 3924 12174
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2608 11354 2636 11562
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2976 11257 3004 11630
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 2962 11248 3018 11257
rect 2504 11212 2556 11218
rect 3436 11218 3464 11494
rect 3804 11218 3832 11494
rect 2962 11183 3018 11192
rect 3424 11212 3476 11218
rect 2504 11154 2556 11160
rect 3424 11154 3476 11160
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 2412 11144 2464 11150
rect 2688 11144 2740 11150
rect 2412 11086 2464 11092
rect 2686 11112 2688 11121
rect 2872 11144 2924 11150
rect 2740 11112 2742 11121
rect 2424 10742 2452 11086
rect 2872 11086 2924 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 4252 11144 4304 11150
rect 4356 11132 4384 13262
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4618 11928 4674 11937
rect 4724 11898 4752 12106
rect 4618 11863 4674 11872
rect 4712 11892 4764 11898
rect 4632 11830 4660 11863
rect 4712 11834 4764 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4816 11694 4844 12174
rect 5000 11898 5028 13874
rect 5184 13394 5212 14470
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5080 12776 5132 12782
rect 5078 12744 5080 12753
rect 5132 12744 5134 12753
rect 5078 12679 5134 12688
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4304 11104 4384 11132
rect 4252 11086 4304 11092
rect 2686 11047 2742 11056
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1596 9586 1624 10610
rect 2608 10130 2636 10950
rect 2884 10266 2912 11086
rect 2976 10810 3004 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3344 10266 3372 10746
rect 4264 10674 4292 10950
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 1398 9551 1454 9560
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1596 8634 1624 9522
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1780 8634 1808 9386
rect 2148 9178 2176 9454
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2240 8974 2268 9318
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 1860 8832 1912 8838
rect 2608 8820 2636 10066
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9722 2912 9862
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 9178 2820 9454
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2780 8832 2832 8838
rect 2608 8792 2780 8820
rect 1860 8774 1912 8780
rect 2780 8774 2832 8780
rect 1872 8634 1900 8774
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 6390 1440 7822
rect 1596 7546 1624 8570
rect 2792 8430 2820 8774
rect 2976 8430 3004 9930
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2792 8090 2820 8366
rect 3068 8294 3096 9590
rect 3528 9178 3556 10610
rect 4724 10554 4752 11222
rect 4816 10742 4844 11630
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4724 10526 4844 10554
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4356 10266 4384 10406
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4356 10062 4384 10202
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 8634 3648 9318
rect 3896 9042 3924 9318
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8634 4200 8910
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 8566 4292 8978
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3620 8090 3648 8298
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 3252 6866 3280 7754
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3528 6798 3556 7482
rect 3804 7478 3832 7822
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 7002 3832 7278
rect 3896 7274 3924 8366
rect 4264 8090 4292 8502
rect 4356 8498 4384 9998
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4448 9586 4476 9930
rect 4816 9586 4844 10526
rect 4908 10266 4936 10610
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5000 9466 5028 10610
rect 4816 9438 5028 9466
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4816 7834 4844 9438
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 8634 4936 8910
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5092 8378 5120 12679
rect 5184 12050 5212 13330
rect 5276 12238 5304 14350
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5531 14340 5583 14346
rect 5531 14282 5583 14288
rect 5368 13938 5396 14282
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5368 13394 5396 13874
rect 5552 13530 5580 14282
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5368 12442 5396 13330
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5552 12646 5580 13194
rect 5644 12986 5672 13806
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13530 5764 13670
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5828 12918 5856 14214
rect 5920 13938 5948 14962
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13394 6132 13670
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6288 13190 6316 17614
rect 6380 17202 6408 17847
rect 6644 17818 6696 17824
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6472 16590 6500 17070
rect 6748 16998 6776 17614
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6840 16726 6868 17274
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6932 16590 6960 16934
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6932 16114 6960 16526
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6380 15162 6408 15506
rect 6564 15162 6592 15982
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6748 15706 6776 15846
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6932 14890 6960 15370
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14482 6408 14758
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6748 14278 6776 14826
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5184 12022 5304 12050
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5000 8350 5120 8378
rect 4896 8016 4948 8022
rect 5000 7970 5028 8350
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4948 7964 5028 7970
rect 4896 7958 5028 7964
rect 4908 7942 5028 7958
rect 5092 7954 5120 8230
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 4172 7002 4200 7346
rect 4356 7342 4384 7686
rect 4632 7546 4660 7822
rect 4816 7806 4936 7834
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4356 6934 4384 7278
rect 4908 7274 4936 7806
rect 5000 7410 5028 7942
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5184 7750 5212 11834
rect 5276 10674 5304 12022
rect 5354 11792 5410 11801
rect 5354 11727 5410 11736
rect 5368 10810 5396 11727
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11150 5488 11494
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10062 5304 10474
rect 5368 10062 5396 10746
rect 5552 10674 5580 11222
rect 5644 10810 5672 12718
rect 6288 12714 6316 13126
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6380 12170 6408 13874
rect 6748 13870 6776 14214
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 12986 6684 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6748 12866 6776 13806
rect 6656 12850 6776 12866
rect 6644 12844 6776 12850
rect 6696 12838 6776 12844
rect 6644 12786 6696 12792
rect 6840 12442 6868 13874
rect 6932 12850 6960 13942
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11552 6328 11558
rect 6196 11500 6276 11506
rect 6196 11494 6328 11500
rect 6196 11478 6316 11494
rect 6196 11150 6224 11478
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5736 10266 5764 11086
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6104 10538 6132 10746
rect 6380 10742 6408 11630
rect 6656 11354 6684 12174
rect 6840 11665 6868 12174
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6826 11656 6882 11665
rect 6826 11591 6882 11600
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6748 11218 6776 11290
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10266 5948 10406
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5276 9042 5304 9386
rect 5368 9178 5396 9454
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5368 8974 5396 9114
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 5276 7002 5304 7278
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 5170 6896 5226 6905
rect 3884 6860 3936 6866
rect 5170 6831 5226 6840
rect 3884 6802 3936 6808
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1412 5710 1440 6326
rect 2792 6118 2820 6734
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2332 5710 2360 6054
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 1412 5234 1440 5646
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 4690 1440 5170
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 2446 1440 3878
rect 1872 3534 1900 5646
rect 2792 5370 2820 6054
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2884 5234 2912 6598
rect 3436 5914 3464 6734
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5234 3096 5510
rect 3528 5234 3556 6598
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 5914 3832 6258
rect 3896 6186 3924 6802
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2148 4826 2176 5170
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 3534 1992 4558
rect 2148 4146 2176 4626
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1676 3528 1728 3534
rect 1860 3528 1912 3534
rect 1676 3470 1728 3476
rect 1858 3496 1860 3505
rect 1952 3528 2004 3534
rect 1912 3496 1914 3505
rect 1688 3058 1716 3470
rect 1952 3470 2004 3476
rect 1858 3431 1914 3440
rect 2148 3126 2176 4082
rect 2332 3398 2360 4558
rect 3160 3738 3188 5102
rect 3896 4826 3924 6122
rect 4172 6118 4200 6598
rect 5000 6322 5028 6598
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5710 4200 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5370 5120 5646
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 5092 4622 5120 5102
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4264 4282 4292 4490
rect 4724 4282 4752 4558
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3738 3280 4082
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3160 3590 3648 3618
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2320 3392 2372 3398
rect 2516 3369 2544 3470
rect 3160 3466 3188 3590
rect 3620 3534 3648 3590
rect 4264 3534 4292 3878
rect 4356 3738 4384 4014
rect 4816 4010 4844 4422
rect 5000 4146 5028 4422
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 2320 3334 2372 3340
rect 2502 3360 2558 3369
rect 3252 3346 3280 3470
rect 3436 3398 3464 3470
rect 3424 3392 3476 3398
rect 3252 3318 3372 3346
rect 3424 3334 3476 3340
rect 3790 3360 3846 3369
rect 2502 3295 2558 3304
rect 3344 3194 3372 3318
rect 3790 3295 3846 3304
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 2446 1716 2994
rect 2148 2650 2176 3062
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2650 2544 2790
rect 3252 2650 3280 3130
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2056 2106 2084 2518
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 3240 2440 3292 2446
rect 3424 2440 3476 2446
rect 3292 2400 3424 2428
rect 3240 2382 3292 2388
rect 3424 2382 3476 2388
rect 2148 2106 2176 2382
rect 3148 2304 3200 2310
rect 3528 2292 3556 2450
rect 3200 2264 3556 2292
rect 3148 2246 3200 2252
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2136 2100 2188 2106
rect 2136 2042 2188 2048
rect 3804 800 3832 3295
rect 4080 3058 4108 3470
rect 4724 3058 4752 3606
rect 5092 3482 5120 4558
rect 5184 3670 5212 6831
rect 5368 6798 5396 7686
rect 5460 6866 5488 9998
rect 5552 9722 5580 10066
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5644 9654 5672 9998
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5736 8906 5764 9862
rect 6104 9654 6132 10474
rect 6840 10112 6868 11591
rect 6932 10810 6960 12038
rect 7024 11898 7052 17546
rect 7668 17202 7696 18226
rect 8312 17746 8340 19110
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8404 17746 8432 18566
rect 8496 17814 8524 18566
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8208 17672 8260 17678
rect 8260 17620 8340 17626
rect 8208 17614 8340 17620
rect 8220 17598 8340 17614
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17270 7788 17478
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 8312 17202 8340 17598
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16794 7144 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11014 7144 16118
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7208 12850 7236 14010
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7392 13802 7420 13942
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7208 11914 7236 12650
rect 7392 12646 7420 12718
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12442 7420 12582
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7208 11886 7420 11914
rect 7392 11694 7420 11886
rect 7484 11762 7512 17002
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16794 7604 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7668 15994 7696 17138
rect 8404 17082 8432 17206
rect 8220 17054 8432 17082
rect 8220 16998 8248 17054
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16658 8432 16934
rect 8496 16658 8524 17750
rect 8588 17134 8616 18702
rect 8680 18358 8708 22034
rect 8772 22030 8800 24006
rect 9232 23594 9260 24278
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9220 23588 9272 23594
rect 9220 23530 9272 23536
rect 9232 23118 9260 23530
rect 9324 23118 9352 24006
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9508 23118 9536 23462
rect 9600 23118 9628 24142
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9508 22794 9536 23054
rect 9692 22953 9720 25214
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 24954 10088 25094
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 10336 24886 10364 25230
rect 10324 24880 10376 24886
rect 10324 24822 10376 24828
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10244 23866 10272 24006
rect 10336 23866 10364 24074
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10428 23662 10456 24550
rect 10520 24138 10548 27270
rect 10980 27130 11008 27270
rect 11072 27130 11100 27270
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10784 26852 10836 26858
rect 10784 26794 10836 26800
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 10704 24410 10732 24822
rect 10796 24698 10824 26794
rect 11164 26330 11192 27406
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12912 27130 12940 27338
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13004 27130 13032 27270
rect 13740 27130 13768 27270
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 12452 26518 12480 26794
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 11072 26302 11192 26330
rect 11244 26376 11296 26382
rect 12360 26353 12388 26386
rect 11244 26318 11296 26324
rect 12346 26344 12402 26353
rect 11072 25226 11100 26302
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11164 25294 11192 26182
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 11072 24954 11100 25162
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10796 24670 11192 24698
rect 10876 24608 10928 24614
rect 10928 24568 11100 24596
rect 10876 24550 10928 24556
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 9876 23118 9904 23598
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 9772 22976 9824 22982
rect 9678 22944 9734 22953
rect 9772 22918 9824 22924
rect 9678 22879 9734 22888
rect 9508 22766 9720 22794
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9496 22568 9548 22574
rect 9494 22536 9496 22545
rect 9548 22536 9550 22545
rect 9494 22471 9550 22480
rect 9128 22432 9180 22438
rect 9180 22392 9260 22420
rect 9128 22374 9180 22380
rect 8850 22128 8906 22137
rect 8850 22063 8852 22072
rect 8904 22063 8906 22072
rect 8852 22034 8904 22040
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21622 8984 21830
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9126 21448 9182 21457
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8772 19990 8800 20402
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8772 17814 8800 19654
rect 8864 18766 8892 21286
rect 8956 20466 8984 21422
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 18834 8984 20402
rect 9048 19854 9076 21422
rect 9126 21383 9182 21392
rect 9140 21350 9168 21383
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 20262 9168 20810
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9048 19514 9076 19790
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8956 18426 8984 18770
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8956 17882 8984 18158
rect 9048 18086 9076 19110
rect 9140 18222 9168 19790
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 9048 17218 9076 18022
rect 9140 17882 9168 18158
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8772 17190 9076 17218
rect 8772 17134 8800 17190
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16250 7788 16390
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8496 16250 8524 16594
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8864 16114 8892 17070
rect 8956 16794 8984 17070
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 7576 15966 7696 15994
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7576 15042 7604 15966
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15434 7696 15846
rect 7760 15706 7788 15982
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8680 15706 8708 15846
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7760 15162 7788 15370
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7576 15014 7788 15042
rect 8312 15026 8340 15506
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 14074 7604 14282
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13394 7696 13670
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12986 7604 13262
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7760 12434 7788 15014
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8036 14618 8064 14962
rect 8496 14822 8524 15438
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8022 13968 8078 13977
rect 8022 13903 8024 13912
rect 8076 13903 8078 13912
rect 8024 13874 8076 13880
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7852 13326 7880 13670
rect 7944 13530 7972 13670
rect 8128 13530 8156 13806
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7576 12406 7788 12434
rect 8036 12434 8064 12854
rect 8404 12850 8432 14010
rect 8496 13977 8524 14758
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8482 13968 8538 13977
rect 8482 13903 8538 13912
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13530 8524 13806
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8588 13326 8616 14214
rect 9048 13802 9076 17190
rect 9232 16046 9260 22392
rect 9508 20754 9536 22471
rect 9600 22234 9628 22646
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9692 22114 9720 22766
rect 9600 22086 9720 22114
rect 9600 21690 9628 22086
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9600 20806 9628 21626
rect 9692 21078 9720 21898
rect 9784 21894 9812 22918
rect 10152 22166 10180 22986
rect 9864 22160 9916 22166
rect 9862 22128 9864 22137
rect 10140 22160 10192 22166
rect 9916 22128 9918 22137
rect 10140 22102 10192 22108
rect 9862 22063 9918 22072
rect 10046 21992 10102 22001
rect 9956 21956 10008 21962
rect 10244 21978 10272 23122
rect 10152 21962 10272 21978
rect 10046 21927 10102 21936
rect 10140 21956 10272 21962
rect 9956 21898 10008 21904
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9968 21690 9996 21898
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10060 21570 10088 21927
rect 10192 21950 10272 21956
rect 10140 21898 10192 21904
rect 10060 21542 10180 21570
rect 9864 21344 9916 21350
rect 9784 21304 9864 21332
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9324 20726 9536 20754
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9324 20380 9352 20726
rect 9508 20590 9628 20618
rect 9508 20482 9536 20590
rect 9600 20584 9628 20590
rect 9784 20584 9812 21304
rect 9864 21286 9916 21292
rect 10046 21040 10102 21049
rect 10046 20975 10102 20984
rect 10060 20874 10088 20975
rect 10048 20868 10100 20874
rect 9600 20556 9812 20584
rect 9876 20828 10048 20856
rect 9508 20466 9628 20482
rect 9508 20460 9640 20466
rect 9508 20454 9588 20460
rect 9588 20402 9640 20408
rect 9324 20352 9536 20380
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 18426 9352 19790
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9416 14940 9444 19382
rect 9508 18034 9536 20352
rect 9770 20360 9826 20369
rect 9600 20318 9770 20346
rect 9600 19990 9628 20318
rect 9770 20295 9826 20304
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9876 19378 9904 20828
rect 10048 20810 10100 20816
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 18834 9904 19110
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9508 18006 9812 18034
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 16794 9720 17478
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16250 9720 16526
rect 9784 16454 9812 18006
rect 9876 17338 9904 18634
rect 9968 18290 9996 19926
rect 10060 19378 10088 20198
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10152 18850 10180 21542
rect 10060 18822 10180 18850
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9876 16794 9904 17274
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16114 9812 16390
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9600 15502 9628 15846
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9496 14952 9548 14958
rect 9416 14912 9496 14940
rect 9496 14894 9548 14900
rect 9508 14006 9536 14894
rect 9968 14498 9996 18090
rect 10060 17882 10088 18822
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10060 16658 10088 17818
rect 10152 17678 10180 18702
rect 10244 18290 10272 21950
rect 10336 21894 10364 23190
rect 10888 22710 10916 24006
rect 10968 23588 11020 23594
rect 10968 23530 11020 23536
rect 10980 23050 11008 23530
rect 11072 23050 11100 24568
rect 11164 24426 11192 24670
rect 11256 24614 11284 26318
rect 11704 26308 11756 26314
rect 12346 26279 12402 26288
rect 11704 26250 11756 26256
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11716 25498 11744 26250
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 12360 25294 12388 25842
rect 12452 25838 12480 26454
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12544 25362 12572 26318
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12636 26042 12664 26250
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12728 25838 12756 26522
rect 12820 25838 12848 26930
rect 13268 26920 13320 26926
rect 13268 26862 13320 26868
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 26586 13216 26726
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13280 26382 13308 26862
rect 13924 26586 13952 27406
rect 14660 27130 14688 27406
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 13912 26580 13964 26586
rect 13912 26522 13964 26528
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13910 26344 13966 26353
rect 13910 26279 13966 26288
rect 13924 25922 13952 26279
rect 14188 26240 14240 26246
rect 14188 26182 14240 26188
rect 14200 25974 14228 26182
rect 14292 25974 14320 26930
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14370 26072 14426 26081
rect 14370 26007 14372 26016
rect 14424 26007 14426 26016
rect 14556 26036 14608 26042
rect 14372 25978 14424 25984
rect 14556 25978 14608 25984
rect 13832 25894 13952 25922
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14280 25968 14332 25974
rect 14280 25910 14332 25916
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11164 24398 11284 24426
rect 11256 24206 11284 24398
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 11164 23322 11192 24074
rect 11532 23594 11560 24346
rect 11716 23866 11744 24686
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11256 23186 11284 23530
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 10968 23044 11020 23050
rect 10968 22986 11020 22992
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 10876 22704 10928 22710
rect 10876 22646 10928 22652
rect 10980 22574 11008 22986
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10414 21992 10470 22001
rect 10414 21927 10416 21936
rect 10468 21927 10470 21936
rect 10416 21898 10468 21904
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10428 21078 10456 21490
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10336 20398 10364 21014
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10428 19961 10456 20810
rect 10612 20369 10640 21354
rect 10704 20874 10732 21422
rect 10980 21010 11008 22034
rect 11072 21690 11100 22442
rect 11256 22438 11284 23122
rect 11716 22794 11744 23462
rect 11808 23050 11836 24550
rect 11900 24410 11928 24754
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12176 24410 12204 24686
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11992 23066 12020 24142
rect 12268 23662 12296 24686
rect 12452 24138 12480 25094
rect 12544 24750 12572 25298
rect 12716 24880 12768 24886
rect 12820 24868 12848 25774
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12768 24840 12848 24868
rect 12716 24822 12768 24828
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12440 24132 12492 24138
rect 12440 24074 12492 24080
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 12084 23186 12112 23530
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11716 22766 11836 22794
rect 11900 22778 11928 23054
rect 11992 23038 12112 23066
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11716 22234 11744 22646
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11808 22012 11836 22766
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 12084 22094 12112 23038
rect 12268 22574 12296 23598
rect 12728 23508 12756 24822
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 23866 12848 24550
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12808 23520 12860 23526
rect 12728 23480 12808 23508
rect 12728 23168 12756 23480
rect 12808 23462 12860 23468
rect 12808 23180 12860 23186
rect 12728 23140 12808 23168
rect 12808 23122 12860 23128
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12268 22098 12296 22510
rect 11992 22066 12112 22094
rect 12256 22092 12308 22098
rect 11888 22024 11940 22030
rect 11808 21984 11888 22012
rect 11888 21966 11940 21972
rect 11992 21842 12020 22066
rect 12256 22034 12308 22040
rect 12820 22030 12848 23122
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 11900 21814 12020 21842
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11072 21418 11100 21626
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10888 20466 10916 20742
rect 11256 20534 11284 20878
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 10598 20360 10654 20369
rect 10598 20295 10654 20304
rect 10414 19952 10470 19961
rect 10414 19887 10416 19896
rect 10468 19887 10470 19896
rect 10416 19858 10468 19864
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10336 18970 10364 19246
rect 10520 18970 10548 19790
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10336 18426 10364 18906
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10612 18290 10640 20295
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10704 19514 10732 20198
rect 10796 20058 10824 20402
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10980 19786 11008 20198
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11334 19816 11390 19825
rect 10968 19780 11020 19786
rect 11334 19751 11336 19760
rect 10968 19722 11020 19728
rect 11388 19751 11390 19760
rect 11336 19722 11388 19728
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 11348 19446 11376 19722
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18766 11100 19178
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11808 18970 11836 20402
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11796 18692 11848 18698
rect 11900 18680 11928 21814
rect 12912 21622 12940 24006
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12268 20262 12296 21422
rect 13004 20942 13032 21490
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 19922 12756 20198
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18970 12480 19314
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11848 18652 11928 18680
rect 11796 18634 11848 18640
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10796 18426 10824 18566
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 11072 17921 11100 18566
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11058 17912 11114 17921
rect 11058 17847 11114 17856
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17202 10180 17614
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10060 16182 10088 16458
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 10060 15570 10088 16118
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10152 15706 10180 15982
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14618 10088 14758
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9876 14470 9996 14498
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12850 8616 13126
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8588 12442 8616 12650
rect 8576 12436 8628 12442
rect 8036 12406 8156 12434
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 11688 7432 11694
rect 7576 11642 7604 12406
rect 7760 12374 7788 12406
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11898 7788 12174
rect 8128 12102 8156 12406
rect 8576 12378 8628 12384
rect 9048 12306 9076 13738
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 13190 9260 13262
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9692 12850 9720 13194
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9586 12472 9642 12481
rect 9586 12407 9642 12416
rect 9036 12300 9088 12306
rect 8956 12260 9036 12288
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 7380 11630 7432 11636
rect 7484 11614 7604 11642
rect 8300 11620 8352 11626
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7116 10470 7144 10950
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6748 10084 6868 10112
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 6380 8362 6408 9046
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 5828 7886 5856 8298
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5644 7585 5672 7686
rect 5630 7576 5686 7585
rect 5630 7511 5686 7520
rect 5920 7410 5948 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5460 6322 5488 6802
rect 6012 6458 6040 7890
rect 6380 7886 6408 8298
rect 6748 7886 6776 10084
rect 7012 10056 7064 10062
rect 6840 10016 7012 10044
rect 6840 8974 6868 10016
rect 7012 9998 7064 10004
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6932 9450 6960 9862
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6932 9042 6960 9386
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6104 7546 6132 7822
rect 6366 7576 6422 7585
rect 6092 7540 6144 7546
rect 6366 7511 6422 7520
rect 6092 7482 6144 7488
rect 6380 7410 6408 7511
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6748 6730 6776 7210
rect 6840 7002 6868 8910
rect 7024 8566 7052 9862
rect 7208 9110 7236 10610
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 9178 7420 9522
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7196 9104 7248 9110
rect 7484 9058 7512 11614
rect 8300 11562 8352 11568
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7576 11150 7604 11494
rect 7852 11218 7880 11494
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10062 7604 10950
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7196 9046 7248 9052
rect 7392 9030 7512 9058
rect 7576 9042 7604 9454
rect 7564 9036 7616 9042
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6866 6960 7142
rect 7024 7002 7052 7958
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7206 7144 7754
rect 7300 7750 7328 8230
rect 7392 8022 7420 9030
rect 7564 8978 7616 8984
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 8634 7512 8842
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8430 7604 8978
rect 7668 8566 7696 10134
rect 7760 10062 7788 10746
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 7852 10266 7880 10542
rect 8036 10266 8064 10542
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 8312 9178 8340 11562
rect 8390 11248 8446 11257
rect 8390 11183 8446 11192
rect 8404 11082 8432 11183
rect 8496 11150 8524 11698
rect 8484 11144 8536 11150
rect 8482 11112 8484 11121
rect 8536 11112 8538 11121
rect 8392 11076 8444 11082
rect 8538 11070 8616 11098
rect 8482 11047 8538 11056
rect 8392 11018 8444 11024
rect 8404 10606 8432 11018
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8404 9654 8432 10134
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8496 9382 8524 9998
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7484 7834 7512 8366
rect 7484 7806 7604 7834
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7478 7512 7686
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6380 6458 6408 6666
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 7116 6322 7144 7142
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5234 5304 6190
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 5828 5914 5856 6054
rect 7484 5914 7512 6054
rect 7576 5914 7604 7806
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8404 7426 8432 8774
rect 8312 7410 8432 7426
rect 8300 7404 8432 7410
rect 8352 7398 8432 7404
rect 8300 7346 8352 7352
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6798 8156 7142
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5234 6316 5510
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4826 5304 4966
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5460 4282 5488 5170
rect 5920 4758 5948 5170
rect 6564 5098 6592 5646
rect 6748 5370 6776 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5370 7144 5510
rect 7484 5370 7512 5646
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6656 4826 6684 5102
rect 7576 4826 7604 5646
rect 7668 5234 7696 6054
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7760 5166 7788 5714
rect 8220 5556 8248 6190
rect 8312 5710 8340 6938
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8220 5528 8340 5556
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8312 5302 8340 5528
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4282 5856 4422
rect 6932 4282 6960 4694
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6736 4208 6788 4214
rect 5354 4176 5410 4185
rect 5276 4134 5354 4162
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5170 3496 5226 3505
rect 5092 3454 5170 3482
rect 5170 3431 5172 3440
rect 5224 3431 5226 3440
rect 5172 3402 5224 3408
rect 5276 3194 5304 4134
rect 6736 4150 6788 4156
rect 5354 4111 5410 4120
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5368 3738 5396 4014
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4342 2952 4398 2961
rect 4540 2938 4568 2994
rect 4540 2910 4844 2938
rect 4342 2887 4344 2896
rect 4396 2887 4398 2896
rect 4344 2858 4396 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4172 2514 4200 2790
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4816 2038 4844 2910
rect 5368 2650 5396 3674
rect 5460 2854 5488 4082
rect 5644 3890 5672 4082
rect 6644 4072 6696 4078
rect 6274 4040 6330 4049
rect 6644 4014 6696 4020
rect 6274 3975 6330 3984
rect 5816 3936 5868 3942
rect 5644 3862 5764 3890
rect 5816 3878 5868 3884
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5644 3534 5672 3606
rect 5736 3534 5764 3862
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5828 2514 5856 3878
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6012 3466 6040 3606
rect 6288 3534 6316 3975
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 6472 3194 6500 3878
rect 6550 3768 6606 3777
rect 6550 3703 6606 3712
rect 6564 3448 6592 3703
rect 6656 3602 6684 4014
rect 6748 3602 6776 4150
rect 7024 4010 7052 4626
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 8312 4146 8340 4966
rect 8404 4826 8432 4966
rect 8496 4826 8524 9046
rect 8588 8838 8616 11070
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 8974 8708 9522
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 7886 8616 8298
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8680 6254 8708 8910
rect 8956 8498 8984 12260
rect 9036 12242 9088 12248
rect 9600 11150 9628 12407
rect 9692 11898 9720 12786
rect 9876 12782 9904 14470
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 13530 9996 14282
rect 10060 13870 10088 14554
rect 10244 14482 10272 17546
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10612 17134 10640 17206
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10612 16998 10640 17070
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10230 14376 10286 14385
rect 10152 14006 10180 14350
rect 10230 14311 10286 14320
rect 10244 14278 10272 14311
rect 10336 14278 10364 14894
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12986 9996 13194
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9864 12776 9916 12782
rect 9862 12744 9864 12753
rect 9916 12744 9918 12753
rect 9862 12679 9918 12688
rect 10060 12434 10088 13126
rect 9968 12406 10088 12434
rect 9968 12238 9996 12406
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9784 12050 9812 12174
rect 10152 12050 10180 13942
rect 10336 13394 10364 14214
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 13530 10456 13806
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10520 13530 10548 13738
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12918 10548 13262
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12434 10548 12854
rect 9784 12022 10180 12050
rect 10244 12406 10548 12434
rect 10612 12434 10640 16934
rect 10888 16794 10916 17070
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10704 14618 10732 14758
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10796 13326 10824 16594
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15706 10916 15846
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 14074 10916 14214
rect 10876 14068 10928 14074
rect 11072 14056 11100 16662
rect 11164 16522 11192 18226
rect 11900 18222 11928 18652
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11992 18154 12020 18566
rect 12084 18426 12112 18702
rect 12452 18426 12480 18906
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 11980 18148 12032 18154
rect 11980 18090 12032 18096
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11348 17270 11376 17750
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11624 17542 11652 17614
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11624 17202 11652 17478
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11808 16794 11836 17070
rect 11900 16794 11928 17546
rect 12176 17338 12204 18158
rect 12452 17678 12480 18158
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17338 12296 17478
rect 12636 17338 12664 18702
rect 12728 17746 12756 19858
rect 12912 19514 12940 20742
rect 13004 20330 13032 20878
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19514 13032 19790
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 13096 18970 13124 19654
rect 13188 19394 13216 25638
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13556 24206 13584 24550
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23866 13400 24006
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13280 21146 13308 21898
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13556 20466 13584 20538
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13188 19366 13308 19394
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13188 18426 13216 19246
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 12176 16674 12204 17274
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12176 16646 12296 16674
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 12164 16584 12216 16590
rect 12268 16574 12296 16646
rect 12268 16546 12480 16574
rect 12164 16526 12216 16532
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11256 15502 11284 16526
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11440 15910 11468 16458
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11716 15366 11744 16390
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11072 14028 11284 14056
rect 10876 14010 10928 14016
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12850 10824 13126
rect 10888 12850 10916 13262
rect 10980 12986 11008 13874
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13190 11100 13670
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10612 12406 10824 12434
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9722 9628 9998
rect 9784 9994 9812 12022
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 11694 10088 11834
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 10674 9904 11494
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10810 10088 11086
rect 10152 10810 10180 11290
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 9178 9076 9522
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9178 9260 9318
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8498 9076 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 7954 9352 8298
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7410 9076 7686
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6458 8800 6734
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9048 6322 9076 6666
rect 9508 6662 9536 8434
rect 9588 8016 9640 8022
rect 9586 7984 9588 7993
rect 9640 7984 9642 7993
rect 9586 7919 9642 7928
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7410 9628 7754
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6798 9628 7346
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9692 6662 9720 8502
rect 9784 7888 9812 9930
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 9518 10088 9862
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9178 10088 9454
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10244 8294 10272 12406
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11898 10732 12174
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10796 11150 10824 12406
rect 10888 11762 10916 12786
rect 10980 12714 11008 12922
rect 10968 12708 11020 12714
rect 11020 12668 11100 12696
rect 10968 12650 11020 12656
rect 11072 12442 11100 12668
rect 11256 12481 11284 14028
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11808 12782 11836 13806
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11532 12628 11560 12718
rect 11532 12600 11744 12628
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11242 12472 11298 12481
rect 11369 12475 11677 12484
rect 11060 12436 11112 12442
rect 11716 12442 11744 12600
rect 11242 12407 11298 12416
rect 11704 12436 11756 12442
rect 11060 12378 11112 12384
rect 11256 12374 11284 12407
rect 11900 12434 11928 16458
rect 12176 15502 12204 16526
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11900 12406 12020 12434
rect 11704 12378 11756 12384
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11256 12186 11284 12310
rect 11992 12238 12020 12406
rect 11164 12158 11284 12186
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11060 11688 11112 11694
rect 11058 11656 11060 11665
rect 11112 11656 11114 11665
rect 11058 11591 11114 11600
rect 11164 11218 11192 12158
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11762 11284 12038
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10796 10606 10824 11086
rect 10980 10810 11008 11086
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11518 10704 11574 10713
rect 11518 10639 11574 10648
rect 11532 10606 11560 10639
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11808 10266 11836 10542
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11900 10130 11928 11290
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 10336 8566 10364 9998
rect 10428 8974 10456 9998
rect 11716 9722 11744 9998
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11808 9586 11836 9862
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9178 10640 9318
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10520 8430 10548 8774
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10232 8288 10284 8294
rect 10152 8248 10232 8276
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9772 7882 9824 7888
rect 9772 7824 9824 7830
rect 9784 7478 9812 7824
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9876 7002 9904 7414
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9232 6458 9260 6598
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8956 5370 8984 6258
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9508 5370 9536 6190
rect 9600 6118 9628 6190
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5914 9628 6054
rect 9968 5914 9996 6190
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10060 5817 10088 8026
rect 10046 5808 10102 5817
rect 10046 5743 10048 5752
rect 10100 5743 10102 5752
rect 10048 5714 10100 5720
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 10048 5160 10100 5166
rect 10152 5148 10180 8248
rect 10232 8230 10284 8236
rect 10612 7546 10640 8842
rect 10888 8634 10916 9454
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11900 9042 11928 9862
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11072 8634 11100 8910
rect 11716 8634 11744 8910
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10520 5658 10548 6190
rect 10612 5778 10640 7482
rect 10704 7478 10732 8366
rect 10980 8072 11008 8434
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 10980 8044 11100 8072
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10244 5370 10272 5646
rect 10520 5630 10640 5658
rect 10612 5574 10640 5630
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5370 10640 5510
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10100 5137 10180 5148
rect 10100 5128 10194 5137
rect 10100 5120 10138 5128
rect 10048 5102 10100 5108
rect 10704 5098 10732 7414
rect 10980 6866 11008 7890
rect 11072 6866 11100 8044
rect 11164 7886 11192 8366
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11886 7984 11942 7993
rect 11886 7919 11888 7928
rect 11940 7919 11942 7928
rect 11888 7890 11940 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7750 11192 7822
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7546 11284 7686
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 7002 11192 7142
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11992 6866 12020 12174
rect 12084 11694 12112 15302
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12360 14482 12388 14554
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 14074 12204 14350
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 14074 12296 14214
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12452 13734 12480 16546
rect 12636 16250 12664 17070
rect 12728 16658 12756 17682
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12728 15706 12756 16594
rect 13280 16114 13308 19366
rect 13372 18766 13400 20266
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 20058 13492 20198
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13556 19378 13584 20402
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13648 19310 13676 21286
rect 13740 21146 13768 21490
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20890 13860 25894
rect 13912 25764 13964 25770
rect 13912 25706 13964 25712
rect 13924 25498 13952 25706
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14016 24206 14044 24346
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 13924 21894 13952 24142
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 23186 14044 24006
rect 14108 23866 14136 25230
rect 14200 24954 14228 25910
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14200 23866 14228 24006
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14108 23202 14136 23802
rect 14004 23180 14056 23186
rect 14108 23174 14228 23202
rect 14004 23122 14056 23128
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14108 22234 14136 23054
rect 14200 22642 14228 23174
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14292 21690 14320 23054
rect 14384 22778 14412 24142
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 14476 22506 14504 24074
rect 14568 23032 14596 25978
rect 14660 24800 14688 26250
rect 14752 25838 14780 27270
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15120 26228 15148 26794
rect 15212 26382 15240 27270
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15120 26200 15240 26228
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 15212 25294 15240 26200
rect 15304 25906 15332 26726
rect 15396 25906 15424 27542
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15488 25650 15516 26454
rect 15764 25838 15792 27542
rect 18708 27538 18736 29200
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 19156 27600 19208 27606
rect 19156 27542 19208 27548
rect 21364 27600 21416 27606
rect 21364 27542 21416 27548
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15856 26586 15884 27406
rect 16488 27396 16540 27402
rect 16488 27338 16540 27344
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16316 26994 16344 27270
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 16500 26450 16528 27338
rect 16868 27130 16896 27474
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 17420 26994 17448 27270
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 16120 25696 16172 25702
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 14752 24954 14780 25094
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 15212 24818 15240 25094
rect 15304 24818 15332 25638
rect 15488 25622 15608 25650
rect 16120 25638 16172 25644
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15200 24812 15252 24818
rect 14660 24772 14780 24800
rect 14752 24732 14780 24772
rect 15200 24754 15252 24760
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 14924 24744 14976 24750
rect 14752 24704 14924 24732
rect 14924 24686 14976 24692
rect 15396 24614 15424 25298
rect 15488 24954 15516 25434
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 15016 24336 15068 24342
rect 15016 24278 15068 24284
rect 14752 23866 14780 24278
rect 15028 24206 15056 24278
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 15396 23866 15424 24142
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 14568 23004 14688 23032
rect 14554 22944 14610 22953
rect 14554 22879 14610 22888
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 13832 20862 13952 20890
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13648 18290 13676 19246
rect 13740 19242 13768 20198
rect 13832 19854 13860 20742
rect 13924 20262 13952 20862
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13924 19990 13952 20198
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13728 18760 13780 18766
rect 13832 18748 13860 19246
rect 13780 18720 13860 18748
rect 13728 18702 13780 18708
rect 13740 18358 13768 18702
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13648 17542 13676 18226
rect 13740 17678 13768 18294
rect 13832 18154 13860 18566
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13464 17338 13492 17478
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13648 17202 13676 17478
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 16590 13676 17138
rect 13740 16590 13768 17614
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12728 15094 12756 15642
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 14074 12940 14214
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12986 12204 13126
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12360 12442 12388 13398
rect 12452 12730 12480 13670
rect 12544 13530 12572 13806
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 12866 12572 13466
rect 12728 12986 12756 13806
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 12986 12940 13330
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12544 12838 12848 12866
rect 12452 12702 12664 12730
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12440 12096 12492 12102
rect 12544 12084 12572 12582
rect 12636 12434 12664 12702
rect 12820 12442 12848 12838
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12436 12860 12442
rect 12636 12406 12756 12434
rect 12544 12056 12664 12084
rect 12440 12038 12492 12044
rect 12176 11898 12204 12038
rect 12452 11898 12480 12038
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12636 11762 12664 12056
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 7342 12112 11630
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10606 12664 11086
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12360 10130 12388 10406
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9722 12572 9998
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12728 9586 12756 12406
rect 12808 12378 12860 12384
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 11898 12848 12242
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12808 11756 12860 11762
rect 12912 11744 12940 12718
rect 13004 12442 13032 16050
rect 13648 16046 13676 16526
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14550 13492 14758
rect 13740 14618 13768 14962
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13832 14498 13860 18090
rect 14016 17814 14044 20402
rect 14568 19446 14596 22879
rect 14660 20466 14688 23004
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 14752 22778 14780 22918
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 15212 22574 15240 22918
rect 15488 22778 15516 24006
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15200 22568 15252 22574
rect 15120 22528 15200 22556
rect 15120 22234 15148 22528
rect 15200 22510 15252 22516
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 15580 22094 15608 25622
rect 16132 25498 16160 25638
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15672 24954 15700 25094
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15764 22574 15792 24006
rect 16040 23730 16068 24754
rect 16316 24206 16344 25162
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 16040 22642 16068 23666
rect 16316 23662 16344 24142
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16316 22642 16344 23598
rect 16500 23050 16528 25366
rect 16592 23118 16620 26726
rect 17500 26512 17552 26518
rect 17500 26454 17552 26460
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16684 25702 16712 26318
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 16960 25294 16988 26182
rect 17052 25498 17080 26318
rect 17512 25906 17540 26454
rect 17696 26450 17724 27270
rect 18340 27130 18368 27406
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18892 27130 18920 27270
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18880 27124 18932 27130
rect 18880 27066 18932 27072
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 24818 16804 25094
rect 17236 24886 17264 25638
rect 17328 25362 17356 25638
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17420 25276 17448 25774
rect 17500 25288 17552 25294
rect 17420 25248 17500 25276
rect 17500 25230 17552 25236
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24410 16988 24550
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 17052 23186 17080 23462
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 17224 23112 17276 23118
rect 17512 23100 17540 25230
rect 17604 24682 17632 26250
rect 17788 25922 17816 26862
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 17788 25894 17908 25922
rect 18524 25906 18552 26250
rect 18892 26246 18920 26522
rect 19168 26382 19196 27542
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 19260 26586 19288 26726
rect 19352 26586 19380 27270
rect 19536 27130 19564 27406
rect 19616 27328 19668 27334
rect 19616 27270 19668 27276
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19628 26586 19656 27270
rect 20824 27062 20852 27270
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 19248 26580 19300 26586
rect 19248 26522 19300 26528
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 20180 25974 20208 26318
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17788 25498 17816 25774
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17880 25294 17908 25894
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18696 25832 18748 25838
rect 20536 25832 20588 25838
rect 18696 25774 18748 25780
rect 20534 25800 20536 25809
rect 20588 25800 20590 25809
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18708 25498 18736 25774
rect 20534 25735 20590 25744
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 20352 25696 20404 25702
rect 20548 25684 20576 25735
rect 20404 25656 20576 25684
rect 20352 25638 20404 25644
rect 18800 25498 18828 25638
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 17696 25158 17724 25230
rect 17684 25152 17736 25158
rect 17684 25094 17736 25100
rect 17880 24954 17908 25230
rect 19076 24954 19104 25230
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 17592 24676 17644 24682
rect 17592 24618 17644 24624
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 18248 24410 18276 24550
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 19536 24410 19564 24550
rect 19628 24410 19656 24550
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 19524 24404 19576 24410
rect 19524 24346 19576 24352
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23730 17632 24006
rect 18248 23866 18276 24346
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18892 23798 18920 24006
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17604 23322 17632 23666
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 23322 18092 23598
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17592 23112 17644 23118
rect 17512 23072 17592 23100
rect 17224 23054 17276 23060
rect 17592 23054 17644 23060
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 16316 22234 16344 22578
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 15304 22066 15608 22094
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14936 21146 14964 21286
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 15028 20924 15056 21490
rect 15212 21049 15240 21490
rect 15198 21040 15254 21049
rect 15198 20975 15254 20984
rect 15304 20942 15332 22066
rect 15580 21962 15608 22066
rect 16592 22030 16620 23054
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17144 22778 17172 22918
rect 17236 22778 17264 23054
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17604 22574 17632 23054
rect 19352 23050 19380 23530
rect 19628 23050 19656 24006
rect 19720 23798 19748 25094
rect 20640 24818 20668 26726
rect 21100 26586 21128 27406
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21284 26586 21312 27270
rect 21376 27130 21404 27542
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 22388 27130 22416 27406
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 27130 22784 27270
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 21376 26586 21404 27066
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21284 26382 21312 26522
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21468 25974 21496 26930
rect 22744 26920 22796 26926
rect 22742 26888 22744 26897
rect 22796 26888 22798 26897
rect 22742 26823 22798 26832
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21560 26586 21588 26726
rect 21548 26580 21600 26586
rect 21548 26522 21600 26528
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 22296 26042 22324 26182
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 21192 25498 21220 25774
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 24954 20760 25230
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19720 23186 19748 23734
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19616 23044 19668 23050
rect 19616 22986 19668 22992
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18524 22778 18552 22918
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 18144 22568 18196 22574
rect 18328 22568 18380 22574
rect 18144 22510 18196 22516
rect 18248 22528 18328 22556
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17696 22030 17724 22374
rect 18156 22234 18184 22510
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15764 21146 15792 21422
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15200 20936 15252 20942
rect 15028 20896 15200 20924
rect 15200 20878 15252 20884
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 15212 20602 15240 20878
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 20058 14872 20266
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 15366 14044 17614
rect 14200 16590 14228 19314
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18970 14504 19246
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17338 14320 17614
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14108 15502 14136 16050
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13924 14618 13952 15098
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14016 14618 14044 14894
rect 14108 14822 14136 15438
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13832 14470 14044 14498
rect 13084 14408 13136 14414
rect 13360 14408 13412 14414
rect 13136 14356 13360 14362
rect 13084 14350 13412 14356
rect 13096 14334 13400 14350
rect 13372 14074 13400 14334
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13188 12832 13216 13330
rect 13372 12986 13400 14010
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13530 13584 13874
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 12986 13492 13194
rect 13648 12986 13676 13262
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13360 12844 13412 12850
rect 13188 12804 13360 12832
rect 13188 12714 13216 12804
rect 13360 12786 13412 12792
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13912 12640 13964 12646
rect 14016 12628 14044 14470
rect 14200 14278 14228 15846
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14292 14074 14320 16050
rect 14476 15094 14504 16730
rect 14568 15978 14596 19382
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15162 14596 15914
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 14482 14596 14894
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14385 14596 14418
rect 14554 14376 14610 14385
rect 14554 14311 14610 14320
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12986 14136 13126
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12918 14228 13942
rect 14660 13462 14688 18702
rect 15304 18630 15332 20878
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15396 20058 15424 20334
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15396 19514 15424 19790
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14752 16454 14780 17614
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 16130 14780 16390
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 15212 16250 15240 16934
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15304 16250 15332 16458
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14752 16102 15056 16130
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14936 15706 14964 15846
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15028 15638 15056 16102
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 14832 15428 14884 15434
rect 14752 15388 14832 15416
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14096 12708 14148 12714
rect 14200 12696 14228 12854
rect 14292 12782 14320 13126
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14148 12668 14228 12696
rect 14096 12650 14148 12656
rect 13964 12600 14044 12628
rect 13912 12582 13964 12588
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13004 11880 13032 12378
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13464 11898 13492 12174
rect 13452 11892 13504 11898
rect 13004 11852 13216 11880
rect 13084 11756 13136 11762
rect 12860 11716 13084 11744
rect 12808 11698 12860 11704
rect 13084 11698 13136 11704
rect 13188 11150 13216 11852
rect 13452 11834 13504 11840
rect 13556 11762 13584 12174
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12820 10606 12848 10746
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 9110 12756 9522
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 13004 8498 13032 10610
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10062 13768 10542
rect 13924 10198 13952 12582
rect 14108 12374 14136 12650
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14292 12238 14320 12718
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14108 11150 14136 12038
rect 14200 11898 14228 12038
rect 14292 11898 14320 12174
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14476 11898 14504 12106
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 11286 14504 11630
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14476 10606 14504 11222
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10810 14596 11086
rect 14660 10810 14688 11222
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9178 13216 9454
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6186 10824 6734
rect 11072 6186 11100 6802
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5914 11100 6122
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11716 5914 11744 6734
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 10138 5063 10194 5072
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7288 4072 7340 4078
rect 8128 4049 8156 4082
rect 8208 4072 8260 4078
rect 7288 4014 7340 4020
rect 8114 4040 8170 4049
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3505 6776 3538
rect 6828 3528 6880 3534
rect 6734 3496 6790 3505
rect 6644 3460 6696 3466
rect 6564 3420 6644 3448
rect 6828 3470 6880 3476
rect 6734 3431 6790 3440
rect 6644 3402 6696 3408
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6840 2990 6868 3470
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7024 2650 7052 3946
rect 7300 3738 7328 4014
rect 8208 4014 8260 4020
rect 8114 3975 8170 3984
rect 8220 3738 8248 4014
rect 8588 3942 8616 4558
rect 8680 4486 8708 4966
rect 8772 4690 8800 4966
rect 10244 4690 10364 4706
rect 11256 4690 11284 5782
rect 11808 5642 11836 6258
rect 11992 5710 12020 6666
rect 12084 6458 12112 6666
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12072 6316 12124 6322
rect 12176 6304 12204 8434
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 8090 12756 8230
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13556 7886 13584 9522
rect 13740 8974 13768 9998
rect 13924 9722 13952 10134
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14108 9722 14136 9862
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9178 14136 9318
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 12268 7002 12296 7822
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12452 7002 12480 7754
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7478 13216 7686
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12360 6458 12388 6870
rect 12544 6458 12572 7278
rect 13096 7002 13124 7278
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13464 6934 13492 7346
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12124 6276 12204 6304
rect 12440 6316 12492 6322
rect 12072 6258 12124 6264
rect 12440 6258 12492 6264
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11532 5370 11560 5578
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11808 5234 11836 5578
rect 12084 5302 12112 6258
rect 12452 6186 12480 6258
rect 13556 6254 13584 7822
rect 13740 6882 13768 7890
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13648 6854 13768 6882
rect 13648 6798 13676 6854
rect 14016 6798 14044 7822
rect 14108 7546 14136 8434
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5914 12848 6122
rect 13096 5914 13124 6190
rect 13188 5914 13216 6190
rect 13372 5914 13400 6190
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 10232 4684 10364 4690
rect 10284 4678 10364 4684
rect 10232 4626 10284 4632
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4146 10180 4422
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 9140 3777 9168 4014
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9126 3768 9182 3777
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 8208 3732 8260 3738
rect 9324 3738 9352 3878
rect 9692 3738 9720 3878
rect 9876 3738 9904 3878
rect 9126 3703 9182 3712
rect 9312 3732 9364 3738
rect 8208 3674 8260 3680
rect 9312 3674 9364 3680
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3194 7788 3334
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 8680 3194 8708 3470
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6274 2544 6330 2553
rect 5816 2508 5868 2514
rect 6274 2479 6330 2488
rect 5816 2450 5868 2456
rect 6288 2446 6316 2479
rect 6276 2440 6328 2446
rect 5998 2408 6054 2417
rect 6276 2382 6328 2388
rect 8036 2378 8064 2994
rect 8220 2514 8248 3062
rect 8588 2650 8616 3130
rect 9692 2774 9720 3402
rect 9692 2746 9904 2774
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 5998 2343 6054 2352
rect 8024 2372 8076 2378
rect 6012 2310 6040 2343
rect 8024 2314 8076 2320
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 9876 1834 9904 2746
rect 10060 2650 10088 3470
rect 10336 3466 10364 4678
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10336 2650 10364 3402
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10428 2038 10456 2518
rect 10520 2446 10548 4014
rect 10612 3942 10640 4558
rect 11256 4146 11284 4626
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4146 11376 4490
rect 11808 4486 11836 5170
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3058 10640 3334
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10888 2650 10916 3470
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 2650 11192 3402
rect 11256 3058 11284 4082
rect 11348 4026 11376 4082
rect 11348 3998 11744 4026
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11716 3602 11744 3998
rect 12452 3738 12480 5102
rect 12544 3942 12572 5102
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4826 12848 4966
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13096 4758 13124 5238
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12820 3738 12848 4490
rect 13096 4282 13124 4694
rect 13372 4282 13400 4966
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13464 4554 13492 4762
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 13096 3534 13124 4218
rect 13556 4214 13584 5102
rect 13648 4826 13676 6394
rect 14108 5273 14136 6598
rect 14200 6458 14228 9046
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14292 7886 14320 8570
rect 14568 8090 14596 9862
rect 14660 9722 14688 10746
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6798 14320 7346
rect 14476 6798 14504 7822
rect 14568 7002 14596 7822
rect 14660 7546 14688 8230
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14646 6896 14702 6905
rect 14646 6831 14702 6840
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14188 6316 14240 6322
rect 14292 6304 14320 6734
rect 14660 6662 14688 6831
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14240 6276 14320 6304
rect 14188 6258 14240 6264
rect 14094 5264 14150 5273
rect 14094 5199 14150 5208
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 11428 3528 11480 3534
rect 13084 3528 13136 3534
rect 11428 3470 11480 3476
rect 12346 3496 12402 3505
rect 11440 3194 11468 3470
rect 13084 3470 13136 3476
rect 13556 3466 13584 4150
rect 13740 4078 13768 4694
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13832 3738 13860 4014
rect 14108 3738 14136 4422
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 12346 3431 12402 3440
rect 13544 3460 13596 3466
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 12360 3126 12388 3431
rect 13544 3402 13596 3408
rect 14016 3194 14044 3606
rect 14200 3534 14228 6258
rect 14660 6118 14688 6598
rect 14752 6225 14780 15388
rect 14832 15370 14884 15376
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 15304 14482 15332 15846
rect 15396 15026 15424 19110
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15580 18426 15608 18702
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15672 17882 15700 20810
rect 15750 20632 15806 20641
rect 15750 20567 15806 20576
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15672 17626 15700 17818
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15580 17598 15700 17626
rect 15488 17202 15516 17546
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15488 16794 15516 17138
rect 15580 17134 15608 17598
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17338 15700 17478
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15672 16046 15700 17070
rect 15764 16658 15792 20567
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19990 15884 20198
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15856 19718 15884 19926
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15856 17678 15884 18158
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15948 15178 15976 21490
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16132 21146 16160 21286
rect 16316 21146 16344 21966
rect 16592 21622 16620 21966
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 17512 21554 17540 21830
rect 18248 21690 18276 22528
rect 18328 22510 18380 22516
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18786 22128 18842 22137
rect 18786 22063 18842 22072
rect 18800 21894 18828 22063
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18708 21554 18736 21830
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 16488 21480 16540 21486
rect 16486 21448 16488 21457
rect 16540 21448 16542 21457
rect 16486 21383 16542 21392
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 16500 20602 16528 20878
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 17052 20466 17080 20742
rect 17236 20602 17264 20878
rect 17512 20602 17540 20878
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17972 20466 18000 20742
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 20058 16252 20198
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16316 19938 16344 20402
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16224 19910 16344 19938
rect 16224 19854 16252 19910
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16224 19378 16252 19790
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16316 19446 16344 19722
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18426 16068 18566
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16040 17746 16068 18362
rect 16224 18290 16252 19314
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 17338 16160 17614
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16114 16252 16730
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16316 15366 16344 19382
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17746 16528 18022
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16794 16436 16934
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16500 16522 16528 17138
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15580 15150 15976 15178
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15488 14958 15516 15098
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 15304 12986 15332 13262
rect 15580 13258 15608 15150
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15764 13410 15792 14962
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 14074 15884 14214
rect 15948 14074 15976 14894
rect 16132 14550 16160 15302
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 14074 16068 14350
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16040 13530 16068 14010
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15672 13382 15792 13410
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 15304 10266 15332 12174
rect 15580 11898 15608 12174
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11082 15700 13382
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12850 15792 13194
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 11898 16252 12174
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15396 10198 15424 10610
rect 15672 10606 15700 11018
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10674 15884 10950
rect 16040 10810 16068 11086
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16040 10266 16068 10406
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 16040 9586 16068 10202
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15120 9178 15148 9454
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 7857 15148 8434
rect 15106 7848 15162 7857
rect 15106 7783 15162 7792
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 15212 7546 15240 7686
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15108 6724 15160 6730
rect 15160 6684 15240 6712
rect 15108 6666 15160 6672
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 15212 6458 15240 6684
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15304 6458 15332 6598
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 14738 6216 14794 6225
rect 14738 6151 14794 6160
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 15396 5930 15424 6598
rect 15304 5902 15424 5930
rect 14370 5808 14426 5817
rect 15304 5778 15332 5902
rect 15488 5794 15516 9318
rect 15856 9178 15884 9454
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8838 15976 8910
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16040 8548 16068 8842
rect 15948 8520 16068 8548
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 7002 15608 7346
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 14370 5743 14372 5752
rect 14424 5743 14426 5752
rect 15292 5772 15344 5778
rect 14372 5714 14424 5720
rect 15292 5714 15344 5720
rect 15396 5766 15516 5794
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 14384 5522 14412 5578
rect 14556 5568 14608 5574
rect 14384 5494 14504 5522
rect 14556 5510 14608 5516
rect 14280 5160 14332 5166
rect 14278 5128 14280 5137
rect 14372 5160 14424 5166
rect 14332 5128 14334 5137
rect 14372 5102 14424 5108
rect 14278 5063 14334 5072
rect 14384 4826 14412 5102
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3194 14228 3470
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2514 11284 2994
rect 13360 2848 13412 2854
rect 13188 2796 13360 2802
rect 13188 2790 13412 2796
rect 13188 2774 13400 2790
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11348 2038 11376 2382
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 11256 870 11376 898
rect 11256 800 11284 870
rect 3790 0 3846 800
rect 11242 0 11298 800
rect 11348 762 11376 870
rect 11624 762 11652 1974
rect 13096 1834 13124 2518
rect 13188 2446 13216 2774
rect 14476 2650 14504 5494
rect 14568 5302 14596 5510
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14936 2446 14964 3130
rect 15212 2650 15240 5578
rect 15396 5030 15424 5766
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5370 15516 5510
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15304 4146 15332 4626
rect 15672 4162 15700 8298
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 8090 15884 8230
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15764 6662 15792 7482
rect 15948 7002 15976 8520
rect 16132 8498 16160 9998
rect 16316 9994 16344 15302
rect 16592 14074 16620 20266
rect 16868 20058 16896 20334
rect 17604 20058 17632 20402
rect 17972 20058 18000 20402
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 17236 19718 17264 19790
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 18064 19514 18092 19790
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17316 19372 17368 19378
rect 18064 19334 18092 19450
rect 18248 19394 18276 20810
rect 18340 20602 18368 21014
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 17316 19314 17368 19320
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18426 17264 18566
rect 17328 18426 17356 19314
rect 17880 19306 18092 19334
rect 18144 19372 18196 19378
rect 18248 19366 18368 19394
rect 18144 19314 18196 19320
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17604 18766 17632 19110
rect 17880 18970 17908 19306
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17236 16794 17264 17546
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17328 16794 17356 16934
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16684 15910 16712 16526
rect 17236 16250 17264 16730
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17512 16114 17540 16934
rect 17604 16794 17632 18702
rect 17880 18426 17908 18906
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17788 17610 17816 18022
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17972 17338 18000 18158
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 18064 17542 18092 18090
rect 18156 17814 18184 19314
rect 18340 19310 18368 19366
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18708 18766 18736 19654
rect 18892 19242 18920 20878
rect 18984 20398 19012 22986
rect 19352 22574 19380 22986
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 22234 19656 22374
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19812 21622 19840 24686
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 23798 20116 24550
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 19996 23526 20024 23734
rect 20640 23662 20668 24074
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19904 22710 19932 22918
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19890 22264 19946 22273
rect 19890 22199 19946 22208
rect 19904 22030 19932 22199
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19996 21690 20024 21966
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 19812 20942 19840 21558
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 20942 20116 21286
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19812 20534 19840 20878
rect 20272 20602 20300 23598
rect 20640 23118 20668 23598
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20732 23050 20760 24142
rect 21008 23866 21036 24142
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20996 23248 21048 23254
rect 20996 23190 21048 23196
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22642 20760 22986
rect 20720 22636 20772 22642
rect 20640 22596 20720 22624
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20456 22098 20484 22442
rect 20548 22234 20576 22442
rect 20640 22250 20668 22596
rect 20720 22578 20772 22584
rect 20824 22574 20852 23054
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20536 22228 20588 22234
rect 20640 22222 20760 22250
rect 20824 22234 20852 22510
rect 20536 22170 20588 22176
rect 20444 22092 20496 22098
rect 20732 22094 20760 22222
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20732 22066 20852 22094
rect 20444 22034 20496 22040
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 19800 20528 19852 20534
rect 19800 20470 19852 20476
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18984 19310 19012 20334
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19628 19446 19656 19654
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18892 18970 18920 19178
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 19352 17882 19380 18294
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 19628 17678 19656 19382
rect 19904 18426 19932 19450
rect 20088 19378 20116 20266
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20456 18834 20484 22034
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20548 21486 20576 21830
rect 20640 21554 20668 21830
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20824 21010 20852 22066
rect 20916 21554 20944 22918
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19248 17672 19300 17678
rect 19076 17632 19248 17660
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15706 17264 15846
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17224 15496 17276 15502
rect 17130 15464 17186 15473
rect 17224 15438 17276 15444
rect 17130 15399 17186 15408
rect 17144 14890 17172 15399
rect 17236 15162 17264 15438
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17604 15026 17632 15302
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 14482 17172 14826
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16592 12986 16620 13670
rect 16776 12986 16804 14350
rect 17696 14074 17724 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17420 13394 17448 14010
rect 17408 13388 17460 13394
rect 17328 13348 17408 13376
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12374 16712 12718
rect 16776 12442 16804 12922
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16776 10130 16804 10406
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 17052 9926 17080 11834
rect 17328 11218 17356 13348
rect 17408 13330 17460 13336
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10742 17172 10950
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17144 10112 17172 10678
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10266 17264 10542
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17224 10124 17276 10130
rect 17144 10084 17224 10112
rect 17224 10066 17276 10072
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17236 9382 17264 10066
rect 17420 9586 17448 13126
rect 17788 11801 17816 17138
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14618 18000 14758
rect 17960 14612 18012 14618
rect 18012 14572 18092 14600
rect 17960 14554 18012 14560
rect 18064 14328 18092 14572
rect 18156 14482 18184 16050
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18524 14958 18552 15302
rect 18892 15162 18920 15438
rect 18984 15366 19012 16390
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18248 14618 18276 14894
rect 18524 14822 18552 14894
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18064 14300 18644 14328
rect 18616 13938 18644 14300
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18696 13932 18748 13938
rect 18800 13920 18828 14350
rect 18748 13892 18828 13920
rect 18696 13874 18748 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13326 18000 13738
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18800 13326 18828 13892
rect 18892 13870 18920 15098
rect 18984 14414 19012 15302
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18984 13734 19012 13942
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 17972 12850 18000 13262
rect 17960 12844 18012 12850
rect 18012 12804 18092 12832
rect 17960 12786 18012 12792
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17972 12238 18000 12582
rect 18064 12238 18092 12804
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18156 12442 18184 12650
rect 18248 12646 18276 13262
rect 18340 12986 18368 13262
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17774 11792 17830 11801
rect 17774 11727 17830 11736
rect 17498 11656 17554 11665
rect 17498 11591 17554 11600
rect 17512 11218 17540 11591
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17788 11150 17816 11727
rect 18248 11506 18276 12582
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18800 12306 18828 13262
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18064 11478 18276 11506
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17696 9926 17724 11086
rect 18064 10606 18092 11478
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18156 10810 18184 10950
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16868 9042 16896 9318
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16304 8968 16356 8974
rect 16210 8936 16266 8945
rect 16304 8910 16356 8916
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16764 8968 16816 8974
rect 17236 8956 17264 9318
rect 17328 9178 17356 9454
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17316 8968 17368 8974
rect 17236 8928 17316 8956
rect 16764 8910 16816 8916
rect 17316 8910 17368 8916
rect 16210 8871 16266 8880
rect 16224 8838 16252 8871
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16120 8492 16172 8498
rect 16040 8452 16120 8480
rect 16040 7002 16068 8452
rect 16120 8434 16172 8440
rect 16212 7880 16264 7886
rect 16316 7868 16344 8910
rect 16500 8634 16528 8910
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16264 7840 16344 7868
rect 16212 7822 16264 7828
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7206 16160 7686
rect 16224 7546 16252 7822
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 5914 15792 6598
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15764 4826 15792 5850
rect 15856 5545 15884 6734
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15842 5536 15898 5545
rect 15842 5471 15898 5480
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15292 4140 15344 4146
rect 15672 4134 15792 4162
rect 15292 4082 15344 4088
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15672 3942 15700 3975
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15304 2650 15332 2790
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15672 2446 15700 3878
rect 15764 3097 15792 4134
rect 15948 3369 15976 6598
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 16040 5914 16068 6122
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16040 3534 16068 4762
rect 16132 4690 16160 7142
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16500 6610 16528 8570
rect 16592 6866 16620 8910
rect 16776 8090 16804 8910
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16684 7041 16712 7346
rect 16670 7032 16726 7041
rect 16670 6967 16726 6976
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16578 6760 16634 6769
rect 16578 6695 16580 6704
rect 16632 6695 16634 6704
rect 16764 6724 16816 6730
rect 16580 6666 16632 6672
rect 16764 6666 16816 6672
rect 16670 6624 16726 6633
rect 16224 6202 16252 6598
rect 16316 6304 16344 6598
rect 16500 6582 16670 6610
rect 16670 6559 16726 6568
rect 16316 6276 16436 6304
rect 16224 6174 16344 6202
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5914 16252 6054
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16224 4282 16252 4626
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15934 3360 15990 3369
rect 15934 3295 15990 3304
rect 16132 3194 16160 4082
rect 16316 4049 16344 6174
rect 16302 4040 16358 4049
rect 16302 3975 16358 3984
rect 16408 3369 16436 6276
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 5370 16528 5646
rect 16592 5370 16620 5782
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16592 4622 16620 5306
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16684 3670 16712 6559
rect 16776 6390 16804 6666
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16776 5710 16804 6054
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16776 3738 16804 4014
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16672 3664 16724 3670
rect 16776 3641 16804 3674
rect 16672 3606 16724 3612
rect 16762 3632 16818 3641
rect 16762 3567 16818 3576
rect 16868 3534 16896 8774
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17052 6798 17080 8434
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7342 17172 7822
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 7342 17264 7686
rect 17328 7478 17356 8910
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17316 7472 17368 7478
rect 17420 7449 17448 8366
rect 17316 7414 17368 7420
rect 17406 7440 17462 7449
rect 17406 7375 17462 7384
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17328 6798 17356 7210
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4826 16988 5102
rect 17144 4826 17172 5510
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17236 3738 17264 5850
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17328 5234 17356 5306
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17420 4593 17448 6598
rect 17406 4584 17462 4593
rect 17406 4519 17462 4528
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 16856 3528 16908 3534
rect 17328 3505 17356 3878
rect 16856 3470 16908 3476
rect 17314 3496 17370 3505
rect 16764 3460 16816 3466
rect 17314 3431 17370 3440
rect 16764 3402 16816 3408
rect 16580 3392 16632 3398
rect 16394 3360 16450 3369
rect 16580 3334 16632 3340
rect 16394 3295 16450 3304
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15750 3088 15806 3097
rect 16592 3058 16620 3334
rect 16776 3126 16804 3402
rect 17420 3194 17448 3878
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 15750 3023 15806 3032
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16776 2774 16804 3062
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16684 2746 16804 2774
rect 16684 2514 16712 2746
rect 16960 2650 16988 2926
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 13188 2310 13216 2382
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 13648 2038 13676 2246
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 15488 2038 15516 2246
rect 13636 2032 13688 2038
rect 13636 1974 13688 1980
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 16776 1834 16804 2382
rect 17512 1970 17540 8774
rect 17604 8401 17632 8774
rect 17590 8392 17646 8401
rect 17590 8327 17646 8336
rect 17696 7546 17724 9386
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 8498 17816 9318
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8498 17908 8774
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 8378 17908 8434
rect 17788 8350 17908 8378
rect 17788 7886 17816 8350
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 8022 17908 8230
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17590 6896 17646 6905
rect 17590 6831 17592 6840
rect 17644 6831 17646 6840
rect 17592 6802 17644 6808
rect 17696 6118 17724 7278
rect 17972 6934 18000 10202
rect 18156 9586 18184 10746
rect 18248 10674 18276 10950
rect 18708 10742 18736 11494
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 6934 18092 8774
rect 18248 8566 18276 9930
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18708 8786 18736 10542
rect 18800 10062 18828 10950
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18892 9994 18920 12786
rect 19076 11694 19104 17632
rect 19248 17614 19300 17620
rect 19616 17672 19668 17678
rect 20456 17660 20484 18770
rect 20548 17678 20576 20198
rect 20824 20058 20852 20946
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20916 19990 20944 21082
rect 21008 20890 21036 23190
rect 21100 22642 21128 24822
rect 21284 23662 21312 25842
rect 21560 25702 21588 25978
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21548 25696 21600 25702
rect 21548 25638 21600 25644
rect 21376 25498 21404 25638
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21928 25362 21956 25842
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 21468 24750 21496 25298
rect 22020 25294 22048 25774
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22572 25498 22600 25638
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 22204 24834 22232 25094
rect 22112 24818 22232 24834
rect 22100 24812 22232 24818
rect 22152 24806 22232 24812
rect 22100 24754 22152 24760
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21376 22094 21404 24074
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 21468 23730 21496 24006
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21468 23322 21496 23666
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21560 23254 21588 24006
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22204 23610 22232 24006
rect 22112 23582 22232 23610
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 22112 23186 22140 23582
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22204 23322 22232 23462
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 21640 23044 21692 23050
rect 21640 22986 21692 22992
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 21560 22098 21588 22918
rect 21652 22624 21680 22986
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 22296 22642 22324 24210
rect 22480 24206 22508 24550
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22388 23662 22416 24074
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22008 22636 22060 22642
rect 21652 22596 22008 22624
rect 22008 22578 22060 22584
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22388 22574 22416 23598
rect 22480 23118 22508 24142
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22572 23730 22600 24006
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22480 22506 22508 23054
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 21916 22500 21968 22506
rect 21916 22442 21968 22448
rect 22008 22500 22060 22506
rect 22008 22442 22060 22448
rect 22468 22500 22520 22506
rect 22468 22442 22520 22448
rect 21928 22273 21956 22442
rect 21914 22264 21970 22273
rect 21914 22199 21970 22208
rect 21376 22066 21496 22094
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21100 21418 21128 21966
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21376 21350 21404 21966
rect 21468 21434 21496 22066
rect 21548 22092 21600 22098
rect 22020 22094 22048 22442
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 21548 22034 21600 22040
rect 21652 22066 22048 22094
rect 21652 21554 21680 22066
rect 22204 21894 22232 22374
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21468 21406 21588 21434
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21364 20936 21416 20942
rect 21008 20862 21128 20890
rect 21364 20878 21416 20884
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 21008 20398 21036 20742
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20824 18290 20852 19110
rect 20916 18834 20944 19926
rect 21008 19417 21036 20334
rect 20994 19408 21050 19417
rect 20994 19343 20996 19352
rect 21048 19343 21050 19352
rect 20996 19314 21048 19320
rect 21100 19281 21128 20862
rect 21376 20777 21404 20878
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21008 18426 21036 18702
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 19616 17614 19668 17620
rect 19904 17632 20484 17660
rect 20536 17672 20588 17678
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 16250 19288 17138
rect 19536 16998 19564 17478
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19168 15570 19196 15982
rect 19352 15910 19380 16526
rect 19444 15978 19472 16526
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19154 15464 19210 15473
rect 19260 15450 19288 15506
rect 19210 15422 19288 15450
rect 19352 15434 19380 15846
rect 19340 15428 19392 15434
rect 19154 15399 19210 15408
rect 19340 15370 19392 15376
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19168 14618 19196 14894
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19260 14498 19288 14894
rect 19168 14482 19288 14498
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19156 14476 19288 14482
rect 19208 14470 19288 14476
rect 19156 14418 19208 14424
rect 19444 14278 19472 14486
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19260 12442 19288 12718
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19536 11830 19564 16934
rect 19628 16794 19656 17614
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16794 19748 16934
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19628 13938 19656 16730
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19628 13530 19656 13670
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19812 12345 19840 14962
rect 19904 14958 19932 17632
rect 20536 17614 20588 17620
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20442 17232 20498 17241
rect 20442 17167 20444 17176
rect 20496 17167 20498 17176
rect 20444 17138 20496 17144
rect 20732 17134 20760 17546
rect 20916 17270 20944 18226
rect 21100 17490 21128 19207
rect 21008 17462 21128 17490
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20626 16688 20682 16697
rect 20626 16623 20628 16632
rect 20680 16623 20682 16632
rect 20628 16594 20680 16600
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20272 16250 20300 16526
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 16250 20392 16390
rect 20548 16250 20576 16526
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20534 16144 20590 16153
rect 20534 16079 20590 16088
rect 20548 15706 20576 16079
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19904 13530 19932 14894
rect 19996 14006 20024 15302
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20088 14618 20116 14894
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19996 12442 20024 12718
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19798 12336 19854 12345
rect 19798 12271 19854 12280
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19430 11248 19486 11257
rect 19430 11183 19432 11192
rect 19484 11183 19486 11192
rect 19432 11154 19484 11160
rect 19536 10810 19564 11766
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19168 10130 19196 10474
rect 19720 10470 19748 10746
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18892 9654 18920 9930
rect 18984 9926 19012 9998
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 19168 9674 19196 10066
rect 18880 9648 18932 9654
rect 19168 9646 19288 9674
rect 18880 9590 18932 9596
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 9178 18828 9454
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18708 8758 19012 8786
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18156 7002 18184 7346
rect 18144 6996 18196 7002
rect 18248 6984 18276 7754
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18432 7410 18460 7686
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18524 7342 18552 7686
rect 18616 7546 18644 7822
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18248 6956 18368 6984
rect 18144 6938 18196 6944
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5574 17724 6054
rect 17788 5710 17816 6598
rect 17880 5914 17908 6734
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17972 5794 18000 6054
rect 17880 5766 18000 5794
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17880 5166 17908 5766
rect 18248 5574 18276 6598
rect 18340 6118 18368 6956
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18420 6656 18472 6662
rect 18524 6633 18552 6734
rect 18420 6598 18472 6604
rect 18510 6624 18566 6633
rect 18432 6254 18460 6598
rect 18510 6559 18566 6568
rect 18616 6458 18644 6802
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18616 6254 18644 6394
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18604 5840 18656 5846
rect 18326 5808 18382 5817
rect 18604 5782 18656 5788
rect 18326 5743 18382 5752
rect 18340 5710 18368 5743
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18616 5370 18644 5782
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 17592 5160 17644 5166
rect 17868 5160 17920 5166
rect 17592 5102 17644 5108
rect 17774 5128 17830 5137
rect 17604 2990 17632 5102
rect 17868 5102 17920 5108
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17774 5063 17830 5072
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17696 2446 17724 4966
rect 17788 4622 17816 5063
rect 17972 4826 18000 5102
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 18064 4554 18092 4966
rect 18248 4706 18276 5306
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18156 4690 18276 4706
rect 18144 4684 18276 4690
rect 18196 4678 18276 4684
rect 18144 4626 18196 4632
rect 18708 4570 18736 8570
rect 18788 8084 18840 8090
rect 18840 8044 18920 8072
rect 18788 8026 18840 8032
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18800 5137 18828 5238
rect 18786 5128 18842 5137
rect 18786 5063 18842 5072
rect 18432 4554 18736 4570
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18420 4548 18736 4554
rect 18472 4542 18736 4548
rect 18788 4548 18840 4554
rect 18420 4490 18472 4496
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17788 2446 17816 3130
rect 17880 2582 17908 3402
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17972 2514 18000 4150
rect 18064 4078 18092 4490
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18064 3058 18092 3130
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18156 2854 18184 4490
rect 18524 3942 18552 4542
rect 18788 4490 18840 4496
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18512 3936 18564 3942
rect 18708 3913 18736 4082
rect 18512 3878 18564 3884
rect 18694 3904 18750 3913
rect 18315 3836 18623 3845
rect 18694 3839 18750 3848
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18800 3754 18828 4490
rect 18708 3726 18828 3754
rect 18708 3670 18736 3726
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18248 2378 18276 3334
rect 18708 3194 18736 3606
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3194 18828 3334
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 13084 1828 13136 1834
rect 13084 1770 13136 1776
rect 16764 1828 16816 1834
rect 16764 1770 16816 1776
rect 18708 800 18736 2790
rect 18892 2774 18920 8044
rect 18984 7041 19012 8758
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 8090 19104 8230
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19076 7954 19104 8026
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19168 7478 19196 9522
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 18970 7032 19026 7041
rect 18970 6967 19026 6976
rect 19260 6882 19288 9646
rect 19444 9518 19472 10134
rect 19720 10130 19748 10406
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19430 9344 19486 9353
rect 19352 9302 19430 9330
rect 19352 8566 19380 9302
rect 19430 9279 19486 9288
rect 19536 9178 19564 9454
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19614 9208 19670 9217
rect 19524 9172 19576 9178
rect 19614 9143 19670 9152
rect 19524 9114 19576 9120
rect 19628 9042 19656 9143
rect 19720 9042 19748 9318
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19352 7478 19380 8502
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 18984 6854 19288 6882
rect 18984 6338 19012 6854
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6497 19104 6598
rect 19062 6488 19118 6497
rect 19062 6423 19118 6432
rect 18984 6310 19104 6338
rect 19168 6322 19196 6666
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6322 19288 6598
rect 19352 6458 19380 6734
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 6322 19472 8502
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19536 7274 19564 7686
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 18970 5128 19026 5137
rect 18970 5063 19026 5072
rect 18984 3534 19012 5063
rect 19076 4026 19104 6310
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19168 6174 19380 6202
rect 19168 6118 19196 6174
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5914 19288 6054
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19168 4214 19196 5510
rect 19260 5234 19288 5850
rect 19352 5574 19380 6174
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19352 5001 19380 5238
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19340 4820 19392 4826
rect 19260 4780 19340 4808
rect 19156 4208 19208 4214
rect 19156 4150 19208 4156
rect 19260 4078 19288 4780
rect 19340 4762 19392 4768
rect 19248 4072 19300 4078
rect 19076 4020 19248 4026
rect 19076 4014 19300 4020
rect 19076 3998 19288 4014
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19168 3126 19196 3402
rect 19352 3398 19380 3946
rect 19444 3602 19472 6258
rect 19536 5302 19564 7210
rect 19628 7177 19656 8774
rect 19720 8634 19748 8774
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7546 19748 7822
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19614 7168 19670 7177
rect 19614 7103 19670 7112
rect 19614 6488 19670 6497
rect 19614 6423 19670 6432
rect 19628 5710 19656 6423
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19720 5556 19748 7210
rect 19812 5930 19840 10406
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 8974 19932 9998
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19996 8566 20024 10542
rect 20076 9512 20128 9518
rect 20074 9480 20076 9489
rect 20128 9480 20130 9489
rect 20074 9415 20130 9424
rect 20180 9178 20208 14894
rect 20548 13734 20576 15642
rect 20640 15638 20668 15914
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20732 15094 20760 17070
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20824 16250 20852 17002
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16454 20944 16934
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20824 15570 20852 15914
rect 20916 15570 20944 16390
rect 21008 16153 21036 17462
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20994 16144 21050 16153
rect 20994 16079 21050 16088
rect 21100 15570 21128 17274
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20824 15162 20852 15302
rect 21192 15178 21220 20538
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21284 19334 21312 20470
rect 21468 19786 21496 21286
rect 21560 20602 21588 21406
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21454 19408 21510 19417
rect 21364 19346 21416 19352
rect 21284 19306 21364 19334
rect 21454 19343 21456 19352
rect 21508 19343 21510 19352
rect 21456 19314 21508 19320
rect 21364 19288 21416 19294
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 16114 21312 18566
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 21100 15150 21220 15178
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 21100 15026 21128 15150
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20824 14618 20852 14894
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 21008 14414 21036 14758
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20916 14074 20944 14350
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 12850 20300 13126
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20074 9072 20130 9081
rect 20180 9042 20208 9114
rect 20074 9007 20130 9016
rect 20168 9036 20220 9042
rect 20088 8974 20116 9007
rect 20168 8978 20220 8984
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 20088 8412 20116 8502
rect 19996 8384 20116 8412
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 7002 19932 7346
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19996 6798 20024 8384
rect 20074 8120 20130 8129
rect 20074 8055 20076 8064
rect 20128 8055 20130 8064
rect 20076 8026 20128 8032
rect 20180 7970 20208 8978
rect 20088 7954 20208 7970
rect 20076 7948 20208 7954
rect 20128 7942 20208 7948
rect 20076 7890 20128 7896
rect 20272 7546 20300 11630
rect 20350 9616 20406 9625
rect 20456 9602 20484 13466
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20916 12986 20944 13262
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12442 20760 12718
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20824 12306 20852 12582
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20916 11150 20944 11290
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20916 10062 20944 11086
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9722 20760 9930
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20456 9574 20576 9602
rect 20350 9551 20352 9560
rect 20404 9551 20406 9560
rect 20352 9522 20404 9528
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20364 8106 20392 9318
rect 20456 8673 20484 9318
rect 20548 9058 20576 9574
rect 20628 9580 20680 9586
rect 20732 9568 20760 9658
rect 20902 9616 20958 9625
rect 20680 9540 20760 9568
rect 20824 9574 20902 9602
rect 20628 9522 20680 9528
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 9104 20680 9110
rect 20548 9052 20628 9058
rect 20548 9046 20680 9052
rect 20548 9030 20668 9046
rect 20732 9042 20760 9318
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20442 8664 20498 8673
rect 20548 8634 20576 8910
rect 20442 8599 20498 8608
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20364 8078 20576 8106
rect 20640 8090 20668 9030
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20732 8566 20760 8842
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20732 8090 20760 8502
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19812 5902 19932 5930
rect 19904 5778 19932 5902
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19812 5658 19840 5714
rect 19812 5630 19932 5658
rect 19996 5642 20024 6734
rect 19800 5568 19852 5574
rect 19720 5528 19800 5556
rect 19800 5510 19852 5516
rect 19904 5522 19932 5630
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 20088 5522 20116 7346
rect 20272 6390 20300 7482
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 19812 5386 19840 5510
rect 19904 5494 20116 5522
rect 19812 5358 20024 5386
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19720 4282 19748 4558
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3602 19564 4082
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19432 3120 19484 3126
rect 19536 3108 19564 3538
rect 19484 3080 19564 3108
rect 19432 3062 19484 3068
rect 19628 3040 19656 3674
rect 18800 2746 18920 2774
rect 19536 3012 19656 3040
rect 18800 1766 18828 2746
rect 19536 2446 19564 3012
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19812 2038 19840 2926
rect 19904 2650 19932 5238
rect 19996 4842 20024 5358
rect 20074 4856 20130 4865
rect 19996 4814 20074 4842
rect 19996 4146 20024 4814
rect 20074 4791 20130 4800
rect 20272 4554 20300 6326
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20456 5302 20484 5646
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20272 4214 20300 4490
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20272 3602 20300 4150
rect 20260 3596 20312 3602
rect 20180 3556 20260 3584
rect 20180 3126 20208 3556
rect 20260 3538 20312 3544
rect 20364 3398 20392 5034
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20456 3194 20484 3402
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19996 2650 20024 2858
rect 20548 2774 20576 8078
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20824 7970 20852 9574
rect 21008 9586 21036 13398
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10742 21128 10950
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20902 9551 20958 9560
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 9024 21036 9522
rect 20732 7942 20852 7970
rect 20916 8996 21036 9024
rect 20732 5953 20760 7942
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20824 6254 20852 7822
rect 20916 7750 20944 8996
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21008 8634 21036 8842
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21100 8537 21128 9998
rect 21192 9874 21220 15030
rect 21284 14482 21312 15642
rect 21376 15162 21404 17138
rect 21468 16658 21496 18702
rect 21652 18290 21680 19994
rect 21744 19990 21772 20198
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21744 19854 21772 19926
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22204 18426 22232 21490
rect 22296 21146 22324 21966
rect 22572 21570 22600 22714
rect 22664 21894 22692 23598
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22572 21542 22692 21570
rect 22664 21486 22692 21542
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22652 21480 22704 21486
rect 22756 21457 22784 26823
rect 22848 26450 22876 27406
rect 23676 26586 23704 27610
rect 26160 27554 26188 29200
rect 26240 27600 26292 27606
rect 26160 27548 26240 27554
rect 26160 27542 26292 27548
rect 26608 27600 26660 27606
rect 26608 27542 26660 27548
rect 26160 27526 26280 27542
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24044 26926 24072 27338
rect 24136 27010 24164 27406
rect 24136 26994 24256 27010
rect 24136 26988 24268 26994
rect 24136 26982 24216 26988
rect 24216 26930 24268 26936
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22848 25906 22876 26386
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 23112 25832 23164 25838
rect 23112 25774 23164 25780
rect 23124 25498 23152 25774
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23400 25294 23428 26318
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23584 25906 23612 26182
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 24320 25838 24348 26726
rect 24872 26586 24900 26862
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 24964 26042 24992 26454
rect 25056 26450 25084 27406
rect 26068 27130 26096 27406
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26528 26994 26556 27270
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 25688 26920 25740 26926
rect 25686 26888 25688 26897
rect 25740 26888 25742 26897
rect 25686 26823 25742 26832
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 25792 26382 25820 26930
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 26424 26920 26476 26926
rect 26424 26862 26476 26868
rect 26160 26450 26188 26862
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25148 26246 25176 26318
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 25608 26042 25636 26318
rect 25792 26246 25820 26318
rect 25780 26240 25832 26246
rect 25780 26182 25832 26188
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24044 25498 24072 25638
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23124 24614 23152 25230
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 24044 24886 24072 25094
rect 24216 24948 24268 24954
rect 24216 24890 24268 24896
rect 24032 24880 24084 24886
rect 24032 24822 24084 24828
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23124 24206 23152 24550
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 23186 22876 24006
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 23124 23050 23152 24142
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23798 23244 24006
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23492 23730 23520 24550
rect 23584 24410 23612 24550
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23664 24336 23716 24342
rect 23664 24278 23716 24284
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23400 23322 23428 23462
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 22928 21480 22980 21486
rect 22652 21422 22704 21428
rect 22742 21448 22798 21457
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22282 20632 22338 20641
rect 22282 20567 22284 20576
rect 22336 20567 22338 20576
rect 22284 20538 22336 20544
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22296 18426 22324 20334
rect 22388 19922 22416 21422
rect 22928 21422 22980 21428
rect 22742 21383 22798 21392
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22480 19514 22508 19654
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22480 18426 22508 18634
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 21640 18284 21692 18290
rect 21560 18244 21640 18272
rect 21560 17882 21588 18244
rect 21640 18226 21692 18232
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 22008 17672 22060 17678
rect 22112 17660 22140 18226
rect 22060 17632 22140 17660
rect 22008 17614 22060 17620
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22204 16794 22232 17478
rect 22572 17202 22600 19722
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22756 18630 22784 19654
rect 22848 19242 22876 20470
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 22940 19122 22968 21422
rect 23032 21010 23060 22374
rect 23308 22098 23336 23190
rect 23492 23186 23520 23666
rect 23584 23322 23612 23802
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23676 23118 23704 24278
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23768 23866 23796 24006
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23860 23322 23888 24074
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23584 22778 23612 23054
rect 24136 22778 24164 23054
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23492 22030 23520 22374
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23400 21554 23428 21830
rect 23768 21690 23796 22170
rect 24044 22030 24072 22578
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23124 19446 23152 20402
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 22848 19094 22968 19122
rect 22848 18630 22876 19094
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22756 18290 22784 18566
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22848 18170 22876 18566
rect 23216 18222 23244 21422
rect 23676 21146 23704 21422
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23492 20466 23520 21082
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23492 18970 23520 19722
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23768 18850 23796 21422
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 20942 23980 21286
rect 24044 20942 24072 21966
rect 24136 21010 24164 22374
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20602 24072 20742
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23860 19922 23888 20470
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23676 18822 23796 18850
rect 22756 18142 22876 18170
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 16130 21588 16526
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21652 16250 21680 16390
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21468 16114 21588 16130
rect 21456 16108 21588 16114
rect 21508 16102 21588 16108
rect 21456 16050 21508 16056
rect 21468 15434 21496 16050
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21652 14958 21680 15438
rect 21836 15434 21864 15982
rect 22204 15502 22232 16730
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22296 15706 22324 16390
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 22388 15094 22416 16458
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22020 14618 22048 14894
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21468 14074 21496 14282
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 13326 21496 13874
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21284 11830 21312 13194
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12374 21404 13126
rect 21468 12850 21496 13262
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21468 10606 21496 12310
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21364 10192 21416 10198
rect 21362 10160 21364 10169
rect 21416 10160 21418 10169
rect 21362 10095 21418 10104
rect 21192 9846 21404 9874
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21086 8528 21142 8537
rect 20996 8492 21048 8498
rect 21086 8463 21142 8472
rect 20996 8434 21048 8440
rect 21008 7970 21036 8434
rect 21192 8106 21220 9658
rect 21270 9616 21326 9625
rect 21270 9551 21272 9560
rect 21324 9551 21326 9560
rect 21272 9522 21324 9528
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21284 8401 21312 9318
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 21192 8078 21312 8106
rect 21008 7942 21128 7970
rect 21284 7954 21312 8078
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20718 5944 20774 5953
rect 20718 5879 20774 5888
rect 20824 5658 20852 6190
rect 20916 5914 20944 6802
rect 21008 6322 21036 7686
rect 21100 7206 21128 7942
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 7546 21220 7686
rect 21284 7546 21312 7890
rect 21376 7546 21404 9846
rect 21468 8498 21496 10406
rect 21560 8974 21588 13806
rect 21652 11830 21680 14214
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22204 12986 22232 13738
rect 22296 13394 22324 14418
rect 22480 14362 22508 15438
rect 22572 14618 22600 15438
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22664 14550 22692 16118
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22388 14334 22508 14362
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21836 12646 21864 12854
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12442 22140 12582
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21652 11150 21680 11494
rect 22020 11354 22048 11766
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21652 10742 21680 11086
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22296 10742 22324 10950
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22190 10568 22246 10577
rect 22190 10503 22246 10512
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10266 22140 10406
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21640 10192 21692 10198
rect 21640 10134 21692 10140
rect 21730 10160 21786 10169
rect 21652 9722 21680 10134
rect 21730 10095 21732 10104
rect 21784 10095 21786 10104
rect 21732 10066 21784 10072
rect 22204 10062 22232 10503
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21822 9616 21878 9625
rect 21822 9551 21878 9560
rect 22008 9580 22060 9586
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21744 9217 21772 9454
rect 21730 9208 21786 9217
rect 21640 9172 21692 9178
rect 21730 9143 21786 9152
rect 21640 9114 21692 9120
rect 21652 8974 21680 9114
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21836 8820 21864 9551
rect 22008 9522 22060 9528
rect 22020 8838 22048 9522
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22112 9178 22140 9454
rect 22296 9217 22324 9454
rect 22282 9208 22338 9217
rect 22100 9172 22152 9178
rect 22282 9143 22338 9152
rect 22100 9114 22152 9120
rect 21560 8792 21864 8820
rect 22008 8832 22060 8838
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 8294 21496 8434
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21454 8120 21510 8129
rect 21454 8055 21510 8064
rect 21468 8022 21496 8055
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21560 7426 21588 8792
rect 22112 8820 22140 9114
rect 22112 8792 22232 8820
rect 22008 8774 22060 8780
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 22204 8634 22232 8792
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22020 8090 22048 8434
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22204 7546 22232 7822
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 21284 7398 21588 7426
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21284 6633 21312 7398
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21468 6866 21496 7142
rect 21560 7002 21588 7142
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21270 6624 21326 6633
rect 21270 6559 21326 6568
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20640 5630 20852 5658
rect 20640 5370 20668 5630
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20732 4826 20760 5170
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20640 3942 20668 4558
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20364 2746 20576 2774
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20364 2514 20392 2746
rect 20640 2514 20668 3606
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20824 2446 20852 5306
rect 21284 5234 21312 6559
rect 21376 5914 21404 6666
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21560 5817 21588 6734
rect 21546 5808 21602 5817
rect 21546 5743 21602 5752
rect 21454 5536 21510 5545
rect 21454 5471 21510 5480
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21100 4758 21128 5102
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21192 4214 21220 4966
rect 21468 4282 21496 5471
rect 21652 5234 21680 7414
rect 22006 7032 22062 7041
rect 22204 7002 22232 7482
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22006 6967 22062 6976
rect 22192 6996 22244 7002
rect 22020 6662 22048 6967
rect 22192 6938 22244 6944
rect 22296 6934 22324 7278
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 22296 6458 22324 6870
rect 22388 6866 22416 14334
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12986 22508 13262
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22572 12850 22600 13670
rect 22664 12986 22692 14486
rect 22756 13326 22784 18142
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17338 23152 17614
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23216 16697 23244 18158
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23492 17678 23520 18022
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23308 17202 23336 17546
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23202 16688 23258 16697
rect 23202 16623 23258 16632
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 23032 16046 23060 16390
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23032 15502 23060 15982
rect 23216 15570 23244 16623
rect 23400 16590 23428 16934
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23400 16114 23428 16390
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23492 16046 23520 17070
rect 23584 16046 23612 17750
rect 23676 17626 23704 18822
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23768 18426 23796 18702
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23952 18222 23980 19110
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23768 17882 23796 18158
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23860 17814 23888 18022
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23676 17598 23796 17626
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23676 17338 23704 17478
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23768 17202 23796 17598
rect 23860 17338 23888 17750
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 14822 22968 15302
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 23032 14634 23060 15438
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 22940 14606 23060 14634
rect 22940 13938 22968 14606
rect 23124 14414 23152 15302
rect 23216 14414 23244 15370
rect 23400 15026 23428 15846
rect 23492 15366 23520 15982
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23032 13938 23060 14350
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22756 11694 22784 12106
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22756 9586 22784 11630
rect 22848 9586 22876 13738
rect 22940 12850 22968 13874
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 23032 12434 23060 13262
rect 23216 12986 23244 13262
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23308 12850 23336 14214
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 22940 12406 23060 12434
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22756 9466 22784 9522
rect 22756 9438 22876 9466
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9178 22784 9318
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22480 8498 22508 8910
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8634 22600 8774
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22756 8498 22784 9114
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22480 8294 22508 8434
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22558 7576 22614 7585
rect 22664 7546 22692 8230
rect 22848 8090 22876 9438
rect 22940 8430 22968 12406
rect 23296 12232 23348 12238
rect 23584 12186 23612 15846
rect 24044 15706 24072 15846
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13326 23704 13670
rect 23952 13462 23980 15438
rect 24044 15026 24072 15642
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14414 24072 14758
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23676 12714 23704 13262
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12986 23796 13126
rect 23860 12986 23888 13398
rect 24044 13326 24072 14350
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23952 12714 23980 13262
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 24044 12238 24072 13262
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 23296 12174 23348 12180
rect 23308 11830 23336 12174
rect 23400 12158 23612 12186
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 11150 23060 11494
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23308 10742 23336 11766
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23124 10130 23152 10678
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23032 9466 23060 10066
rect 23216 9586 23244 10202
rect 23308 10062 23336 10678
rect 23400 10674 23428 12158
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23492 10962 23520 11562
rect 23584 11150 23612 12038
rect 24030 11928 24086 11937
rect 24030 11863 24086 11872
rect 24044 11762 24072 11863
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23756 11688 23808 11694
rect 24136 11642 24164 12242
rect 23756 11630 23808 11636
rect 23676 11354 23704 11630
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23492 10934 23704 10962
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23584 9994 23612 10406
rect 23572 9988 23624 9994
rect 23572 9930 23624 9936
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23032 9450 23152 9466
rect 23032 9444 23164 9450
rect 23032 9438 23112 9444
rect 23112 9386 23164 9392
rect 23124 9042 23152 9386
rect 23308 9353 23336 9522
rect 23294 9344 23350 9353
rect 23294 9279 23350 9288
rect 23492 9110 23520 9862
rect 23480 9104 23532 9110
rect 23480 9046 23532 9052
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22756 7546 22784 7686
rect 22558 7511 22614 7520
rect 22652 7540 22704 7546
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21928 4865 21956 5170
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 21914 4856 21970 4865
rect 22112 4826 22140 5034
rect 22204 5001 22232 5034
rect 22190 4992 22246 5001
rect 22190 4927 22246 4936
rect 22388 4826 22416 5034
rect 21914 4791 21970 4800
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21180 4208 21232 4214
rect 21180 4150 21232 4156
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21376 3738 21404 3878
rect 21468 3738 21496 3878
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 20994 3632 21050 3641
rect 20994 3567 21050 3576
rect 21008 2922 21036 3567
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21284 3058 21312 3334
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20916 2530 20944 2790
rect 21560 2582 21588 4082
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 21914 2680 21970 2689
rect 21914 2615 21970 2624
rect 21548 2576 21600 2582
rect 20916 2514 21128 2530
rect 21548 2518 21600 2524
rect 21928 2514 21956 2615
rect 22572 2553 22600 7511
rect 22652 7482 22704 7488
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22664 5234 22692 6258
rect 22756 5794 22784 7482
rect 22940 6866 22968 7686
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 23032 6390 23060 8774
rect 23492 8634 23520 8910
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23216 8090 23244 8366
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 22834 6216 22890 6225
rect 22890 6174 22968 6202
rect 22834 6151 22890 6160
rect 22756 5778 22876 5794
rect 22756 5772 22888 5778
rect 22756 5766 22836 5772
rect 22836 5714 22888 5720
rect 22940 5710 22968 6174
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22664 3890 22692 5170
rect 22744 3936 22796 3942
rect 22664 3884 22744 3890
rect 22940 3913 22968 5646
rect 22664 3878 22796 3884
rect 22926 3904 22982 3913
rect 22664 3862 22784 3878
rect 22664 3194 22692 3862
rect 22926 3839 22982 3848
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22940 2774 22968 3839
rect 22848 2746 22968 2774
rect 22558 2544 22614 2553
rect 20916 2508 21140 2514
rect 20916 2502 21088 2508
rect 21088 2450 21140 2456
rect 21916 2508 21968 2514
rect 22848 2514 22876 2746
rect 23124 2514 23152 8026
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 5370 23244 7890
rect 23400 7721 23428 8298
rect 23386 7712 23442 7721
rect 23386 7647 23442 7656
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23492 7410 23520 7482
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23216 3942 23244 4558
rect 23308 4486 23336 7142
rect 23400 6934 23428 7278
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23584 6866 23612 8298
rect 23676 7426 23704 10934
rect 23768 9722 23796 11630
rect 24044 11614 24164 11642
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23952 10062 23980 10678
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23860 9722 23888 9998
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23846 9072 23902 9081
rect 23846 9007 23902 9016
rect 23860 8401 23888 9007
rect 23952 8566 23980 9998
rect 24044 9674 24072 11614
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11354 24164 11494
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24136 11150 24164 11290
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24228 11014 24256 24890
rect 24412 24410 24440 25842
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24596 25226 24624 25638
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24872 24818 24900 25162
rect 25792 25158 25820 26182
rect 26068 26042 26096 26182
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26252 25838 26280 26182
rect 26344 25906 26372 26726
rect 26436 26450 26464 26862
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26240 25832 26292 25838
rect 25870 25800 25926 25809
rect 26240 25774 26292 25780
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 25870 25735 25926 25744
rect 25884 25362 25912 25735
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24596 23730 24624 24550
rect 24688 24410 24716 24618
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24688 23594 24716 24142
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24688 23186 24716 23530
rect 24872 23526 24900 24074
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 24320 20602 24348 21014
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24412 19666 24440 21966
rect 24688 21622 24716 23122
rect 24872 22778 24900 23462
rect 24964 23118 24992 24006
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 25056 23526 25084 23734
rect 25148 23662 25176 24754
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25608 24206 25636 25094
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25700 24410 25728 24686
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25516 24052 25544 24142
rect 25792 24052 25820 25094
rect 25976 24410 26004 25230
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 26068 24206 26096 24754
rect 26252 24682 26280 25094
rect 26528 24954 26556 25774
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26528 24206 26556 24754
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 25516 24024 25820 24052
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24780 22098 24808 22374
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24676 21616 24728 21622
rect 24676 21558 24728 21564
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24504 21146 24532 21422
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24688 20534 24716 21558
rect 24872 21554 24900 22714
rect 25608 22642 25636 24024
rect 26068 23730 26096 24142
rect 26620 24018 26648 27542
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 27804 27396 27856 27402
rect 27804 27338 27856 27344
rect 27252 27056 27304 27062
rect 27252 26998 27304 27004
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26712 26450 26740 26726
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 26804 24954 26832 25230
rect 26792 24948 26844 24954
rect 26792 24890 26844 24896
rect 26792 24132 26844 24138
rect 26792 24074 26844 24080
rect 26528 23990 26648 24018
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 26068 23322 26096 23666
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26068 22778 26096 23258
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 22778 26372 22918
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 26240 22500 26292 22506
rect 26240 22442 26292 22448
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24964 21690 24992 22034
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 24860 21548 24912 21554
rect 24780 21508 24860 21536
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24780 20466 24808 21508
rect 24860 21490 24912 21496
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 20602 24900 20742
rect 25056 20602 25084 20946
rect 25148 20641 25176 21966
rect 25332 21690 25360 21966
rect 25516 21962 25544 22102
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25320 21684 25372 21690
rect 25320 21626 25372 21632
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25792 20942 25820 22374
rect 26252 21894 26280 22442
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26252 21690 26280 21830
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26344 21554 26372 22374
rect 26436 22098 26464 22374
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25134 20632 25190 20641
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 25044 20596 25096 20602
rect 26528 20618 26556 23990
rect 26804 23866 26832 24074
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26988 23338 27016 26522
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27080 24818 27108 26318
rect 27160 25220 27212 25226
rect 27160 25162 27212 25168
rect 27172 24886 27200 25162
rect 27160 24880 27212 24886
rect 27160 24822 27212 24828
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 27172 24070 27200 24686
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 26988 23310 27108 23338
rect 27172 23322 27200 24006
rect 26976 23248 27028 23254
rect 26976 23190 27028 23196
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26804 22778 26832 22918
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26620 21554 26648 22578
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26804 21690 26832 21966
rect 26988 21690 27016 23190
rect 26792 21684 26844 21690
rect 26792 21626 26844 21632
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26606 21448 26662 21457
rect 26662 21406 26740 21434
rect 26606 21383 26662 21392
rect 26528 20590 26648 20618
rect 25134 20567 25190 20576
rect 25044 20538 25096 20544
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 25056 19922 25084 20538
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24768 19712 24820 19718
rect 24320 18358 24348 19654
rect 24412 19638 24532 19666
rect 24768 19654 24820 19660
rect 24400 19304 24452 19310
rect 24504 19281 24532 19638
rect 24400 19246 24452 19252
rect 24490 19272 24546 19281
rect 24412 18426 24440 19246
rect 24490 19207 24546 19216
rect 24504 18834 24532 19207
rect 24780 18970 24808 19654
rect 24872 19310 24900 19790
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18970 24900 19110
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24596 18426 24624 18702
rect 24964 18426 24992 19654
rect 25148 19378 25176 20567
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19378 25268 19654
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25044 19304 25096 19310
rect 25332 19258 25360 19858
rect 25608 19446 25636 20334
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25044 19246 25096 19252
rect 25056 18902 25084 19246
rect 25148 19230 25360 19258
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 25148 18714 25176 19230
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25056 18686 25176 18714
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 24676 18284 24728 18290
rect 24952 18284 25004 18290
rect 24728 18244 24900 18272
rect 24676 18226 24728 18232
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24504 16114 24532 18022
rect 24872 17882 24900 18244
rect 25056 18272 25084 18686
rect 25332 18426 25360 18702
rect 25608 18426 25636 19110
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25004 18244 25084 18272
rect 24952 18226 25004 18232
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24964 17762 24992 18226
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24780 17734 24992 17762
rect 24780 17678 24808 17734
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24596 15570 24624 16390
rect 24964 16182 24992 16390
rect 25056 16250 25084 17478
rect 25148 17202 25176 18158
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24872 15706 24900 15914
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24412 14618 24440 14894
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24412 13530 24440 13806
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24412 12986 24440 13466
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12442 24348 12786
rect 24308 12436 24360 12442
rect 24504 12434 24532 14282
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24596 13841 24624 13874
rect 24582 13832 24638 13841
rect 24582 13767 24638 13776
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24504 12406 24624 12434
rect 24308 12378 24360 12384
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24136 10169 24164 10202
rect 24122 10160 24178 10169
rect 24122 10095 24178 10104
rect 24228 10062 24256 10950
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24044 9646 24164 9674
rect 24030 9208 24086 9217
rect 24030 9143 24032 9152
rect 24084 9143 24086 9152
rect 24032 9114 24084 9120
rect 23940 8560 23992 8566
rect 23940 8502 23992 8508
rect 23846 8392 23902 8401
rect 23846 8327 23902 8336
rect 23952 8294 23980 8502
rect 23860 8266 23980 8294
rect 23860 7886 23888 8266
rect 24136 8072 24164 9646
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 23952 8044 24164 8072
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23860 7546 23888 7822
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23846 7440 23902 7449
rect 23676 7398 23796 7426
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23400 6633 23428 6666
rect 23386 6624 23442 6633
rect 23386 6559 23442 6568
rect 23584 5914 23612 6802
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23768 5030 23796 7398
rect 23846 7375 23902 7384
rect 23860 7002 23888 7375
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23952 6905 23980 8044
rect 24228 7954 24256 8434
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 23938 6896 23994 6905
rect 23938 6831 23994 6840
rect 23952 6497 23980 6831
rect 23938 6488 23994 6497
rect 23938 6423 23994 6432
rect 24044 6322 24072 7890
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7041 24164 7686
rect 24320 7449 24348 12038
rect 24504 11393 24532 12038
rect 24490 11384 24546 11393
rect 24490 11319 24546 11328
rect 24400 11280 24452 11286
rect 24400 11222 24452 11228
rect 24412 8906 24440 11222
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24504 10810 24532 11086
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 10266 24532 10542
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24490 9072 24546 9081
rect 24596 9058 24624 12406
rect 24546 9030 24624 9058
rect 24490 9007 24546 9016
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24596 8634 24624 8910
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24412 8129 24440 8366
rect 24398 8120 24454 8129
rect 24596 8090 24624 8366
rect 24398 8055 24454 8064
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24688 7936 24716 13398
rect 24780 12646 24808 15302
rect 25148 15094 25176 17138
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25700 16114 25728 20334
rect 25792 20058 25820 20334
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 25976 20058 26004 20198
rect 26344 20058 26372 20198
rect 26528 20058 26556 20402
rect 26620 20398 26648 20590
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 25780 20052 25832 20058
rect 25780 19994 25832 20000
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26424 19780 26476 19786
rect 26424 19722 26476 19728
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25792 15994 25820 19382
rect 26056 19236 26108 19242
rect 26056 19178 26108 19184
rect 26068 17678 26096 19178
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26344 18970 26372 19110
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26436 18442 26464 19722
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26528 18834 26556 19110
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26436 18414 26556 18442
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26068 17202 26096 17614
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26252 16794 26280 17546
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26344 16726 26372 17750
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26436 17338 26464 17614
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26528 16998 26556 18414
rect 26620 17728 26648 20334
rect 26712 19378 26740 21406
rect 26976 21072 27028 21078
rect 26976 21014 27028 21020
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26896 20534 26924 20878
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26988 20058 27016 21014
rect 27080 20466 27108 23310
rect 27160 23316 27212 23322
rect 27160 23258 27212 23264
rect 27172 23118 27200 23258
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 26976 20052 27028 20058
rect 26976 19994 27028 20000
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26792 17740 26844 17746
rect 26620 17700 26740 17728
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 26620 16250 26648 17546
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 25608 15966 25820 15994
rect 25964 15972 26016 15978
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25608 15638 25636 15966
rect 25964 15914 26016 15920
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25792 15706 25820 15846
rect 25976 15706 26004 15914
rect 25780 15700 25832 15706
rect 25780 15642 25832 15648
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24964 13394 24992 14758
rect 25148 14482 25176 15030
rect 25792 15026 25820 15642
rect 26344 15570 26372 16050
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26436 15706 26464 15846
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26712 15570 26740 17700
rect 26792 17682 26844 17688
rect 26804 17082 26832 17682
rect 26896 17270 26924 18022
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 26988 17202 27016 19994
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19378 27108 19654
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27172 18290 27200 19858
rect 27264 19786 27292 26998
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27632 26586 27660 26862
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27724 26586 27752 26726
rect 27816 26586 27844 27338
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27620 26580 27672 26586
rect 27620 26522 27672 26528
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27712 26308 27764 26314
rect 27712 26250 27764 26256
rect 27724 25906 27752 26250
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27356 25498 27384 25638
rect 27908 25498 27936 26930
rect 28080 26512 28132 26518
rect 28080 26454 28132 26460
rect 27988 25696 28040 25702
rect 27988 25638 28040 25644
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 28000 25430 28028 25638
rect 27988 25424 28040 25430
rect 27988 25366 28040 25372
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27540 24410 27568 25230
rect 28000 24970 28028 25366
rect 27908 24942 28028 24970
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27908 24138 27936 24942
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 27896 24132 27948 24138
rect 27896 24074 27948 24080
rect 28000 23866 28028 24550
rect 28092 24138 28120 26454
rect 28184 25362 28212 27406
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 27033 28488 27270
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28446 27024 28502 27033
rect 28264 26988 28316 26994
rect 28446 26959 28502 26968
rect 28264 26930 28316 26936
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28184 24954 28212 25298
rect 28172 24948 28224 24954
rect 28172 24890 28224 24896
rect 28276 24682 28304 26930
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 28368 25906 28396 26726
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28552 25498 28580 26318
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28540 25492 28592 25498
rect 28540 25434 28592 25440
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28172 24608 28224 24614
rect 28172 24550 28224 24556
rect 28080 24132 28132 24138
rect 28080 24074 28132 24080
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27988 23180 28040 23186
rect 27988 23122 28040 23128
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27540 22098 27568 22918
rect 27724 22574 27752 23054
rect 27896 23044 27948 23050
rect 27896 22986 27948 22992
rect 27908 22778 27936 22986
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27896 22568 27948 22574
rect 27896 22510 27948 22516
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27448 20890 27476 21966
rect 27908 21962 27936 22510
rect 28000 22137 28028 23122
rect 28184 23050 28212 24550
rect 28264 24132 28316 24138
rect 28264 24074 28316 24080
rect 28276 23526 28304 24074
rect 28368 23866 28396 24754
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28276 23254 28304 23462
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 27986 22128 28042 22137
rect 27986 22063 28042 22072
rect 27896 21956 27948 21962
rect 27896 21898 27948 21904
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 27356 20862 27476 20890
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27356 20058 27384 20862
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27448 20466 27476 20742
rect 27540 20602 27568 20878
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27632 20466 27660 20742
rect 27724 20602 27752 20810
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27712 20392 27764 20398
rect 27764 20352 27844 20380
rect 27712 20334 27764 20340
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 27540 19854 27568 20198
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27540 18834 27568 19314
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26804 17054 26924 17082
rect 26896 16522 26924 17054
rect 27172 16658 27200 18226
rect 27264 17882 27292 18566
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27436 17604 27488 17610
rect 27436 17546 27488 17552
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26884 16516 26936 16522
rect 26884 16458 26936 16464
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25884 14618 25912 14962
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 13977 25268 14282
rect 25226 13968 25282 13977
rect 25226 13903 25228 13912
rect 25280 13903 25282 13912
rect 25228 13874 25280 13880
rect 25332 13734 25360 14350
rect 26252 14090 26280 15302
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26620 14618 26648 14962
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26424 14340 26476 14346
rect 26424 14282 26476 14288
rect 26068 14062 26280 14090
rect 26068 13954 26096 14062
rect 25792 13938 26096 13954
rect 25780 13932 26096 13938
rect 25832 13926 26096 13932
rect 25780 13874 25832 13880
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25056 13530 25084 13670
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 25516 13138 25544 13466
rect 25516 13110 25636 13138
rect 24952 12776 25004 12782
rect 24872 12724 24952 12730
rect 24872 12718 25004 12724
rect 24872 12702 24992 12718
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24780 11150 24808 12582
rect 24872 11558 24900 12702
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25608 12306 25636 13110
rect 25792 12918 25820 13670
rect 25976 13394 26004 13670
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25136 12164 25188 12170
rect 25136 12106 25188 12112
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24872 11218 24900 11494
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24872 10606 24900 11154
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 25056 10810 25084 10950
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 24952 10736 25004 10742
rect 24952 10678 25004 10684
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24780 9081 24808 10474
rect 24872 9654 24900 10542
rect 24964 10010 24992 10678
rect 25056 10130 25084 10746
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25148 10010 25176 12106
rect 25516 11540 25544 12174
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25516 11512 25636 11540
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25608 11354 25636 11512
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25226 11248 25282 11257
rect 25226 11183 25282 11192
rect 25240 10674 25268 11183
rect 25976 11121 26004 12038
rect 25962 11112 26018 11121
rect 25962 11047 26018 11056
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 24964 9982 25084 10010
rect 25148 9982 25452 10010
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9722 24992 9862
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24766 9072 24822 9081
rect 24872 9042 24900 9590
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24766 9007 24822 9016
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24780 8566 24808 8910
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24872 8566 24900 8842
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24766 8392 24822 8401
rect 24766 8327 24822 8336
rect 24780 8090 24808 8327
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24964 7954 24992 9454
rect 25056 9382 25084 9982
rect 25424 9926 25452 9982
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25148 9178 25176 9862
rect 25964 9648 26016 9654
rect 25792 9608 25964 9636
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8566 25084 8774
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 25792 8430 25820 9608
rect 25964 9590 26016 9596
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25134 8120 25190 8129
rect 25261 8123 25569 8132
rect 25134 8055 25190 8064
rect 25320 8084 25372 8090
rect 24952 7948 25004 7954
rect 24688 7908 24900 7936
rect 24492 7880 24544 7886
rect 24544 7840 24808 7868
rect 24492 7822 24544 7828
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24306 7440 24362 7449
rect 24306 7375 24362 7384
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24306 7304 24362 7313
rect 24122 7032 24178 7041
rect 24122 6967 24178 6976
rect 24228 6798 24256 7278
rect 24306 7239 24362 7248
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23952 5370 23980 6258
rect 24044 6118 24072 6258
rect 24032 6112 24084 6118
rect 24216 6112 24268 6118
rect 24084 6072 24164 6100
rect 24032 6054 24084 6060
rect 24136 5710 24164 6072
rect 24216 6054 24268 6060
rect 24228 5914 24256 6054
rect 24320 5930 24348 7239
rect 24504 6746 24532 7482
rect 24582 7440 24638 7449
rect 24582 7375 24638 7384
rect 24412 6718 24532 6746
rect 24412 6390 24440 6718
rect 24490 6488 24546 6497
rect 24490 6423 24546 6432
rect 24504 6390 24532 6423
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24216 5908 24268 5914
rect 24320 5902 24532 5930
rect 24216 5850 24268 5856
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23676 4758 23704 4966
rect 23860 4758 23888 5306
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23848 4752 23900 4758
rect 23848 4694 23900 4700
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23386 4176 23442 4185
rect 23386 4111 23388 4120
rect 23440 4111 23442 4120
rect 23388 4082 23440 4088
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23400 3754 23428 3878
rect 23400 3726 23520 3754
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 23400 2938 23428 3538
rect 23308 2922 23428 2938
rect 23296 2916 23428 2922
rect 23348 2910 23428 2916
rect 23296 2858 23348 2864
rect 23308 2666 23336 2858
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23216 2638 23336 2666
rect 22558 2479 22614 2488
rect 22836 2508 22888 2514
rect 21916 2450 21968 2456
rect 22836 2450 22888 2456
rect 23112 2508 23164 2514
rect 23112 2450 23164 2456
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21548 2372 21600 2378
rect 21548 2314 21600 2320
rect 19800 2032 19852 2038
rect 19800 1974 19852 1980
rect 21560 1970 21588 2314
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 23216 1970 23244 2638
rect 23400 2530 23428 2790
rect 23492 2564 23520 3726
rect 23584 2774 23612 4490
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23676 3670 23704 4014
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23676 3058 23704 3606
rect 23768 3194 23796 4626
rect 24044 4162 24072 5646
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24228 4706 24256 4966
rect 24320 4826 24348 5782
rect 24398 5264 24454 5273
rect 24398 5199 24400 5208
rect 24452 5199 24454 5208
rect 24400 5170 24452 5176
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24228 4678 24348 4706
rect 24320 4554 24348 4678
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 24412 4282 24440 4558
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 23952 4134 24072 4162
rect 23952 3670 23980 4134
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23860 3194 23888 3538
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23952 3074 23980 3606
rect 24044 3097 24072 4014
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23768 3046 23980 3074
rect 24030 3088 24086 3097
rect 23584 2746 23704 2774
rect 23572 2576 23624 2582
rect 23492 2536 23572 2564
rect 23308 2502 23428 2530
rect 23572 2518 23624 2524
rect 23308 2446 23336 2502
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 23400 2106 23428 2314
rect 23676 2310 23704 2746
rect 23768 2446 23796 3046
rect 24030 3023 24086 3032
rect 23846 2680 23902 2689
rect 23846 2615 23902 2624
rect 23860 2446 23888 2615
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23572 2304 23624 2310
rect 23572 2246 23624 2252
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23492 2106 23520 2246
rect 23584 2106 23612 2246
rect 23388 2100 23440 2106
rect 23388 2042 23440 2048
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 21548 1964 21600 1970
rect 21548 1906 21600 1912
rect 23204 1964 23256 1970
rect 23204 1906 23256 1912
rect 18788 1760 18840 1766
rect 18788 1702 18840 1708
rect 24228 1698 24256 4014
rect 24320 3738 24348 4218
rect 24412 3738 24440 4218
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24504 3534 24532 5902
rect 24596 4758 24624 7375
rect 24780 6866 24808 7840
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24872 6798 24900 7908
rect 24952 7890 25004 7896
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24688 5710 24716 6598
rect 24964 6390 24992 7890
rect 25148 7528 25176 8055
rect 25320 8026 25372 8032
rect 25148 7500 25268 7528
rect 25240 7188 25268 7500
rect 25332 7206 25360 8026
rect 25976 7886 26004 8230
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25424 7546 25820 7562
rect 25424 7540 25832 7546
rect 25424 7534 25780 7540
rect 25424 7342 25452 7534
rect 25780 7482 25832 7488
rect 25792 7410 25820 7482
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25148 7160 25268 7188
rect 25320 7200 25372 7206
rect 25148 6866 25176 7160
rect 25320 7142 25372 7148
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25042 6624 25098 6633
rect 25042 6559 25098 6568
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 25056 6186 25084 6559
rect 25240 6458 25268 6666
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 6180 25096 6186
rect 25044 6122 25096 6128
rect 25148 5914 25176 6190
rect 25424 6186 25452 6666
rect 25700 6633 25728 7346
rect 26068 7290 26096 13926
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26146 13832 26202 13841
rect 26146 13767 26202 13776
rect 26160 13734 26188 13767
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26252 13326 26280 13874
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26252 12714 26280 13262
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26252 12170 26280 12650
rect 26344 12442 26372 13874
rect 26436 13530 26464 14282
rect 26608 13728 26660 13734
rect 26608 13670 26660 13676
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26528 13002 26556 13126
rect 26436 12974 26556 13002
rect 26620 12986 26648 13670
rect 26804 13546 26832 15846
rect 26896 14940 26924 16458
rect 27172 16114 27200 16594
rect 27448 16232 27476 17546
rect 27632 17218 27660 19722
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27724 19310 27752 19654
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27816 19122 27844 20352
rect 27908 19990 27936 20878
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 27908 19854 27936 19926
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27908 19446 27936 19790
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 27896 19440 27948 19446
rect 27896 19382 27948 19388
rect 27540 17202 27660 17218
rect 27528 17196 27660 17202
rect 27580 17190 27660 17196
rect 27724 19094 27844 19122
rect 27528 17138 27580 17144
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27448 16204 27568 16232
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 26988 15094 27016 16050
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 27080 15638 27108 15982
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 27172 15008 27200 16050
rect 27356 15366 27384 16050
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27252 15020 27304 15026
rect 27172 14980 27252 15008
rect 27252 14962 27304 14968
rect 26896 14912 27200 14940
rect 26976 14816 27028 14822
rect 26976 14758 27028 14764
rect 26988 14618 27016 14758
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 27066 13968 27122 13977
rect 27066 13903 27068 13912
rect 27120 13903 27122 13912
rect 27068 13874 27120 13880
rect 26712 13518 26832 13546
rect 26608 12980 26660 12986
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26240 12164 26292 12170
rect 26240 12106 26292 12112
rect 26436 11830 26464 12974
rect 26608 12922 26660 12928
rect 26712 12730 26740 13518
rect 26620 12702 26740 12730
rect 26804 13394 27016 13410
rect 26804 13388 27028 13394
rect 26804 13382 26976 13388
rect 26620 11937 26648 12702
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12306 26740 12582
rect 26804 12306 26832 13382
rect 26976 13330 27028 13336
rect 27080 13274 27108 13874
rect 26896 13246 27108 13274
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 26606 11928 26662 11937
rect 26606 11863 26662 11872
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 26804 11642 26832 12242
rect 26712 11614 26832 11642
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11286 26648 11494
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26712 11132 26740 11614
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 26620 11104 26740 11132
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26160 10810 26188 11018
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26238 10160 26294 10169
rect 26148 10124 26200 10130
rect 26238 10095 26240 10104
rect 26148 10066 26200 10072
rect 26292 10095 26294 10104
rect 26240 10066 26292 10072
rect 26160 8294 26188 10066
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26252 9489 26280 9522
rect 26238 9480 26294 9489
rect 26238 9415 26294 9424
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26344 8634 26372 9318
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26436 8514 26464 10610
rect 26620 9625 26648 11104
rect 26804 10742 26832 11494
rect 26896 11150 26924 13246
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 27080 11898 27108 12718
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26884 10668 26936 10674
rect 26884 10610 26936 10616
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26712 10130 26740 10406
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26712 9722 26740 10066
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26606 9616 26662 9625
rect 26606 9551 26662 9560
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26436 8486 26556 8514
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 8090 26188 8230
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26422 7984 26478 7993
rect 26528 7954 26556 8486
rect 26422 7919 26478 7928
rect 26516 7948 26568 7954
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26160 7410 26188 7686
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 25976 7262 26096 7290
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25686 6624 25742 6633
rect 25686 6559 25742 6568
rect 25780 6384 25832 6390
rect 25780 6326 25832 6332
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24780 4282 24808 5170
rect 24872 4622 24900 5578
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25056 5302 25084 5510
rect 25148 5370 25176 5646
rect 25516 5370 25544 5850
rect 25792 5778 25820 6326
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25504 5364 25556 5370
rect 25504 5306 25556 5312
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4622 24992 4966
rect 25148 4826 25176 5306
rect 25320 5160 25372 5166
rect 25318 5128 25320 5137
rect 25372 5128 25374 5137
rect 25318 5063 25374 5072
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 25504 4616 25556 4622
rect 25504 4558 25556 4564
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 25424 4146 25452 4422
rect 25516 4214 25544 4558
rect 25504 4208 25556 4214
rect 25504 4150 25556 4156
rect 25136 4140 25188 4146
rect 25136 4082 25188 4088
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 24860 4072 24912 4078
rect 25148 4026 25176 4082
rect 24860 4014 24912 4020
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24584 3528 24636 3534
rect 24872 3505 24900 4014
rect 24964 3998 25176 4026
rect 24584 3470 24636 3476
rect 24858 3496 24914 3505
rect 24412 2961 24440 3470
rect 24398 2952 24454 2961
rect 24398 2887 24454 2896
rect 24596 2650 24624 3470
rect 24676 3460 24728 3466
rect 24858 3431 24914 3440
rect 24676 3402 24728 3408
rect 24688 2854 24716 3402
rect 24872 3194 24900 3431
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24780 2378 24808 2518
rect 24964 2446 24992 3998
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25148 3058 25176 3878
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25608 2650 25636 5646
rect 25700 4146 25728 5646
rect 25780 5092 25832 5098
rect 25780 5034 25832 5040
rect 25792 4826 25820 5034
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25792 3913 25820 4014
rect 25778 3904 25834 3913
rect 25778 3839 25834 3848
rect 25884 3738 25912 7142
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25870 3632 25926 3641
rect 25700 3398 25728 3606
rect 25870 3567 25872 3576
rect 25924 3567 25926 3576
rect 25872 3538 25924 3544
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25700 2514 25728 3334
rect 25976 2774 26004 7262
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 26068 6390 26096 7142
rect 26056 6384 26108 6390
rect 26056 6326 26108 6332
rect 26160 5710 26188 7346
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26252 6390 26280 6938
rect 26332 6656 26384 6662
rect 26330 6624 26332 6633
rect 26384 6624 26386 6633
rect 26330 6559 26386 6568
rect 26436 6474 26464 7919
rect 26516 7890 26568 7896
rect 26620 7834 26648 9114
rect 26712 8276 26740 9318
rect 26804 8945 26832 9522
rect 26896 9382 26924 10610
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26790 8936 26846 8945
rect 26790 8871 26846 8880
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26896 8430 26924 8774
rect 26988 8498 27016 11698
rect 27172 10674 27200 14912
rect 27448 14618 27476 16050
rect 27540 15026 27568 16204
rect 27632 15570 27660 16934
rect 27724 16046 27752 19094
rect 28000 18834 28028 19654
rect 28092 19310 28120 21830
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 28092 18426 28120 18566
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 27896 18216 27948 18222
rect 27896 18158 27948 18164
rect 27802 17232 27858 17241
rect 27802 17167 27858 17176
rect 27816 16794 27844 17167
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27816 15570 27844 16390
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27804 15564 27856 15570
rect 27804 15506 27856 15512
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27724 15162 27752 15302
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27620 14952 27672 14958
rect 27620 14894 27672 14900
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27356 13870 27384 14486
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27264 12986 27292 13466
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27448 11762 27476 12582
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27344 11688 27396 11694
rect 27540 11642 27568 14418
rect 27632 14006 27660 14894
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 27724 12782 27752 15098
rect 27816 14482 27844 15302
rect 27908 15162 27936 18158
rect 28092 17134 28120 18362
rect 28080 17128 28132 17134
rect 28080 17070 28132 17076
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 28092 15706 28120 15846
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 28184 15366 28212 19246
rect 28368 18290 28396 21830
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28368 17338 28396 17478
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 27816 12434 27844 14010
rect 28092 13938 28120 14758
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28184 13870 28212 14350
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27724 12406 27844 12434
rect 27724 12306 27752 12406
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27344 11630 27396 11636
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27264 10674 27292 11494
rect 27356 10810 27384 11630
rect 27448 11614 27568 11642
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27448 10538 27476 11614
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27540 10606 27568 10950
rect 27528 10600 27580 10606
rect 27526 10568 27528 10577
rect 27580 10568 27582 10577
rect 27436 10532 27488 10538
rect 27526 10503 27582 10512
rect 27436 10474 27488 10480
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27080 9586 27108 10202
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27080 9178 27108 9318
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 27066 8528 27122 8537
rect 26976 8492 27028 8498
rect 27066 8463 27122 8472
rect 26976 8434 27028 8440
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26712 8248 26924 8276
rect 26344 6446 26464 6474
rect 26528 7806 26648 7834
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26238 6216 26294 6225
rect 26238 6151 26294 6160
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 26252 5234 26280 6151
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26148 4616 26200 4622
rect 26054 4584 26110 4593
rect 26148 4558 26200 4564
rect 26054 4519 26110 4528
rect 26068 3602 26096 4519
rect 26160 4078 26188 4558
rect 26252 4486 26280 5170
rect 26344 4622 26372 6446
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26436 5234 26464 5714
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26240 4480 26292 4486
rect 26528 4434 26556 7806
rect 26606 7712 26662 7721
rect 26606 7647 26662 7656
rect 26620 7002 26648 7647
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26620 6866 26648 6938
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26240 4422 26292 4428
rect 26344 4406 26556 4434
rect 26344 4078 26372 4406
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26332 4072 26384 4078
rect 26516 4072 26568 4078
rect 26332 4014 26384 4020
rect 26514 4040 26516 4049
rect 26568 4040 26570 4049
rect 26160 3738 26188 4014
rect 26514 3975 26570 3984
rect 26620 3738 26648 6394
rect 26712 5370 26740 7822
rect 26804 5914 26832 7822
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26896 5302 26924 8248
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 27080 4978 27108 8463
rect 27250 7848 27306 7857
rect 27250 7783 27306 7792
rect 27264 6798 27292 7783
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27250 5536 27306 5545
rect 27250 5471 27306 5480
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 26988 4950 27108 4978
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26988 4570 27016 4950
rect 27066 4720 27122 4729
rect 27066 4655 27068 4664
rect 27120 4655 27122 4664
rect 27068 4626 27120 4632
rect 26804 4486 26832 4558
rect 26988 4542 27108 4570
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26804 4146 26832 4422
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26804 3738 26832 4082
rect 26988 3913 27016 4082
rect 26974 3904 27030 3913
rect 26974 3839 27030 3848
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 25976 2746 26096 2774
rect 26068 2650 26096 2746
rect 26712 2650 26740 2994
rect 27080 2836 27108 4542
rect 27172 3602 27200 5170
rect 27264 4690 27292 5471
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27356 3738 27384 9454
rect 27632 9178 27660 9862
rect 27724 9722 27752 10406
rect 27908 10146 27936 13194
rect 28000 12374 28028 13806
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12986 28120 13126
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 28092 12434 28120 12922
rect 28092 12406 28212 12434
rect 27988 12368 28040 12374
rect 27988 12310 28040 12316
rect 28000 11762 28028 12310
rect 28184 11898 28212 12406
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28276 11778 28304 16390
rect 28368 15706 28396 16458
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 28368 14074 28396 15370
rect 28460 15162 28488 20742
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28552 16250 28580 18702
rect 28644 16658 28672 21286
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 28540 14816 28592 14822
rect 28540 14758 28592 14764
rect 28448 14340 28500 14346
rect 28448 14282 28500 14288
rect 28356 14068 28408 14074
rect 28356 14010 28408 14016
rect 28460 11898 28488 14282
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 28184 11750 28304 11778
rect 28552 11762 28580 14758
rect 28644 13462 28672 16594
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28630 12336 28686 12345
rect 28630 12271 28686 12280
rect 28540 11756 28592 11762
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 28092 10282 28120 11494
rect 28184 11150 28212 11750
rect 28540 11698 28592 11704
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28276 10674 28304 11154
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28092 10254 28212 10282
rect 27908 10118 28120 10146
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27804 9920 27856 9926
rect 27804 9862 27856 9868
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27816 8974 27844 9862
rect 28000 9722 28028 9998
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27436 8016 27488 8022
rect 27436 7958 27488 7964
rect 27448 7410 27476 7958
rect 27436 7404 27488 7410
rect 27436 7346 27488 7352
rect 27540 6934 27568 8230
rect 27528 6928 27580 6934
rect 27528 6870 27580 6876
rect 27632 6202 27660 8910
rect 27908 8430 27936 9590
rect 27988 9444 28040 9450
rect 27988 9386 28040 9392
rect 28000 8430 28028 9386
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 28092 8090 28120 10118
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 28184 8022 28212 10254
rect 28264 10124 28316 10130
rect 28264 10066 28316 10072
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 28276 7290 28304 10066
rect 28540 9988 28592 9994
rect 28540 9930 28592 9936
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 9722 28488 9862
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 28368 8634 28396 8774
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28184 7262 28304 7290
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27908 6798 27936 7142
rect 27896 6792 27948 6798
rect 27988 6792 28040 6798
rect 27896 6734 27948 6740
rect 27986 6760 27988 6769
rect 28040 6760 28042 6769
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27816 6254 27844 6598
rect 27908 6458 27936 6734
rect 27986 6695 28042 6704
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27804 6248 27856 6254
rect 27632 6174 27752 6202
rect 27804 6190 27856 6196
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27632 5914 27660 6054
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27540 5302 27568 5578
rect 27618 5400 27674 5409
rect 27618 5335 27674 5344
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 27632 4690 27660 5335
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27632 4282 27660 4490
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27724 4146 27752 6174
rect 27816 4826 27844 6190
rect 28184 5574 28212 7262
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 28276 6497 28304 7142
rect 28262 6488 28318 6497
rect 28262 6423 28318 6432
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 27172 3194 27200 3538
rect 27988 3460 28040 3466
rect 27988 3402 28040 3408
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27252 3052 27304 3058
rect 27252 2994 27304 3000
rect 27160 2848 27212 2854
rect 27080 2808 27160 2836
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 27080 2514 27108 2808
rect 27160 2790 27212 2796
rect 27264 2650 27292 2994
rect 28000 2650 28028 3402
rect 27252 2644 27304 2650
rect 27252 2586 27304 2592
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 28368 2446 28396 7686
rect 28552 5914 28580 9930
rect 28644 7886 28672 12271
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 28540 5908 28592 5914
rect 28540 5850 28592 5856
rect 28538 5808 28594 5817
rect 28538 5743 28594 5752
rect 28552 5370 28580 5743
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 28552 2514 28580 5306
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 28540 2508 28592 2514
rect 28540 2450 28592 2456
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 24216 1692 24268 1698
rect 24216 1634 24268 1640
rect 11348 734 11652 762
rect 18694 0 18750 800
rect 26146 0 26202 800
<< via2 >>
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 938 27276 940 27296
rect 940 27276 992 27296
rect 992 27276 994 27296
rect 938 27240 994 27276
rect 2594 27004 2596 27024
rect 2596 27004 2648 27024
rect 2648 27004 2650 27024
rect 2594 26968 2650 27004
rect 3790 26832 3846 26888
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 3422 25780 3424 25800
rect 3424 25780 3476 25800
rect 3476 25780 3478 25800
rect 3422 25744 3478 25780
rect 1582 23704 1638 23760
rect 1950 24928 2006 24984
rect 2962 20304 3018 20360
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 1306 16632 1362 16688
rect 5262 22092 5318 22128
rect 5262 22072 5264 22092
rect 5264 22072 5316 22092
rect 5316 22072 5318 22092
rect 6826 27376 6882 27432
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 6366 26288 6422 26344
rect 6366 24928 6422 24984
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 938 13096 994 13152
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4526 15272 4582 15328
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 5538 21428 5540 21448
rect 5540 21428 5592 21448
rect 5592 21428 5594 21448
rect 5538 21392 5594 21428
rect 7286 26324 7288 26344
rect 7288 26324 7340 26344
rect 7340 26324 7342 26344
rect 7286 26288 7342 26324
rect 5998 21972 6000 21992
rect 6000 21972 6052 21992
rect 6052 21972 6054 21992
rect 5998 21936 6054 21972
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 8482 25764 8538 25800
rect 8482 25744 8484 25764
rect 8484 25744 8536 25764
rect 8536 25744 8538 25764
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 10046 26968 10102 27024
rect 10230 27376 10286 27432
rect 9862 26016 9918 26072
rect 10046 26852 10102 26888
rect 10046 26832 10048 26852
rect 10048 26832 10100 26852
rect 10100 26832 10102 26852
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 8298 22516 8300 22536
rect 8300 22516 8352 22536
rect 8352 22516 8354 22536
rect 8298 22480 8354 22516
rect 8114 22208 8170 22264
rect 8206 22072 8262 22128
rect 7286 19896 7342 19952
rect 5446 17992 5502 18048
rect 6366 17856 6422 17912
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 8390 19760 8446 19816
rect 8666 22208 8722 22264
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 5446 17176 5502 17232
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 2962 11192 3018 11248
rect 2686 11092 2688 11112
rect 2688 11092 2740 11112
rect 2740 11092 2742 11112
rect 2686 11056 2742 11092
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 4618 11872 4674 11928
rect 5078 12724 5080 12744
rect 5080 12724 5132 12744
rect 5132 12724 5134 12744
rect 5078 12688 5134 12724
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 1398 9560 1454 9616
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 5354 11736 5410 11792
rect 6826 11600 6882 11656
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 5170 6840 5226 6896
rect 1858 3476 1860 3496
rect 1860 3476 1912 3496
rect 1912 3476 1914 3496
rect 1858 3440 1914 3476
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 2502 3304 2558 3360
rect 3790 3304 3846 3360
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 9678 22888 9734 22944
rect 9494 22516 9496 22536
rect 9496 22516 9548 22536
rect 9548 22516 9550 22536
rect 9494 22480 9550 22516
rect 8850 22092 8906 22128
rect 8850 22072 8852 22092
rect 8852 22072 8904 22092
rect 8904 22072 8906 22092
rect 9126 21392 9182 21448
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 8022 13932 8078 13968
rect 8022 13912 8024 13932
rect 8024 13912 8076 13932
rect 8076 13912 8078 13932
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 8482 13912 8538 13968
rect 9862 22108 9864 22128
rect 9864 22108 9916 22128
rect 9916 22108 9918 22128
rect 9862 22072 9918 22108
rect 10046 21936 10102 21992
rect 10046 20984 10102 21040
rect 9770 20304 9826 20360
rect 12346 26288 12402 26344
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 13910 26288 13966 26344
rect 14370 26036 14426 26072
rect 14370 26016 14372 26036
rect 14372 26016 14424 26036
rect 14424 26016 14426 26036
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 10414 21956 10470 21992
rect 10414 21936 10416 21956
rect 10416 21936 10468 21956
rect 10468 21936 10470 21956
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 10598 20304 10654 20360
rect 10414 19916 10470 19952
rect 10414 19896 10416 19916
rect 10416 19896 10468 19916
rect 10468 19896 10470 19916
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11334 19780 11390 19816
rect 11334 19760 11336 19780
rect 11336 19760 11388 19780
rect 11388 19760 11390 19780
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11058 17856 11114 17912
rect 9586 12416 9642 12472
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 5630 7520 5686 7576
rect 6366 7520 6422 7576
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 8390 11192 8446 11248
rect 8482 11092 8484 11112
rect 8484 11092 8536 11112
rect 8536 11092 8538 11112
rect 8482 11056 8538 11092
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 5170 3460 5226 3496
rect 5170 3440 5172 3460
rect 5172 3440 5224 3460
rect 5224 3440 5226 3460
rect 5354 4120 5410 4176
rect 4342 2916 4398 2952
rect 4342 2896 4344 2916
rect 4344 2896 4396 2916
rect 4396 2896 4398 2916
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 6274 3984 6330 4040
rect 6550 3712 6606 3768
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 10230 14320 10286 14376
rect 9862 12724 9864 12744
rect 9864 12724 9916 12744
rect 9916 12724 9918 12744
rect 9862 12688 9918 12724
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 9586 7964 9588 7984
rect 9588 7964 9640 7984
rect 9640 7964 9642 7984
rect 9586 7928 9642 7964
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11242 12416 11298 12472
rect 11058 11636 11060 11656
rect 11060 11636 11112 11656
rect 11112 11636 11114 11656
rect 11058 11600 11114 11636
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11518 10648 11574 10704
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 10046 5772 10102 5808
rect 10046 5752 10048 5772
rect 10048 5752 10100 5772
rect 10100 5752 10102 5772
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 10138 5072 10194 5128
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11886 7948 11942 7984
rect 11886 7928 11888 7948
rect 11888 7928 11940 7948
rect 11940 7928 11942 7948
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14554 22888 14610 22944
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 20534 25780 20536 25800
rect 20536 25780 20588 25800
rect 20588 25780 20590 25800
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 20534 25744 20590 25780
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 15198 20984 15254 21040
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 22742 26868 22744 26888
rect 22744 26868 22796 26888
rect 22796 26868 22798 26888
rect 22742 26832 22798 26868
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14554 14320 14610 14376
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 6734 3440 6790 3496
rect 8114 3984 8170 4040
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 9126 3712 9182 3768
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 6274 2488 6330 2544
rect 5998 2352 6054 2408
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 14646 6840 14702 6896
rect 14094 5208 14150 5264
rect 12346 3440 12402 3496
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 15750 20576 15806 20632
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18786 22072 18842 22128
rect 16486 21428 16488 21448
rect 16488 21428 16540 21448
rect 16540 21428 16542 21448
rect 16486 21392 16542 21428
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 15106 7792 15162 7848
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14738 6160 14794 6216
rect 14370 5772 14426 5808
rect 14370 5752 14372 5772
rect 14372 5752 14424 5772
rect 14424 5752 14426 5772
rect 14278 5108 14280 5128
rect 14280 5108 14332 5128
rect 14332 5108 14334 5128
rect 14278 5072 14334 5108
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 19890 22208 19946 22264
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 17130 15408 17186 15464
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 17774 11736 17830 11792
rect 17498 11600 17554 11656
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 16210 8880 16266 8936
rect 15842 5480 15898 5536
rect 15658 3984 15714 4040
rect 16670 6976 16726 7032
rect 16578 6724 16634 6760
rect 16578 6704 16580 6724
rect 16580 6704 16632 6724
rect 16632 6704 16634 6724
rect 16670 6568 16726 6624
rect 15934 3304 15990 3360
rect 16302 3984 16358 4040
rect 16762 3576 16818 3632
rect 17406 7384 17462 7440
rect 17406 4528 17462 4584
rect 17314 3440 17370 3496
rect 16394 3304 16450 3360
rect 15750 3032 15806 3088
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 17590 8336 17646 8392
rect 17590 6860 17646 6896
rect 17590 6840 17592 6860
rect 17592 6840 17644 6860
rect 17644 6840 17646 6860
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21914 22208 21970 22264
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 20994 19372 21050 19408
rect 20994 19352 20996 19372
rect 20996 19352 21048 19372
rect 21048 19352 21050 19372
rect 21362 20712 21418 20768
rect 21086 19216 21142 19272
rect 19154 15408 19210 15464
rect 20442 17196 20498 17232
rect 20442 17176 20444 17196
rect 20444 17176 20496 17196
rect 20496 17176 20498 17196
rect 20626 16652 20682 16688
rect 20626 16632 20628 16652
rect 20628 16632 20680 16652
rect 20680 16632 20682 16652
rect 20534 16088 20590 16144
rect 19798 12280 19854 12336
rect 19430 11212 19486 11248
rect 19430 11192 19432 11212
rect 19432 11192 19484 11212
rect 19484 11192 19486 11212
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18510 6568 18566 6624
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18326 5752 18382 5808
rect 17774 5072 17830 5128
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18786 5072 18842 5128
rect 18694 3848 18750 3904
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 18970 6976 19026 7032
rect 19430 9288 19486 9344
rect 19614 9152 19670 9208
rect 19062 6432 19118 6488
rect 18970 5072 19026 5128
rect 19338 4936 19394 4992
rect 19614 7112 19670 7168
rect 19614 6432 19670 6488
rect 20074 9460 20076 9480
rect 20076 9460 20128 9480
rect 20128 9460 20130 9480
rect 20074 9424 20130 9460
rect 20994 16088 21050 16144
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21454 19372 21510 19408
rect 21454 19352 21456 19372
rect 21456 19352 21508 19372
rect 21508 19352 21510 19372
rect 20074 9016 20130 9072
rect 20074 8084 20130 8120
rect 20074 8064 20076 8084
rect 20076 8064 20128 8084
rect 20128 8064 20130 8084
rect 20350 9580 20406 9616
rect 20350 9560 20352 9580
rect 20352 9560 20404 9580
rect 20404 9560 20406 9580
rect 20442 8608 20498 8664
rect 20074 4800 20130 4856
rect 20902 9560 20958 9616
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 25686 26868 25688 26888
rect 25688 26868 25740 26888
rect 25740 26868 25742 26888
rect 25686 26832 25742 26868
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 22282 20596 22338 20632
rect 22282 20576 22284 20596
rect 22284 20576 22336 20596
rect 22336 20576 22338 20596
rect 22742 21392 22798 21448
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21362 10140 21364 10160
rect 21364 10140 21416 10160
rect 21416 10140 21418 10160
rect 21362 10104 21418 10140
rect 21086 8472 21142 8528
rect 21270 9580 21326 9616
rect 21270 9560 21272 9580
rect 21272 9560 21324 9580
rect 21324 9560 21326 9580
rect 21270 8336 21326 8392
rect 20718 5888 20774 5944
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 22190 10512 22246 10568
rect 21730 10124 21786 10160
rect 21730 10104 21732 10124
rect 21732 10104 21784 10124
rect 21784 10104 21786 10124
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 21822 9560 21878 9616
rect 21730 9152 21786 9208
rect 22282 9152 22338 9208
rect 21454 8064 21510 8120
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 21270 6568 21326 6624
rect 21546 5752 21602 5808
rect 21454 5480 21510 5536
rect 22006 6976 22062 7032
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 23202 16632 23258 16688
rect 22558 7520 22614 7576
rect 24030 11872 24086 11928
rect 23294 9288 23350 9344
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 21914 4800 21970 4856
rect 22190 4936 22246 4992
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 20994 3576 21050 3632
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21914 2624 21970 2680
rect 22834 6160 22890 6216
rect 22926 3848 22982 3904
rect 22558 2488 22614 2544
rect 23386 7656 23442 7712
rect 23846 9016 23902 9072
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25870 25744 25926 25800
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25134 20576 25190 20632
rect 26606 21392 26662 21448
rect 24490 19216 24546 19272
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 24582 13776 24638 13832
rect 24122 10104 24178 10160
rect 24030 9172 24086 9208
rect 24030 9152 24032 9172
rect 24032 9152 24084 9172
rect 24084 9152 24086 9172
rect 23846 8336 23902 8392
rect 23386 6568 23442 6624
rect 23846 7384 23902 7440
rect 23938 6840 23994 6896
rect 23938 6432 23994 6488
rect 24490 11328 24546 11384
rect 24490 9016 24546 9072
rect 24398 8064 24454 8120
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28446 26968 28502 27024
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 27986 22072 28042 22128
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25226 13932 25282 13968
rect 25226 13912 25228 13932
rect 25228 13912 25280 13932
rect 25280 13912 25282 13932
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 25226 11192 25282 11248
rect 25962 11056 26018 11112
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 24766 9016 24822 9072
rect 24766 8336 24822 8392
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25134 8064 25190 8120
rect 24306 7384 24362 7440
rect 24122 6976 24178 7032
rect 24306 7248 24362 7304
rect 24582 7384 24638 7440
rect 24490 6432 24546 6488
rect 23386 4140 23442 4176
rect 23386 4120 23388 4140
rect 23388 4120 23440 4140
rect 23440 4120 23442 4140
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 24398 5228 24454 5264
rect 24398 5208 24400 5228
rect 24400 5208 24452 5228
rect 24452 5208 24454 5228
rect 24030 3032 24086 3088
rect 23846 2624 23902 2680
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25042 6568 25098 6624
rect 26146 13776 26202 13832
rect 27066 13932 27122 13968
rect 27066 13912 27068 13932
rect 27068 13912 27120 13932
rect 27120 13912 27122 13932
rect 26606 11872 26662 11928
rect 26238 10124 26294 10160
rect 26238 10104 26240 10124
rect 26240 10104 26292 10124
rect 26292 10104 26294 10124
rect 26238 9424 26294 9480
rect 26606 9560 26662 9616
rect 26422 7928 26478 7984
rect 25686 6568 25742 6624
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25318 5108 25320 5128
rect 25320 5108 25372 5128
rect 25372 5108 25374 5128
rect 25318 5072 25374 5108
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 24398 2896 24454 2952
rect 24858 3440 24914 3496
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 25778 3848 25834 3904
rect 25870 3596 25926 3632
rect 25870 3576 25872 3596
rect 25872 3576 25924 3596
rect 25924 3576 25926 3596
rect 26330 6604 26332 6624
rect 26332 6604 26384 6624
rect 26384 6604 26386 6624
rect 26330 6568 26386 6604
rect 26790 8880 26846 8936
rect 27802 17176 27858 17232
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 27526 10548 27528 10568
rect 27528 10548 27580 10568
rect 27580 10548 27582 10568
rect 27526 10512 27582 10548
rect 27066 8472 27122 8528
rect 26238 6160 26294 6216
rect 26054 4528 26110 4584
rect 26606 7656 26662 7712
rect 26514 4020 26516 4040
rect 26516 4020 26568 4040
rect 26568 4020 26570 4040
rect 26514 3984 26570 4020
rect 27250 7792 27306 7848
rect 27250 5480 27306 5536
rect 27066 4684 27122 4720
rect 27066 4664 27068 4684
rect 27068 4664 27120 4684
rect 27120 4664 27122 4684
rect 26974 3848 27030 3904
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28630 12280 28686 12336
rect 27986 6740 27988 6760
rect 27988 6740 28040 6760
rect 28040 6740 28042 6760
rect 27986 6704 28042 6740
rect 27618 5344 27674 5400
rect 28262 6432 28318 6488
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28538 5752 28594 5808
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 6821 27434 6887 27437
rect 10225 27434 10291 27437
rect 6821 27432 10291 27434
rect 6821 27376 6826 27432
rect 6882 27376 10230 27432
rect 10286 27376 10291 27432
rect 6821 27374 10291 27376
rect 6821 27371 6887 27374
rect 10225 27371 10291 27374
rect 0 27298 800 27328
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 0 27208 800 27238
rect 933 27235 999 27238
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 2589 27026 2655 27029
rect 10041 27026 10107 27029
rect 2589 27024 10107 27026
rect 2589 26968 2594 27024
rect 2650 26968 10046 27024
rect 10102 26968 10107 27024
rect 2589 26966 10107 26968
rect 2589 26963 2655 26966
rect 10041 26963 10107 26966
rect 28441 27026 28507 27029
rect 29200 27026 30000 27056
rect 28441 27024 30000 27026
rect 28441 26968 28446 27024
rect 28502 26968 30000 27024
rect 28441 26966 30000 26968
rect 28441 26963 28507 26966
rect 29200 26936 30000 26966
rect 3785 26890 3851 26893
rect 10041 26890 10107 26893
rect 3785 26888 10107 26890
rect 3785 26832 3790 26888
rect 3846 26832 10046 26888
rect 10102 26832 10107 26888
rect 3785 26830 10107 26832
rect 3785 26827 3851 26830
rect 10041 26827 10107 26830
rect 22737 26890 22803 26893
rect 25681 26890 25747 26893
rect 22737 26888 25747 26890
rect 22737 26832 22742 26888
rect 22798 26832 25686 26888
rect 25742 26832 25747 26888
rect 22737 26830 25747 26832
rect 22737 26827 22803 26830
rect 25681 26827 25747 26830
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 6361 26346 6427 26349
rect 7281 26346 7347 26349
rect 6361 26344 7347 26346
rect 6361 26288 6366 26344
rect 6422 26288 7286 26344
rect 7342 26288 7347 26344
rect 6361 26286 7347 26288
rect 6361 26283 6427 26286
rect 7281 26283 7347 26286
rect 12341 26346 12407 26349
rect 13905 26346 13971 26349
rect 12341 26344 13971 26346
rect 12341 26288 12346 26344
rect 12402 26288 13910 26344
rect 13966 26288 13971 26344
rect 12341 26286 13971 26288
rect 12341 26283 12407 26286
rect 13905 26283 13971 26286
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 9857 26074 9923 26077
rect 14365 26074 14431 26077
rect 9857 26072 14431 26074
rect 9857 26016 9862 26072
rect 9918 26016 14370 26072
rect 14426 26016 14431 26072
rect 9857 26014 14431 26016
rect 9857 26011 9923 26014
rect 14365 26011 14431 26014
rect 3417 25802 3483 25805
rect 8477 25802 8543 25805
rect 3417 25800 8543 25802
rect 3417 25744 3422 25800
rect 3478 25744 8482 25800
rect 8538 25744 8543 25800
rect 3417 25742 8543 25744
rect 3417 25739 3483 25742
rect 8477 25739 8543 25742
rect 20529 25802 20595 25805
rect 25865 25802 25931 25805
rect 20529 25800 25931 25802
rect 20529 25744 20534 25800
rect 20590 25744 25870 25800
rect 25926 25744 25931 25800
rect 20529 25742 25931 25744
rect 20529 25739 20595 25742
rect 25865 25739 25931 25742
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 1945 24986 2011 24989
rect 6361 24986 6427 24989
rect 1945 24984 6427 24986
rect 1945 24928 1950 24984
rect 2006 24928 6366 24984
rect 6422 24928 6427 24984
rect 1945 24926 6427 24928
rect 1945 24923 2011 24926
rect 6361 24923 6427 24926
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 0 23762 800 23792
rect 1577 23762 1643 23765
rect 0 23760 1643 23762
rect 0 23704 1582 23760
rect 1638 23704 1643 23760
rect 0 23702 1643 23704
rect 0 23672 800 23702
rect 1577 23699 1643 23702
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 9673 22946 9739 22949
rect 14549 22946 14615 22949
rect 9673 22944 14615 22946
rect 9673 22888 9678 22944
rect 9734 22888 14554 22944
rect 14610 22888 14615 22944
rect 9673 22886 14615 22888
rect 9673 22883 9739 22886
rect 14549 22883 14615 22886
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 8293 22538 8359 22541
rect 9489 22538 9555 22541
rect 8293 22536 9555 22538
rect 8293 22480 8298 22536
rect 8354 22480 9494 22536
rect 9550 22480 9555 22536
rect 8293 22478 9555 22480
rect 8293 22475 8359 22478
rect 9489 22475 9555 22478
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 8109 22266 8175 22269
rect 8661 22266 8727 22269
rect 8109 22264 8727 22266
rect 8109 22208 8114 22264
rect 8170 22208 8666 22264
rect 8722 22208 8727 22264
rect 8109 22206 8727 22208
rect 8109 22203 8175 22206
rect 8661 22203 8727 22206
rect 19885 22266 19951 22269
rect 21909 22266 21975 22269
rect 19885 22264 21975 22266
rect 19885 22208 19890 22264
rect 19946 22208 21914 22264
rect 21970 22208 21975 22264
rect 19885 22206 21975 22208
rect 19885 22203 19951 22206
rect 21909 22203 21975 22206
rect 5257 22130 5323 22133
rect 8201 22130 8267 22133
rect 8845 22130 8911 22133
rect 5257 22128 8911 22130
rect 5257 22072 5262 22128
rect 5318 22072 8206 22128
rect 8262 22072 8850 22128
rect 8906 22072 8911 22128
rect 5257 22070 8911 22072
rect 5257 22067 5323 22070
rect 8201 22067 8267 22070
rect 8845 22067 8911 22070
rect 9857 22130 9923 22133
rect 18781 22130 18847 22133
rect 9857 22128 18847 22130
rect 9857 22072 9862 22128
rect 9918 22072 18786 22128
rect 18842 22072 18847 22128
rect 9857 22070 18847 22072
rect 9857 22067 9923 22070
rect 18781 22067 18847 22070
rect 27981 22130 28047 22133
rect 29200 22130 30000 22160
rect 27981 22128 30000 22130
rect 27981 22072 27986 22128
rect 28042 22072 30000 22128
rect 27981 22070 30000 22072
rect 27981 22067 28047 22070
rect 29200 22040 30000 22070
rect 5993 21994 6059 21997
rect 10041 21994 10107 21997
rect 10409 21994 10475 21997
rect 5993 21992 10475 21994
rect 5993 21936 5998 21992
rect 6054 21936 10046 21992
rect 10102 21936 10414 21992
rect 10470 21936 10475 21992
rect 5993 21934 10475 21936
rect 5993 21931 6059 21934
rect 10041 21931 10107 21934
rect 10409 21931 10475 21934
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 5533 21450 5599 21453
rect 9121 21450 9187 21453
rect 5533 21448 9187 21450
rect 5533 21392 5538 21448
rect 5594 21392 9126 21448
rect 9182 21392 9187 21448
rect 5533 21390 9187 21392
rect 5533 21387 5599 21390
rect 9121 21387 9187 21390
rect 16481 21450 16547 21453
rect 22737 21450 22803 21453
rect 26601 21450 26667 21453
rect 16481 21448 26667 21450
rect 16481 21392 16486 21448
rect 16542 21392 22742 21448
rect 22798 21392 26606 21448
rect 26662 21392 26667 21448
rect 16481 21390 26667 21392
rect 16481 21387 16547 21390
rect 22737 21387 22803 21390
rect 26601 21387 26667 21390
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 10041 21042 10107 21045
rect 15193 21042 15259 21045
rect 10041 21040 15259 21042
rect 10041 20984 10046 21040
rect 10102 20984 15198 21040
rect 15254 20984 15259 21040
rect 10041 20982 15259 20984
rect 10041 20979 10107 20982
rect 15193 20979 15259 20982
rect 21357 20770 21423 20773
rect 21222 20768 21423 20770
rect 21222 20712 21362 20768
rect 21418 20712 21423 20768
rect 21222 20710 21423 20712
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 15745 20634 15811 20637
rect 21222 20634 21282 20710
rect 21357 20707 21423 20710
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 15745 20632 21282 20634
rect 15745 20576 15750 20632
rect 15806 20576 21282 20632
rect 15745 20574 21282 20576
rect 22277 20634 22343 20637
rect 25129 20634 25195 20637
rect 22277 20632 25195 20634
rect 22277 20576 22282 20632
rect 22338 20576 25134 20632
rect 25190 20576 25195 20632
rect 22277 20574 25195 20576
rect 15745 20571 15811 20574
rect 22277 20571 22343 20574
rect 25129 20571 25195 20574
rect 2957 20362 3023 20365
rect 2730 20360 3023 20362
rect 2730 20304 2962 20360
rect 3018 20304 3023 20360
rect 2730 20302 3023 20304
rect 0 20226 800 20256
rect 2730 20226 2790 20302
rect 2957 20299 3023 20302
rect 9765 20362 9831 20365
rect 10593 20362 10659 20365
rect 9765 20360 10659 20362
rect 9765 20304 9770 20360
rect 9826 20304 10598 20360
rect 10654 20304 10659 20360
rect 9765 20302 10659 20304
rect 9765 20299 9831 20302
rect 10593 20299 10659 20302
rect 0 20166 2790 20226
rect 0 20136 800 20166
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 7281 19954 7347 19957
rect 10409 19954 10475 19957
rect 7281 19952 10475 19954
rect 7281 19896 7286 19952
rect 7342 19896 10414 19952
rect 10470 19896 10475 19952
rect 7281 19894 10475 19896
rect 7281 19891 7347 19894
rect 10409 19891 10475 19894
rect 8385 19818 8451 19821
rect 11329 19818 11395 19821
rect 8385 19816 11395 19818
rect 8385 19760 8390 19816
rect 8446 19760 11334 19816
rect 11390 19760 11395 19816
rect 8385 19758 11395 19760
rect 8385 19755 8451 19758
rect 11329 19755 11395 19758
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 20989 19410 21055 19413
rect 21449 19410 21515 19413
rect 20989 19408 21515 19410
rect 20989 19352 20994 19408
rect 21050 19352 21454 19408
rect 21510 19352 21515 19408
rect 20989 19350 21515 19352
rect 20989 19347 21055 19350
rect 21449 19347 21515 19350
rect 21081 19274 21147 19277
rect 24485 19274 24551 19277
rect 21081 19272 24551 19274
rect 21081 19216 21086 19272
rect 21142 19216 24490 19272
rect 24546 19216 24551 19272
rect 21081 19214 24551 19216
rect 21081 19211 21147 19214
rect 24485 19211 24551 19214
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 5441 18052 5507 18053
rect 5390 18050 5396 18052
rect 5350 17990 5396 18050
rect 5460 18048 5507 18052
rect 5502 17992 5507 18048
rect 5390 17988 5396 17990
rect 5460 17988 5507 17992
rect 5441 17987 5507 17988
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 6361 17914 6427 17917
rect 11053 17914 11119 17917
rect 6361 17912 11119 17914
rect 6361 17856 6366 17912
rect 6422 17856 11058 17912
rect 11114 17856 11119 17912
rect 6361 17854 11119 17856
rect 6361 17851 6427 17854
rect 11053 17851 11119 17854
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 5441 17234 5507 17237
rect 20437 17234 20503 17237
rect 5441 17232 20503 17234
rect 5441 17176 5446 17232
rect 5502 17176 20442 17232
rect 20498 17176 20503 17232
rect 5441 17174 20503 17176
rect 5441 17171 5507 17174
rect 20437 17171 20503 17174
rect 27797 17234 27863 17237
rect 29200 17234 30000 17264
rect 27797 17232 30000 17234
rect 27797 17176 27802 17232
rect 27858 17176 30000 17232
rect 27797 17174 30000 17176
rect 27797 17171 27863 17174
rect 29200 17144 30000 17174
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 20621 16690 20687 16693
rect 23197 16690 23263 16693
rect 20621 16688 23263 16690
rect 20621 16632 20626 16688
rect 20682 16632 23202 16688
rect 23258 16632 23263 16688
rect 20621 16630 23263 16632
rect 20621 16627 20687 16630
rect 23197 16627 23263 16630
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 20529 16146 20595 16149
rect 20989 16146 21055 16149
rect 20529 16144 21055 16146
rect 20529 16088 20534 16144
rect 20590 16088 20994 16144
rect 21050 16088 21055 16144
rect 20529 16086 21055 16088
rect 20529 16083 20595 16086
rect 20989 16083 21055 16086
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 17125 15466 17191 15469
rect 19149 15466 19215 15469
rect 17125 15464 19215 15466
rect 17125 15408 17130 15464
rect 17186 15408 19154 15464
rect 19210 15408 19215 15464
rect 17125 15406 19215 15408
rect 17125 15403 17191 15406
rect 19149 15403 19215 15406
rect 4521 15330 4587 15333
rect 4838 15330 4844 15332
rect 4521 15328 4844 15330
rect 4521 15272 4526 15328
rect 4582 15272 4844 15328
rect 4521 15270 4844 15272
rect 4521 15267 4587 15270
rect 4838 15268 4844 15270
rect 4908 15268 4914 15332
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 10225 14378 10291 14381
rect 14549 14378 14615 14381
rect 10225 14376 14615 14378
rect 10225 14320 10230 14376
rect 10286 14320 14554 14376
rect 14610 14320 14615 14376
rect 10225 14318 14615 14320
rect 10225 14315 10291 14318
rect 14549 14315 14615 14318
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 8017 13970 8083 13973
rect 8477 13970 8543 13973
rect 8017 13968 8543 13970
rect 8017 13912 8022 13968
rect 8078 13912 8482 13968
rect 8538 13912 8543 13968
rect 8017 13910 8543 13912
rect 8017 13907 8083 13910
rect 8477 13907 8543 13910
rect 25221 13970 25287 13973
rect 27061 13970 27127 13973
rect 25221 13968 27127 13970
rect 25221 13912 25226 13968
rect 25282 13912 27066 13968
rect 27122 13912 27127 13968
rect 25221 13910 27127 13912
rect 25221 13907 25287 13910
rect 27061 13907 27127 13910
rect 24577 13834 24643 13837
rect 26141 13834 26207 13837
rect 24577 13832 26207 13834
rect 24577 13776 24582 13832
rect 24638 13776 26146 13832
rect 26202 13776 26207 13832
rect 24577 13774 26207 13776
rect 24577 13771 24643 13774
rect 26141 13771 26207 13774
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 0 13154 800 13184
rect 933 13154 999 13157
rect 0 13152 999 13154
rect 0 13096 938 13152
rect 994 13096 999 13152
rect 0 13094 999 13096
rect 0 13064 800 13094
rect 933 13091 999 13094
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 5073 12746 5139 12749
rect 9857 12746 9923 12749
rect 5073 12744 9923 12746
rect 5073 12688 5078 12744
rect 5134 12688 9862 12744
rect 9918 12688 9923 12744
rect 5073 12686 9923 12688
rect 5073 12683 5139 12686
rect 9857 12683 9923 12686
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 9581 12474 9647 12477
rect 11237 12474 11303 12477
rect 9581 12472 11303 12474
rect 9581 12416 9586 12472
rect 9642 12416 11242 12472
rect 11298 12416 11303 12472
rect 9581 12414 11303 12416
rect 9581 12411 9647 12414
rect 11237 12411 11303 12414
rect 19793 12338 19859 12341
rect 22870 12338 22876 12340
rect 19793 12336 22876 12338
rect 19793 12280 19798 12336
rect 19854 12280 22876 12336
rect 19793 12278 22876 12280
rect 19793 12275 19859 12278
rect 22870 12276 22876 12278
rect 22940 12276 22946 12340
rect 28625 12338 28691 12341
rect 29200 12338 30000 12368
rect 28625 12336 30000 12338
rect 28625 12280 28630 12336
rect 28686 12280 30000 12336
rect 28625 12278 30000 12280
rect 28625 12275 28691 12278
rect 29200 12248 30000 12278
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 4613 11930 4679 11933
rect 4838 11930 4844 11932
rect 4613 11928 4844 11930
rect 4613 11872 4618 11928
rect 4674 11872 4844 11928
rect 4613 11870 4844 11872
rect 4613 11867 4679 11870
rect 4838 11868 4844 11870
rect 4908 11868 4914 11932
rect 24025 11930 24091 11933
rect 26601 11930 26667 11933
rect 23982 11928 26667 11930
rect 23982 11872 24030 11928
rect 24086 11872 26606 11928
rect 26662 11872 26667 11928
rect 23982 11870 26667 11872
rect 23982 11867 24091 11870
rect 26601 11867 26667 11870
rect 5349 11796 5415 11797
rect 5349 11794 5396 11796
rect 5268 11792 5396 11794
rect 5460 11794 5466 11796
rect 17769 11794 17835 11797
rect 5460 11792 17835 11794
rect 5268 11736 5354 11792
rect 5460 11736 17774 11792
rect 17830 11736 17835 11792
rect 5268 11734 5396 11736
rect 5349 11732 5396 11734
rect 5460 11734 17835 11736
rect 5460 11732 5466 11734
rect 5349 11731 5415 11732
rect 17769 11731 17835 11734
rect 6821 11658 6887 11661
rect 11053 11658 11119 11661
rect 6821 11656 11119 11658
rect 6821 11600 6826 11656
rect 6882 11600 11058 11656
rect 11114 11600 11119 11656
rect 6821 11598 11119 11600
rect 6821 11595 6887 11598
rect 11053 11595 11119 11598
rect 17493 11658 17559 11661
rect 23982 11658 24042 11867
rect 17493 11656 24042 11658
rect 17493 11600 17498 11656
rect 17554 11600 24042 11656
rect 17493 11598 24042 11600
rect 17493 11595 17559 11598
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 24485 11386 24551 11389
rect 24710 11386 24716 11388
rect 24485 11384 24716 11386
rect 24485 11328 24490 11384
rect 24546 11328 24716 11384
rect 24485 11326 24716 11328
rect 24485 11323 24551 11326
rect 24710 11324 24716 11326
rect 24780 11324 24786 11388
rect 2957 11250 3023 11253
rect 8385 11250 8451 11253
rect 2957 11248 8451 11250
rect 2957 11192 2962 11248
rect 3018 11192 8390 11248
rect 8446 11192 8451 11248
rect 2957 11190 8451 11192
rect 2957 11187 3023 11190
rect 8385 11187 8451 11190
rect 19425 11250 19491 11253
rect 25221 11250 25287 11253
rect 19425 11248 25287 11250
rect 19425 11192 19430 11248
rect 19486 11192 25226 11248
rect 25282 11192 25287 11248
rect 19425 11190 25287 11192
rect 19425 11187 19491 11190
rect 25221 11187 25287 11190
rect 2681 11114 2747 11117
rect 8477 11114 8543 11117
rect 2681 11112 8543 11114
rect 2681 11056 2686 11112
rect 2742 11056 8482 11112
rect 8538 11056 8543 11112
rect 2681 11054 8543 11056
rect 2681 11051 2747 11054
rect 8477 11051 8543 11054
rect 25957 11116 26023 11117
rect 25957 11112 26004 11116
rect 26068 11114 26074 11116
rect 25957 11056 25962 11112
rect 25957 11052 26004 11056
rect 26068 11054 26114 11114
rect 26068 11052 26074 11054
rect 25957 11051 26023 11052
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 4838 10644 4844 10708
rect 4908 10706 4914 10708
rect 11513 10706 11579 10709
rect 4908 10704 11579 10706
rect 4908 10648 11518 10704
rect 11574 10648 11579 10704
rect 4908 10646 11579 10648
rect 4908 10644 4914 10646
rect 11513 10643 11579 10646
rect 22185 10570 22251 10573
rect 27521 10570 27587 10573
rect 22185 10568 27587 10570
rect 22185 10512 22190 10568
rect 22246 10512 27526 10568
rect 27582 10512 27587 10568
rect 22185 10510 27587 10512
rect 22185 10507 22251 10510
rect 27521 10507 27587 10510
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 21357 10162 21423 10165
rect 21725 10162 21791 10165
rect 21357 10160 21791 10162
rect 21357 10104 21362 10160
rect 21418 10104 21730 10160
rect 21786 10104 21791 10160
rect 21357 10102 21791 10104
rect 21357 10099 21423 10102
rect 21725 10099 21791 10102
rect 24117 10162 24183 10165
rect 26233 10162 26299 10165
rect 24117 10160 26299 10162
rect 24117 10104 24122 10160
rect 24178 10104 26238 10160
rect 26294 10104 26299 10160
rect 24117 10102 26299 10104
rect 24117 10099 24183 10102
rect 26233 10099 26299 10102
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 20345 9618 20411 9621
rect 20897 9618 20963 9621
rect 20345 9616 20963 9618
rect 20345 9560 20350 9616
rect 20406 9560 20902 9616
rect 20958 9560 20963 9616
rect 20345 9558 20963 9560
rect 20345 9555 20411 9558
rect 20897 9555 20963 9558
rect 21265 9618 21331 9621
rect 21817 9618 21883 9621
rect 26601 9618 26667 9621
rect 21265 9616 26667 9618
rect 21265 9560 21270 9616
rect 21326 9560 21822 9616
rect 21878 9560 26606 9616
rect 26662 9560 26667 9616
rect 21265 9558 26667 9560
rect 21265 9555 21331 9558
rect 21817 9555 21883 9558
rect 26601 9555 26667 9558
rect 20069 9482 20135 9485
rect 26233 9482 26299 9485
rect 20069 9480 26299 9482
rect 20069 9424 20074 9480
rect 20130 9424 26238 9480
rect 26294 9424 26299 9480
rect 20069 9422 26299 9424
rect 20069 9419 20135 9422
rect 26233 9419 26299 9422
rect 19425 9346 19491 9349
rect 23289 9346 23355 9349
rect 19425 9344 23355 9346
rect 19425 9288 19430 9344
rect 19486 9288 23294 9344
rect 23350 9288 23355 9344
rect 19425 9286 23355 9288
rect 19425 9283 19491 9286
rect 23289 9283 23355 9286
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 19609 9210 19675 9213
rect 21725 9210 21791 9213
rect 19609 9208 21791 9210
rect 19609 9152 19614 9208
rect 19670 9152 21730 9208
rect 21786 9152 21791 9208
rect 19609 9150 21791 9152
rect 19609 9147 19675 9150
rect 21725 9147 21791 9150
rect 22277 9210 22343 9213
rect 24025 9210 24091 9213
rect 22277 9208 24091 9210
rect 22277 9152 22282 9208
rect 22338 9152 24030 9208
rect 24086 9152 24091 9208
rect 22277 9150 24091 9152
rect 22277 9147 22343 9150
rect 24025 9147 24091 9150
rect 20069 9074 20135 9077
rect 23841 9074 23907 9077
rect 24485 9074 24551 9077
rect 20069 9072 24551 9074
rect 20069 9016 20074 9072
rect 20130 9016 23846 9072
rect 23902 9016 24490 9072
rect 24546 9016 24551 9072
rect 20069 9014 24551 9016
rect 20069 9011 20135 9014
rect 23841 9011 23907 9014
rect 24485 9011 24551 9014
rect 24761 9074 24827 9077
rect 25814 9074 25820 9076
rect 24761 9072 25820 9074
rect 24761 9016 24766 9072
rect 24822 9016 25820 9072
rect 24761 9014 25820 9016
rect 24761 9011 24827 9014
rect 25814 9012 25820 9014
rect 25884 9012 25890 9076
rect 16205 8938 16271 8941
rect 26785 8938 26851 8941
rect 16205 8936 26851 8938
rect 16205 8880 16210 8936
rect 16266 8880 26790 8936
rect 26846 8880 26851 8936
rect 16205 8878 26851 8880
rect 16205 8875 16271 8878
rect 26785 8875 26851 8878
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 20437 8666 20503 8669
rect 20662 8666 20668 8668
rect 20437 8664 20668 8666
rect 20437 8608 20442 8664
rect 20498 8608 20668 8664
rect 20437 8606 20668 8608
rect 20437 8603 20503 8606
rect 20662 8604 20668 8606
rect 20732 8604 20738 8668
rect 21081 8530 21147 8533
rect 27061 8530 27127 8533
rect 21081 8528 27127 8530
rect 21081 8472 21086 8528
rect 21142 8472 27066 8528
rect 27122 8472 27127 8528
rect 21081 8470 27127 8472
rect 21081 8467 21147 8470
rect 27061 8467 27127 8470
rect 17585 8394 17651 8397
rect 21265 8394 21331 8397
rect 23841 8394 23907 8397
rect 24761 8394 24827 8397
rect 17585 8392 19810 8394
rect 17585 8336 17590 8392
rect 17646 8336 19810 8392
rect 17585 8334 19810 8336
rect 17585 8331 17651 8334
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 9581 7986 9647 7989
rect 11881 7986 11947 7989
rect 9581 7984 11947 7986
rect 9581 7928 9586 7984
rect 9642 7928 11886 7984
rect 11942 7928 11947 7984
rect 9581 7926 11947 7928
rect 9581 7923 9647 7926
rect 11881 7923 11947 7926
rect 15101 7850 15167 7853
rect 19750 7850 19810 8334
rect 21265 8392 22110 8394
rect 21265 8336 21270 8392
rect 21326 8336 22110 8392
rect 21265 8334 22110 8336
rect 21265 8331 21331 8334
rect 20069 8122 20135 8125
rect 21449 8122 21515 8125
rect 20069 8120 21515 8122
rect 20069 8064 20074 8120
rect 20130 8064 21454 8120
rect 21510 8064 21515 8120
rect 20069 8062 21515 8064
rect 20069 8059 20135 8062
rect 21449 8059 21515 8062
rect 22050 7986 22110 8334
rect 23841 8392 24827 8394
rect 23841 8336 23846 8392
rect 23902 8336 24766 8392
rect 24822 8336 24827 8392
rect 23841 8334 24827 8336
rect 23841 8331 23907 8334
rect 24761 8331 24827 8334
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 24393 8122 24459 8125
rect 25129 8122 25195 8125
rect 24393 8120 25195 8122
rect 24393 8064 24398 8120
rect 24454 8064 25134 8120
rect 25190 8064 25195 8120
rect 24393 8062 25195 8064
rect 24393 8059 24459 8062
rect 25129 8059 25195 8062
rect 26417 7986 26483 7989
rect 22050 7984 26483 7986
rect 22050 7928 26422 7984
rect 26478 7928 26483 7984
rect 22050 7926 26483 7928
rect 26417 7923 26483 7926
rect 27245 7850 27311 7853
rect 15101 7848 17234 7850
rect 15101 7792 15106 7848
rect 15162 7792 17234 7848
rect 15101 7790 17234 7792
rect 19750 7848 27311 7850
rect 19750 7792 27250 7848
rect 27306 7792 27311 7848
rect 19750 7790 27311 7792
rect 15101 7787 15167 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 5625 7578 5691 7581
rect 6361 7578 6427 7581
rect 5625 7576 6427 7578
rect 5625 7520 5630 7576
rect 5686 7520 6366 7576
rect 6422 7520 6427 7576
rect 5625 7518 6427 7520
rect 5625 7515 5691 7518
rect 6361 7515 6427 7518
rect 17174 7306 17234 7790
rect 27245 7787 27311 7790
rect 23381 7714 23447 7717
rect 26601 7714 26667 7717
rect 23381 7712 26667 7714
rect 23381 7656 23386 7712
rect 23442 7656 26606 7712
rect 26662 7656 26667 7712
rect 23381 7654 26667 7656
rect 23381 7651 23447 7654
rect 26601 7651 26667 7654
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 22553 7578 22619 7581
rect 22553 7576 24778 7578
rect 22553 7520 22558 7576
rect 22614 7520 24778 7576
rect 22553 7518 24778 7520
rect 22553 7515 22619 7518
rect 17401 7442 17467 7445
rect 23841 7442 23907 7445
rect 17401 7440 23907 7442
rect 17401 7384 17406 7440
rect 17462 7384 23846 7440
rect 23902 7384 23907 7440
rect 17401 7382 23907 7384
rect 17401 7379 17467 7382
rect 23841 7379 23907 7382
rect 24301 7442 24367 7445
rect 24577 7442 24643 7445
rect 24301 7440 24643 7442
rect 24301 7384 24306 7440
rect 24362 7384 24582 7440
rect 24638 7384 24643 7440
rect 24301 7382 24643 7384
rect 24718 7442 24778 7518
rect 29200 7442 30000 7472
rect 24718 7382 30000 7442
rect 24301 7379 24367 7382
rect 24577 7379 24643 7382
rect 29200 7352 30000 7382
rect 24301 7306 24367 7309
rect 17174 7304 24367 7306
rect 17174 7248 24306 7304
rect 24362 7248 24367 7304
rect 17174 7246 24367 7248
rect 24301 7243 24367 7246
rect 19609 7170 19675 7173
rect 24894 7170 24900 7172
rect 19609 7168 24900 7170
rect 19609 7112 19614 7168
rect 19670 7112 24900 7168
rect 19609 7110 24900 7112
rect 19609 7107 19675 7110
rect 24894 7108 24900 7110
rect 24964 7108 24970 7172
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 16665 7034 16731 7037
rect 17902 7034 17908 7036
rect 16665 7032 17908 7034
rect 16665 6976 16670 7032
rect 16726 6976 17908 7032
rect 16665 6974 17908 6976
rect 16665 6971 16731 6974
rect 17902 6972 17908 6974
rect 17972 6972 17978 7036
rect 18965 7034 19031 7037
rect 22001 7034 22067 7037
rect 18965 7032 22067 7034
rect 18965 6976 18970 7032
rect 19026 6976 22006 7032
rect 22062 6976 22067 7032
rect 18965 6974 22067 6976
rect 18965 6971 19031 6974
rect 22001 6971 22067 6974
rect 23422 6972 23428 7036
rect 23492 7034 23498 7036
rect 24117 7034 24183 7037
rect 23492 7032 24183 7034
rect 23492 6976 24122 7032
rect 24178 6976 24183 7032
rect 23492 6974 24183 6976
rect 23492 6972 23498 6974
rect 24117 6971 24183 6974
rect 5165 6898 5231 6901
rect 14641 6898 14707 6901
rect 5165 6896 14707 6898
rect 5165 6840 5170 6896
rect 5226 6840 14646 6896
rect 14702 6840 14707 6896
rect 5165 6838 14707 6840
rect 5165 6835 5231 6838
rect 14641 6835 14707 6838
rect 17585 6898 17651 6901
rect 23933 6898 23999 6901
rect 17585 6896 23999 6898
rect 17585 6840 17590 6896
rect 17646 6840 23938 6896
rect 23994 6840 23999 6896
rect 17585 6838 23999 6840
rect 17585 6835 17651 6838
rect 23933 6835 23999 6838
rect 16573 6762 16639 6765
rect 27981 6762 28047 6765
rect 16573 6760 28047 6762
rect 16573 6704 16578 6760
rect 16634 6704 27986 6760
rect 28042 6704 28047 6760
rect 16573 6702 28047 6704
rect 16573 6699 16639 6702
rect 27981 6699 28047 6702
rect 16665 6626 16731 6629
rect 18505 6626 18571 6629
rect 21265 6626 21331 6629
rect 16665 6624 21331 6626
rect 16665 6568 16670 6624
rect 16726 6568 18510 6624
rect 18566 6568 21270 6624
rect 21326 6568 21331 6624
rect 16665 6566 21331 6568
rect 16665 6563 16731 6566
rect 18505 6563 18571 6566
rect 21265 6563 21331 6566
rect 23381 6626 23447 6629
rect 25037 6626 25103 6629
rect 23381 6624 25103 6626
rect 23381 6568 23386 6624
rect 23442 6568 25042 6624
rect 25098 6568 25103 6624
rect 23381 6566 25103 6568
rect 23381 6563 23447 6566
rect 25037 6563 25103 6566
rect 25681 6626 25747 6629
rect 26325 6626 26391 6629
rect 25681 6624 26391 6626
rect 25681 6568 25686 6624
rect 25742 6568 26330 6624
rect 26386 6568 26391 6624
rect 25681 6566 26391 6568
rect 25681 6563 25747 6566
rect 26325 6563 26391 6566
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 19057 6490 19123 6493
rect 19609 6490 19675 6493
rect 19057 6488 19675 6490
rect 19057 6432 19062 6488
rect 19118 6432 19614 6488
rect 19670 6432 19675 6488
rect 19057 6430 19675 6432
rect 19057 6427 19123 6430
rect 19609 6427 19675 6430
rect 23933 6488 23999 6493
rect 23933 6432 23938 6488
rect 23994 6432 23999 6488
rect 23933 6427 23999 6432
rect 24485 6490 24551 6493
rect 28257 6490 28323 6493
rect 24485 6488 28323 6490
rect 24485 6432 24490 6488
rect 24546 6432 28262 6488
rect 28318 6432 28323 6488
rect 24485 6430 28323 6432
rect 24485 6427 24551 6430
rect 28257 6427 28323 6430
rect 14733 6218 14799 6221
rect 22829 6220 22895 6221
rect 22829 6218 22876 6220
rect 2730 6216 14799 6218
rect 2730 6160 14738 6216
rect 14794 6160 14799 6216
rect 2730 6158 14799 6160
rect 22784 6216 22876 6218
rect 22784 6160 22834 6216
rect 22784 6158 22876 6160
rect 0 6082 800 6112
rect 2730 6082 2790 6158
rect 14733 6155 14799 6158
rect 22829 6156 22876 6158
rect 22940 6156 22946 6220
rect 23936 6218 23996 6427
rect 26233 6218 26299 6221
rect 23936 6216 26299 6218
rect 23936 6160 26238 6216
rect 26294 6160 26299 6216
rect 23936 6158 26299 6160
rect 22829 6155 22895 6156
rect 26233 6155 26299 6158
rect 0 6022 2790 6082
rect 0 5992 800 6022
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 20713 5946 20779 5949
rect 20713 5944 25192 5946
rect 20713 5888 20718 5944
rect 20774 5888 25192 5944
rect 20713 5886 25192 5888
rect 20713 5883 20779 5886
rect 10041 5810 10107 5813
rect 14365 5810 14431 5813
rect 10041 5808 14431 5810
rect 10041 5752 10046 5808
rect 10102 5752 14370 5808
rect 14426 5752 14431 5808
rect 10041 5750 14431 5752
rect 10041 5747 10107 5750
rect 14365 5747 14431 5750
rect 18321 5810 18387 5813
rect 21541 5810 21607 5813
rect 18321 5808 21607 5810
rect 18321 5752 18326 5808
rect 18382 5752 21546 5808
rect 21602 5752 21607 5808
rect 18321 5750 21607 5752
rect 25132 5810 25192 5886
rect 28533 5810 28599 5813
rect 25132 5808 28599 5810
rect 25132 5752 28538 5808
rect 28594 5752 28599 5808
rect 25132 5750 28599 5752
rect 18321 5747 18387 5750
rect 21541 5747 21607 5750
rect 28533 5747 28599 5750
rect 15837 5538 15903 5541
rect 21449 5538 21515 5541
rect 15837 5536 21515 5538
rect 15837 5480 15842 5536
rect 15898 5480 21454 5536
rect 21510 5480 21515 5536
rect 15837 5478 21515 5480
rect 15837 5475 15903 5478
rect 21449 5475 21515 5478
rect 24710 5476 24716 5540
rect 24780 5476 24786 5540
rect 24894 5476 24900 5540
rect 24964 5538 24970 5540
rect 27245 5538 27311 5541
rect 24964 5536 27311 5538
rect 24964 5480 27250 5536
rect 27306 5480 27311 5536
rect 24964 5478 27311 5480
rect 24964 5476 24970 5478
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 24718 5402 24778 5476
rect 27245 5475 27311 5478
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 27613 5402 27679 5405
rect 24718 5400 27679 5402
rect 24718 5344 27618 5400
rect 27674 5344 27679 5400
rect 24718 5342 27679 5344
rect 27613 5339 27679 5342
rect 14089 5266 14155 5269
rect 24393 5266 24459 5269
rect 14089 5264 24459 5266
rect 14089 5208 14094 5264
rect 14150 5208 24398 5264
rect 24454 5208 24459 5264
rect 14089 5206 24459 5208
rect 14089 5203 14155 5206
rect 24393 5203 24459 5206
rect 10133 5130 10199 5133
rect 14273 5130 14339 5133
rect 10133 5128 14339 5130
rect 10133 5072 10138 5128
rect 10194 5072 14278 5128
rect 14334 5072 14339 5128
rect 10133 5070 14339 5072
rect 10133 5067 10199 5070
rect 14273 5067 14339 5070
rect 17769 5130 17835 5133
rect 18781 5130 18847 5133
rect 17769 5128 18847 5130
rect 17769 5072 17774 5128
rect 17830 5072 18786 5128
rect 18842 5072 18847 5128
rect 17769 5070 18847 5072
rect 17769 5067 17835 5070
rect 18781 5067 18847 5070
rect 18965 5130 19031 5133
rect 25313 5130 25379 5133
rect 18965 5128 25379 5130
rect 18965 5072 18970 5128
rect 19026 5072 25318 5128
rect 25374 5072 25379 5128
rect 18965 5070 25379 5072
rect 18965 5067 19031 5070
rect 25313 5067 25379 5070
rect 19333 4994 19399 4997
rect 22185 4994 22251 4997
rect 19333 4992 22251 4994
rect 19333 4936 19338 4992
rect 19394 4936 22190 4992
rect 22246 4936 22251 4992
rect 19333 4934 22251 4936
rect 19333 4931 19399 4934
rect 22185 4931 22251 4934
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 20069 4858 20135 4861
rect 21909 4858 21975 4861
rect 20069 4856 21975 4858
rect 20069 4800 20074 4856
rect 20130 4800 21914 4856
rect 21970 4800 21975 4856
rect 20069 4798 21975 4800
rect 20069 4795 20135 4798
rect 21909 4795 21975 4798
rect 20662 4660 20668 4724
rect 20732 4722 20738 4724
rect 27061 4722 27127 4725
rect 20732 4720 27127 4722
rect 20732 4664 27066 4720
rect 27122 4664 27127 4720
rect 20732 4662 27127 4664
rect 20732 4660 20738 4662
rect 27061 4659 27127 4662
rect 17401 4586 17467 4589
rect 26049 4586 26115 4589
rect 17401 4584 26115 4586
rect 17401 4528 17406 4584
rect 17462 4528 26054 4584
rect 26110 4528 26115 4584
rect 17401 4526 26115 4528
rect 17401 4523 17467 4526
rect 26049 4523 26115 4526
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 5349 4178 5415 4181
rect 23381 4178 23447 4181
rect 5349 4176 23447 4178
rect 5349 4120 5354 4176
rect 5410 4120 23386 4176
rect 23442 4120 23447 4176
rect 5349 4118 23447 4120
rect 5349 4115 5415 4118
rect 23381 4115 23447 4118
rect 6269 4042 6335 4045
rect 8109 4042 8175 4045
rect 15653 4042 15719 4045
rect 6269 4040 15719 4042
rect 6269 3984 6274 4040
rect 6330 3984 8114 4040
rect 8170 3984 15658 4040
rect 15714 3984 15719 4040
rect 6269 3982 15719 3984
rect 6269 3979 6335 3982
rect 8109 3979 8175 3982
rect 15653 3979 15719 3982
rect 16297 4042 16363 4045
rect 26509 4042 26575 4045
rect 16297 4040 26575 4042
rect 16297 3984 16302 4040
rect 16358 3984 26514 4040
rect 26570 3984 26575 4040
rect 16297 3982 26575 3984
rect 16297 3979 16363 3982
rect 26509 3979 26575 3982
rect 18689 3906 18755 3909
rect 22921 3906 22987 3909
rect 25773 3908 25839 3909
rect 25773 3906 25820 3908
rect 18689 3904 22987 3906
rect 18689 3848 18694 3904
rect 18750 3848 22926 3904
rect 22982 3848 22987 3904
rect 18689 3846 22987 3848
rect 25728 3904 25820 3906
rect 25728 3848 25778 3904
rect 25728 3846 25820 3848
rect 18689 3843 18755 3846
rect 22921 3843 22987 3846
rect 25773 3844 25820 3846
rect 25884 3844 25890 3908
rect 25998 3844 26004 3908
rect 26068 3906 26074 3908
rect 26969 3906 27035 3909
rect 26068 3904 27035 3906
rect 26068 3848 26974 3904
rect 27030 3848 27035 3904
rect 26068 3846 27035 3848
rect 26068 3844 26074 3846
rect 25773 3843 25839 3844
rect 26969 3843 27035 3846
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 6545 3770 6611 3773
rect 9121 3770 9187 3773
rect 6545 3768 9187 3770
rect 6545 3712 6550 3768
rect 6606 3712 9126 3768
rect 9182 3712 9187 3768
rect 6545 3710 9187 3712
rect 6545 3707 6611 3710
rect 9121 3707 9187 3710
rect 16757 3634 16823 3637
rect 20989 3634 21055 3637
rect 25865 3634 25931 3637
rect 16757 3632 21055 3634
rect 16757 3576 16762 3632
rect 16818 3576 20994 3632
rect 21050 3576 21055 3632
rect 16757 3574 21055 3576
rect 16757 3571 16823 3574
rect 20989 3571 21055 3574
rect 21222 3632 25931 3634
rect 21222 3576 25870 3632
rect 25926 3576 25931 3632
rect 21222 3574 25931 3576
rect 1853 3498 1919 3501
rect 5165 3498 5231 3501
rect 6729 3498 6795 3501
rect 1853 3496 6795 3498
rect 1853 3440 1858 3496
rect 1914 3440 5170 3496
rect 5226 3440 6734 3496
rect 6790 3440 6795 3496
rect 1853 3438 6795 3440
rect 1853 3435 1919 3438
rect 5165 3435 5231 3438
rect 6729 3435 6795 3438
rect 12341 3498 12407 3501
rect 17309 3498 17375 3501
rect 12341 3496 17375 3498
rect 12341 3440 12346 3496
rect 12402 3440 17314 3496
rect 17370 3440 17375 3496
rect 12341 3438 17375 3440
rect 12341 3435 12407 3438
rect 17309 3435 17375 3438
rect 2497 3362 2563 3365
rect 3785 3362 3851 3365
rect 2497 3360 3851 3362
rect 2497 3304 2502 3360
rect 2558 3304 3790 3360
rect 3846 3304 3851 3360
rect 2497 3302 3851 3304
rect 2497 3299 2563 3302
rect 3785 3299 3851 3302
rect 15929 3362 15995 3365
rect 16389 3362 16455 3365
rect 21222 3362 21282 3574
rect 25865 3571 25931 3574
rect 24853 3498 24919 3501
rect 15929 3360 16314 3362
rect 15929 3304 15934 3360
rect 15990 3304 16314 3360
rect 15929 3302 16314 3304
rect 15929 3299 15995 3302
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 16254 3226 16314 3302
rect 16389 3360 21282 3362
rect 16389 3304 16394 3360
rect 16450 3304 21282 3360
rect 16389 3302 21282 3304
rect 21406 3496 24919 3498
rect 21406 3440 24858 3496
rect 24914 3440 24919 3496
rect 21406 3438 24919 3440
rect 16389 3299 16455 3302
rect 21406 3226 21466 3438
rect 24853 3435 24919 3438
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 16254 3166 21466 3226
rect 15745 3090 15811 3093
rect 24025 3090 24091 3093
rect 15745 3088 24091 3090
rect 15745 3032 15750 3088
rect 15806 3032 24030 3088
rect 24086 3032 24091 3088
rect 15745 3030 24091 3032
rect 15745 3027 15811 3030
rect 24025 3027 24091 3030
rect 4337 2954 4403 2957
rect 24393 2954 24459 2957
rect 4337 2952 24459 2954
rect 4337 2896 4342 2952
rect 4398 2896 24398 2952
rect 24454 2896 24459 2952
rect 4337 2894 24459 2896
rect 4337 2891 4403 2894
rect 24393 2891 24459 2894
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 21909 2682 21975 2685
rect 23841 2682 23907 2685
rect 21909 2680 23907 2682
rect 21909 2624 21914 2680
rect 21970 2624 23846 2680
rect 23902 2624 23907 2680
rect 21909 2622 23907 2624
rect 21909 2619 21975 2622
rect 23841 2619 23907 2622
rect 6269 2546 6335 2549
rect 22553 2546 22619 2549
rect 29200 2546 30000 2576
rect 6269 2544 22619 2546
rect 6269 2488 6274 2544
rect 6330 2488 22558 2544
rect 22614 2488 22619 2544
rect 6269 2486 22619 2488
rect 6269 2483 6335 2486
rect 22553 2483 22619 2486
rect 25638 2486 30000 2546
rect 5993 2410 6059 2413
rect 23422 2410 23428 2412
rect 5993 2408 23428 2410
rect 5993 2352 5998 2408
rect 6054 2352 23428 2408
rect 5993 2350 23428 2352
rect 5993 2347 6059 2350
rect 23422 2348 23428 2350
rect 23492 2348 23498 2412
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 17902 1940 17908 2004
rect 17972 2002 17978 2004
rect 25638 2002 25698 2486
rect 29200 2456 30000 2486
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 17972 1942 25698 2002
rect 17972 1940 17978 1942
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 5396 18048 5460 18052
rect 5396 17992 5446 18048
rect 5446 17992 5460 18048
rect 5396 17988 5460 17992
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 4844 15268 4908 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 22876 12276 22940 12340
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4844 11868 4908 11932
rect 5396 11792 5460 11796
rect 5396 11736 5410 11792
rect 5410 11736 5460 11792
rect 5396 11732 5460 11736
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 24716 11324 24780 11388
rect 26004 11112 26068 11116
rect 26004 11056 26018 11112
rect 26018 11056 26068 11112
rect 26004 11052 26068 11056
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4844 10644 4908 10708
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 25820 9012 25884 9076
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 20668 8604 20732 8668
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 24900 7108 24964 7172
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 17908 6972 17972 7036
rect 23428 6972 23492 7036
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 22876 6216 22940 6220
rect 22876 6160 22890 6216
rect 22890 6160 22940 6216
rect 22876 6156 22940 6160
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 24716 5476 24780 5540
rect 24900 5476 24964 5540
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 20668 4660 20732 4724
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 25820 3904 25884 3908
rect 25820 3848 25834 3904
rect 25834 3848 25884 3904
rect 25820 3844 25884 3848
rect 26004 3844 26068 3908
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 23428 2348 23492 2412
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 17908 1940 17972 2004
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 7890 27232 8210 27792
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4843 15332 4909 15333
rect 4843 15268 4844 15332
rect 4908 15268 4909 15332
rect 4843 15267 4909 15268
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4846 11933 4906 15267
rect 4843 11932 4909 11933
rect 4843 11868 4844 11932
rect 4908 11868 4909 11932
rect 4843 11867 4909 11868
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4846 10709 4906 11867
rect 5398 11797 5458 17987
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 5395 11796 5461 11797
rect 5395 11732 5396 11796
rect 5460 11732 5461 11796
rect 5395 11731 5461 11732
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 4843 10708 4909 10709
rect 4843 10644 4844 10708
rect 4908 10644 4909 10708
rect 4843 10643 4909 10644
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 27232 15156 27792
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 21782 27232 22102 27792
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 22875 12340 22941 12341
rect 22875 12276 22876 12340
rect 22940 12276 22941 12340
rect 22875 12275 22941 12276
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 20667 8668 20733 8669
rect 20667 8604 20668 8668
rect 20732 8604 20733 8668
rect 20667 8603 20733 8604
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 17907 7036 17973 7037
rect 17907 6972 17908 7036
rect 17972 6972 17973 7036
rect 17907 6971 17973 6972
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 17910 2005 17970 6971
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 20670 4725 20730 8603
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 22878 6221 22938 12275
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 24715 11388 24781 11389
rect 24715 11324 24716 11388
rect 24780 11324 24781 11388
rect 24715 11323 24781 11324
rect 23427 7036 23493 7037
rect 23427 6972 23428 7036
rect 23492 6972 23493 7036
rect 23427 6971 23493 6972
rect 22875 6220 22941 6221
rect 22875 6156 22876 6220
rect 22940 6156 22941 6220
rect 22875 6155 22941 6156
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 20667 4724 20733 4725
rect 20667 4660 20668 4724
rect 20732 4660 20733 4724
rect 20667 4659 20733 4660
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 23430 2413 23490 6971
rect 24718 5541 24778 11323
rect 25255 10368 25575 11392
rect 28728 27232 29048 27792
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 26003 11116 26069 11117
rect 26003 11052 26004 11116
rect 26068 11052 26069 11116
rect 26003 11051 26069 11052
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25819 9076 25885 9077
rect 25819 9012 25820 9076
rect 25884 9012 25885 9076
rect 25819 9011 25885 9012
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 24899 7172 24965 7173
rect 24899 7108 24900 7172
rect 24964 7108 24965 7172
rect 24899 7107 24965 7108
rect 24902 5541 24962 7107
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 24715 5540 24781 5541
rect 24715 5476 24716 5540
rect 24780 5476 24781 5540
rect 24715 5475 24781 5476
rect 24899 5540 24965 5541
rect 24899 5476 24900 5540
rect 24964 5476 24965 5540
rect 24899 5475 24965 5476
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25822 3909 25882 9011
rect 26006 3909 26066 11051
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 25819 3908 25885 3909
rect 25819 3844 25820 3908
rect 25884 3844 25885 3908
rect 25819 3843 25885 3844
rect 26003 3908 26069 3909
rect 26003 3844 26004 3908
rect 26068 3844 26069 3908
rect 26003 3843 26069 3844
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 23427 2412 23493 2413
rect 23427 2348 23428 2412
rect 23492 2348 23493 2412
rect 23427 2347 23493 2348
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 2128 25575 2688
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
rect 17907 2004 17973 2005
rect 17907 1940 17908 2004
rect 17972 1940 17973 2004
rect 17907 1939 17973 1940
use sky130_fd_sc_hd__clkinv_4  _0928_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19044 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0929_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0930_
timestamp 1688980957
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0932_
timestamp 1688980957
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1688980957
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1688980957
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0937_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1688980957
transform 1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0942_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1688980957
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0944_
timestamp 1688980957
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1688980957
transform 1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1688980957
transform 1 0 14168 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1688980957
transform 1 0 16468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1688980957
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1688980957
transform 1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0956_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1688980957
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0958_
timestamp 1688980957
transform 1 0 18032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1688980957
transform 1 0 24748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1688980957
transform 1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1688980957
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1688980957
transform 1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0969_
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1688980957
transform 1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1688980957
transform 1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1688980957
transform 1 0 22172 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1688980957
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1688980957
transform 1 0 24104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1688980957
transform 1 0 23000 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1688980957
transform 1 0 23000 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1688980957
transform 1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1688980957
transform 1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1688980957
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1688980957
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1688980957
transform 1 0 20976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1688980957
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1688980957
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1688980957
transform 1 0 23552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1688980957
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1012_
timestamp 1688980957
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1013_
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1688980957
transform 1 0 17020 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1688980957
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1688980957
transform 1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1688980957
transform 1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1024_
timestamp 1688980957
transform 1 0 17572 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1688980957
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1688980957
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1688980957
transform 1 0 17940 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1688980957
transform 1 0 16652 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1688980957
transform 1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1688980957
transform 1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1688980957
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1688980957
transform 1 0 19596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 1688980957
transform 1 0 19872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1688980957
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1688980957
transform 1 0 21344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1688980957
transform 1 0 21344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1688980957
transform 1 0 21528 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1688980957
transform 1 0 19688 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1688980957
transform 1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1688980957
transform 1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1688980957
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1688980957
transform 1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1688980957
transform 1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1067_
timestamp 1688980957
transform 1 0 28060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1688980957
transform 1 0 27232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1069_
timestamp 1688980957
transform 1 0 27232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1071_
timestamp 1688980957
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1688980957
transform 1 0 27048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1073_
timestamp 1688980957
transform 1 0 21896 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1688980957
transform 1 0 27784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1688980957
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1688980957
transform 1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1688980957
transform 1 0 28336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1688980957
transform 1 0 27416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1688980957
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1688980957
transform 1 0 26128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1091_
timestamp 1688980957
transform 1 0 24656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1688980957
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1093_
timestamp 1688980957
transform 1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1096_
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1688980957
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1688980957
transform 1 0 25668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1688980957
transform 1 0 23092 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1688980957
transform 1 0 24932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1688980957
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1688980957
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1688980957
transform 1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1113_
timestamp 1688980957
transform 1 0 26036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1688980957
transform 1 0 27232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1688980957
transform 1 0 28336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1688980957
transform 1 0 28336 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1117_
timestamp 1688980957
transform 1 0 28336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1119_
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1120_
timestamp 1688980957
transform 1 0 27232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1121_
timestamp 1688980957
transform 1 0 28060 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1688980957
transform 1 0 26956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1688980957
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1688980957
transform 1 0 26680 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1688980957
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1127_
timestamp 1688980957
transform 1 0 24656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1134_
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1688980957
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1688980957
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1142_
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1144_
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1688980957
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1688980957
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1150_
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1152_
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1154_
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1688980957
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1688980957
transform 1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1688980957
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1158_
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1688980957
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1161_
timestamp 1688980957
transform 1 0 1472 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1162_
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1688980957
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1688980957
transform 1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1167_
timestamp 1688980957
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1688980957
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1688980957
transform 1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1688980957
transform 1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1688980957
transform 1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1180_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1688980957
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1688980957
transform 1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1688980957
transform 1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1688980957
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1688980957
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1688980957
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1688980957
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1688980957
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1210_
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1688980957
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1688980957
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1216_
timestamp 1688980957
transform 1 0 11592 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1688980957
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1218_
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1221_
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1688980957
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1688980957
transform 1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1228_
timestamp 1688980957
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1234_
timestamp 1688980957
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1235_
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1688980957
transform 1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1238_
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1240_
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1243_
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1244_
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1248_
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1250_
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1688980957
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1254_
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1688980957
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1259_
timestamp 1688980957
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1688980957
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1688980957
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1265_
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1688980957
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1267_
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1268_
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1269_
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1688980957
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1688980957
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1688980957
transform 1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1275_
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1688980957
transform 1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1688980957
transform 1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1280_
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1282_
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1688980957
transform 1 0 15364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1688980957
transform 1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1688980957
transform 1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1288_
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1289_
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1688980957
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1293_
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1688980957
transform 1 0 14996 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1296_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1688980957
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1688980957
transform 1 0 23368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1305_
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1688980957
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1308_
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1309_
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1310_
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1311_
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1312_
timestamp 1688980957
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1688980957
transform 1 0 17020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1688980957
transform 1 0 17296 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1688980957
transform 1 0 7636 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1316_
timestamp 1688980957
transform 1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1688980957
transform 1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1318_
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1688980957
transform 1 0 4600 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1688980957
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1321_
timestamp 1688980957
transform 1 0 2852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1688980957
transform 1 0 2392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1688980957
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1324_
timestamp 1688980957
transform 1 0 2760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1328_
timestamp 1688980957
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1330_
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1688980957
transform 1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1688980957
transform 1 0 3128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1333_
timestamp 1688980957
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 1688980957
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1688980957
transform 1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1336_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 1688980957
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338_
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 1688980957
transform 1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1340_
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1688980957
transform 1 0 8280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1342_
timestamp 1688980957
transform 1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1688980957
transform 1 0 5152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 1688980957
transform 1 0 6348 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1345_
timestamp 1688980957
transform 1 0 4600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1346_
timestamp 1688980957
transform 1 0 5428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1347_
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1348_
timestamp 1688980957
transform 1 0 6624 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1349_
timestamp 1688980957
transform 1 0 2208 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1351_
timestamp 1688980957
transform 1 0 3220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 1688980957
transform 1 0 4324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1354_
timestamp 1688980957
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 1688980957
transform 1 0 1748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1688980957
transform 1 0 2392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1688980957
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1359_
timestamp 1688980957
transform 1 0 5704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1688980957
transform 1 0 5704 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361_
timestamp 1688980957
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1688980957
transform 1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 1688980957
transform 1 0 7636 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1688980957
transform 1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1688980957
transform 1 0 6532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1688980957
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370_
timestamp 1688980957
transform 1 0 7360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1688980957
transform 1 0 8004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1688980957
transform 1 0 7452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374_
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1688980957
transform 1 0 4232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1688980957
transform 1 0 4968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379_
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380_
timestamp 1688980957
transform 1 0 4784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1688980957
transform 1 0 3404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1383_
timestamp 1688980957
transform 1 0 5060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1384_
timestamp 1688980957
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1385_
timestamp 1688980957
transform 1 0 5704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1688980957
transform 1 0 4968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1387_
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388_
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1390_
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1688980957
transform 1 0 3864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1393_
timestamp 1688980957
transform 1 0 2944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1394_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1688980957
transform 1 0 3680 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1396_
timestamp 1688980957
transform 1 0 7820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1397_
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1688980957
transform 1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1400_
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1402_
timestamp 1688980957
transform 1 0 13064 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1403_
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1404_
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1688980957
transform 1 0 11592 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1406_
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1407_
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1409_
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1411_
timestamp 1688980957
transform 1 0 11592 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412_
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1688980957
transform 1 0 11592 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1415_
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1688980957
transform 1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1418_
timestamp 1688980957
transform 1 0 8464 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1419_
timestamp 1688980957
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1420_
timestamp 1688980957
transform 1 0 9936 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1421_
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1423_
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1688980957
transform 1 0 8924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1425_
timestamp 1688980957
transform 1 0 10212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1426_
timestamp 1688980957
transform 1 0 7544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1688980957
transform 1 0 7820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1429_
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1430_
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1431_
timestamp 1688980957
transform 1 0 9016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1432_
timestamp 1688980957
transform 1 0 6992 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1688980957
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1434_
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1435_
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1438_
timestamp 1688980957
transform 1 0 7268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1440_
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1441_
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1442_
timestamp 1688980957
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1688980957
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1444_
timestamp 1688980957
transform 1 0 3128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1688980957
transform 1 0 12972 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1446_
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1448_
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1451_
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1452_
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1455_
timestamp 1688980957
transform 1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1456_
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1688980957
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1460_
timestamp 1688980957
transform 1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1461_
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1462_
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1688980957
transform 1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1464_
timestamp 1688980957
transform 1 0 13524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1465_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1466_
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1688980957
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1688980957
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1473_
timestamp 1688980957
transform 1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1474_
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1476_
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1477_
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1478_
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1688980957
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1688980957
transform 1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1688980957
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1483_
timestamp 1688980957
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1484_
timestamp 1688980957
transform 1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1688980957
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1688980957
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1490_
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1491_
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1492_
timestamp 1688980957
transform 1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1493_
timestamp 1688980957
transform 1 0 6992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1688980957
transform 1 0 7636 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1495_
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1497_
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1498_
timestamp 1688980957
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1499_
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1688980957
transform 1 0 5152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1501_
timestamp 1688980957
transform 1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1502_
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 1688980957
transform 1 0 22540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1505_
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1506_
timestamp 1688980957
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1508_
timestamp 1688980957
transform 1 0 15180 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1509_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1510_
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1511_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1688980957
transform 1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1513_
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1514_
timestamp 1688980957
transform 1 0 16928 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1515_
timestamp 1688980957
transform 1 0 16100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1688980957
transform 1 0 18676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1688980957
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1519_
timestamp 1688980957
transform 1 0 18584 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1520_
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1521_
timestamp 1688980957
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1688980957
transform 1 0 17296 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1524_
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1525_
timestamp 1688980957
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1688980957
transform 1 0 16100 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1528_
timestamp 1688980957
transform 1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1529_
timestamp 1688980957
transform 1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1688980957
transform 1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1688980957
transform 1 0 28336 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1532_
timestamp 1688980957
transform 1 0 28060 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1688980957
transform 1 0 27692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1534_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1535_
timestamp 1688980957
transform 1 0 24656 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1688980957
transform 1 0 25392 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1537_
timestamp 1688980957
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1538_
timestamp 1688980957
transform 1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1688980957
transform 1 0 27416 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1688980957
transform 1 0 25668 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1688980957
transform 1 0 25576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1544_
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1688980957
transform 1 0 24656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1688980957
transform 1 0 25024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1688980957
transform 1 0 27048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1688980957
transform 1 0 26772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1688980957
transform 1 0 23920 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1554_
timestamp 1688980957
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1688980957
transform 1 0 25024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1556_
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1557_
timestamp 1688980957
transform 1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1558_
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1688980957
transform 1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1560_
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1688980957
transform 1 0 24288 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1562_
timestamp 1688980957
transform 1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1688980957
transform 1 0 25760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1564_
timestamp 1688980957
transform 1 0 24932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1688980957
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1566_
timestamp 1688980957
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1567_
timestamp 1688980957
transform 1 0 18400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1568_
timestamp 1688980957
transform 1 0 17204 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1569_
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1688980957
transform 1 0 14168 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 1688980957
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 1688980957
transform 1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1576_
timestamp 1688980957
transform 1 0 14352 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1577_
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1578_
timestamp 1688980957
transform 1 0 24380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1688980957
transform 1 0 23552 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1688980957
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1583_
timestamp 1688980957
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1584_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1585_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1688980957
transform 1 0 22080 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1589_
timestamp 1688980957
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1590_
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1591_
timestamp 1688980957
transform 1 0 19780 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1592_
timestamp 1688980957
transform 1 0 20056 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1688980957
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1594_
timestamp 1688980957
transform 1 0 22356 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1595_
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1596_
timestamp 1688980957
transform 1 0 20240 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1597_
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1598_
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1688980957
transform 1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1601_
timestamp 1688980957
transform 1 0 23736 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1602_
timestamp 1688980957
transform 1 0 23368 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1603_
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1604_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1605_
timestamp 1688980957
transform 1 0 22632 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1606_
timestamp 1688980957
transform 1 0 22448 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1607_
timestamp 1688980957
transform 1 0 21896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1608_
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1609_
timestamp 1688980957
transform 1 0 22172 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1610_
timestamp 1688980957
transform 1 0 23092 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1613_
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1615_
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1616_
timestamp 1688980957
transform 1 0 22264 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1617_
timestamp 1688980957
transform 1 0 22356 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1688980957
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1619_
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1620_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1621_
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1625_
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1688980957
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1627_
timestamp 1688980957
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1628_
timestamp 1688980957
transform 1 0 18768 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1629_
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1630_
timestamp 1688980957
transform 1 0 16192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1688980957
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1632_
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1633_
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1635_
timestamp 1688980957
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1636_
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1637_
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1638_
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1639_
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1640_
timestamp 1688980957
transform 1 0 13616 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1642_
timestamp 1688980957
transform 1 0 13248 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1643_
timestamp 1688980957
transform 1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1644_
timestamp 1688980957
transform 1 0 13156 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1688980957
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1646_
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1647_
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1688980957
transform 1 0 17204 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1688980957
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1650_
timestamp 1688980957
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1652_
timestamp 1688980957
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1654_
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1688980957
transform 1 0 16192 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1656_
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1657_
timestamp 1688980957
transform 1 0 14904 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1658_
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1659_
timestamp 1688980957
transform 1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1688980957
transform 1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1662_
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1688980957
transform 1 0 15180 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1664_
timestamp 1688980957
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1688980957
transform 1 0 17204 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1666_
timestamp 1688980957
transform 1 0 14628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1688980957
transform 1 0 14904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1668_
timestamp 1688980957
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1669_
timestamp 1688980957
transform 1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1688980957
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1688980957
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1673_
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1688980957
transform 1 0 11040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1675_
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1688980957
transform 1 0 9384 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1677_
timestamp 1688980957
transform 1 0 11776 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1679_
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1681_
timestamp 1688980957
transform 1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1682_
timestamp 1688980957
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1688980957
transform 1 0 9752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1688980957
transform 1 0 6624 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1687_
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1688980957
transform 1 0 8280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1688980957
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1690_
timestamp 1688980957
transform 1 0 8004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1688980957
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1688980957
transform 1 0 8004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1688980957
transform 1 0 11592 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1688980957
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1697_
timestamp 1688980957
transform 1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1698_
timestamp 1688980957
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1700_
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1701_
timestamp 1688980957
transform 1 0 8280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1702_
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1703_
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1704_
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1708_
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1711_
timestamp 1688980957
transform 1 0 9752 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1688980957
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1713_
timestamp 1688980957
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1688980957
transform 1 0 9476 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1715_
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1716_
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1717_
timestamp 1688980957
transform 1 0 21344 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1718_
timestamp 1688980957
transform 1 0 22080 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1688980957
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1688980957
transform 1 0 7636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1721_
timestamp 1688980957
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1722_
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1723_
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1725_
timestamp 1688980957
transform 1 0 3956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1727_
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1728_
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1729_
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1730_
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1731_
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1732_
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1733_
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1734_
timestamp 1688980957
transform 1 0 7636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1735_
timestamp 1688980957
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1736_
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1738_
timestamp 1688980957
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1739_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1740_
timestamp 1688980957
transform 1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1741_
timestamp 1688980957
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1742_
timestamp 1688980957
transform 1 0 7544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1743_
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1688980957
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1745_
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1746_
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1688980957
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1748_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1749_
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1750_
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1752_
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1753_
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1754_
timestamp 1688980957
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1688980957
transform 1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1756_
timestamp 1688980957
transform 1 0 6532 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1758_
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1759_
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1761_
timestamp 1688980957
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1762_
timestamp 1688980957
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1763_
timestamp 1688980957
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1688980957
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1688980957
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1766_
timestamp 1688980957
transform 1 0 16744 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1767_
timestamp 1688980957
transform 1 0 17204 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1768_
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1769_
timestamp 1688980957
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1770_
timestamp 1688980957
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1771_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1772_
timestamp 1688980957
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1773_
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1774_
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1775_
timestamp 1688980957
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1776_
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1777_
timestamp 1688980957
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1778_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1779_
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1780_
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1781_
timestamp 1688980957
transform 1 0 19596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1782_
timestamp 1688980957
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1688980957
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1784_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1785_
timestamp 1688980957
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1787_
timestamp 1688980957
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1788_
timestamp 1688980957
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1789_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1790_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1791_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1792_
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp 1688980957
transform 1 0 7176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1794_
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1795_
timestamp 1688980957
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1796_
timestamp 1688980957
transform 1 0 16744 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1797_
timestamp 1688980957
transform 1 0 27876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1798_
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1799_
timestamp 1688980957
transform 1 0 27600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1800_
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1802_
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1803_
timestamp 1688980957
transform 1 0 28336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1804_
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1805_
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1806_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1807_
timestamp 1688980957
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1809_
timestamp 1688980957
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1810_
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1811_
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1813_
timestamp 1688980957
transform 1 0 26956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1814_
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1815_
timestamp 1688980957
transform 1 0 24472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1816_
timestamp 1688980957
transform 1 0 21620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1817_
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1818_
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1819_
timestamp 1688980957
transform 1 0 26128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1820_
timestamp 1688980957
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1821_
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp 1688980957
transform 1 0 23920 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1823_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1824_
timestamp 1688980957
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1825_
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1826_
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1827_
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1828_
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1829_
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1831_
timestamp 1688980957
transform 1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1832_
timestamp 1688980957
transform 1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1833_
timestamp 1688980957
transform 1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1835_
timestamp 1688980957
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1836_
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp 1688980957
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1838_
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1839_
timestamp 1688980957
transform 1 0 1564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1840_
timestamp 1688980957
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1841_
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1842_
timestamp 1688980957
transform 1 0 28244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1843_
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1845_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1846_
timestamp 1688980957
transform 1 0 14444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1688980957
transform 1 0 14168 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1848_
timestamp 1688980957
transform 1 0 15824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1849_
timestamp 1688980957
transform 1 0 12052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1850_
timestamp 1688980957
transform 1 0 14444 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1851_
timestamp 1688980957
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1852_
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1853_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1854_
timestamp 1688980957
transform 1 0 19504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1855_
timestamp 1688980957
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1856_
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1857_
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1858_
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1859_
timestamp 1688980957
transform 1 0 21344 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1860_
timestamp 1688980957
transform 1 0 28060 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1861_
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1862_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1863_
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1864_
timestamp 1688980957
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1865_
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1866_
timestamp 1688980957
transform 1 0 3128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1867_
timestamp 1688980957
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1868_
timestamp 1688980957
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1869_
timestamp 1688980957
transform 1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1870_
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1871_
timestamp 1688980957
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1872_
timestamp 1688980957
transform 1 0 2300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1873_
timestamp 1688980957
transform 1 0 2576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp 1688980957
transform 1 0 2852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1875_
timestamp 1688980957
transform 1 0 3772 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp 1688980957
transform 1 0 4600 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1877_
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1878_
timestamp 1688980957
transform 1 0 1564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1879_
timestamp 1688980957
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1688980957
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1881_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1882_
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1883_
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1884_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1885_
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1886_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1888_
timestamp 1688980957
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1889_
timestamp 1688980957
transform 1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1890_
timestamp 1688980957
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1891_
timestamp 1688980957
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1892_
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1893_
timestamp 1688980957
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1894_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1895_
timestamp 1688980957
transform 1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1896_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1897_
timestamp 1688980957
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1688980957
transform 1 0 28244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1901_
timestamp 1688980957
transform 1 0 19320 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1688980957
transform 1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1903_
timestamp 1688980957
transform 1 0 16744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1688980957
transform 1 0 24472 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1688980957
transform 1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1906_
timestamp 1688980957
transform 1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1907_
timestamp 1688980957
transform 1 0 21068 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1908_
timestamp 1688980957
transform 1 0 16192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1909_
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1910_
timestamp 1688980957
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1911_
timestamp 1688980957
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1912_
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1688980957
transform 1 0 25392 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1914_
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1915_
timestamp 1688980957
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1916_
timestamp 1688980957
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1917_
timestamp 1688980957
transform 1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1918_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1688980957
transform 1 0 21160 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1688980957
transform 1 0 21896 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1688980957
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1688980957
transform 1 0 25392 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1688980957
transform 1 0 27140 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1688980957
transform 1 0 27140 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1688980957
transform 1 0 26404 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1688980957
transform 1 0 24932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1688980957
transform 1 0 25392 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1688980957
transform 1 0 25300 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1688980957
transform 1 0 25208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1688980957
transform 1 0 27140 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1688980957
transform 1 0 27140 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1688980957
transform 1 0 19688 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfbbn_1  _1936_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1688980957
transform 1 0 23460 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1938_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24656 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1688980957
transform 1 0 25944 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1942_
timestamp 1688980957
transform 1 0 20056 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1946_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1688980957
transform 1 0 17480 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1950_
timestamp 1688980957
transform 1 0 9016 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1688980957
transform 1 0 10304 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1688980957
transform 1 0 7360 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1954_
timestamp 1688980957
transform 1 0 5796 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1688980957
transform 1 0 5060 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1958_
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1962_
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1688980957
transform 1 0 13248 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1688980957
transform 1 0 4784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1966_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1688980957
transform 1 0 6900 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1688980957
transform 1 0 6716 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1970_
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1688980957
transform 1 0 2668 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1688980957
transform 1 0 11316 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1974_
timestamp 1688980957
transform 1 0 11408 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1688980957
transform 1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1978_
timestamp 1688980957
transform 1 0 14352 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1688980957
transform 1 0 11776 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1981_
timestamp 1688980957
transform 1 0 19320 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1982_
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1983_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1688980957
transform 1 0 17204 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1688980957
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1986_
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1987_
timestamp 1688980957
transform 1 0 22632 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1988_
timestamp 1688980957
transform 1 0 22724 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1989_
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1990_
timestamp 1688980957
transform 1 0 17572 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1688980957
transform 1 0 19596 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1688980957
transform 1 0 21896 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1994_
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1995_
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1996_
timestamp 1688980957
transform 1 0 24656 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1997_
timestamp 1688980957
transform 1 0 21344 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1998_
timestamp 1688980957
transform 1 0 22724 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1999_
timestamp 1688980957
transform 1 0 25392 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2000_
timestamp 1688980957
transform 1 0 25024 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2001_
timestamp 1688980957
transform 1 0 17848 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2002_
timestamp 1688980957
transform 1 0 16560 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2003_
timestamp 1688980957
transform 1 0 15732 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2004_
timestamp 1688980957
transform 1 0 19596 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2005_
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2006_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2007_
timestamp 1688980957
transform 1 0 15088 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2008_
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2009_
timestamp 1688980957
transform 1 0 13248 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2010_
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2011_
timestamp 1688980957
transform 1 0 12512 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2012_
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2013_
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2014_
timestamp 1688980957
transform 1 0 12972 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2015_
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2016_
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfbbn_1  _2017_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  _2018_
timestamp 1688980957
transform 1 0 5060 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2019_
timestamp 1688980957
transform 1 0 6808 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2020_
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1688980957
transform 1 0 2208 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2023_
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2024_
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2025_
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2026_
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2027_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2028_
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2029_
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2030_
timestamp 1688980957
transform 1 0 1656 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2031_
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2032_
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2033_
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2034_
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2035_
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfbbn_1  _2036_
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  _2037_
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2038_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2039_
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2040_
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2041_
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2042_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2043_
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2044_
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2045_
timestamp 1688980957
transform 1 0 2668 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2046_
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2047_
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2048_
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2049_
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2050_
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2051_
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2052_
timestamp 1688980957
transform 1 0 11684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2053_
timestamp 1688980957
transform 1 0 11960 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2054_
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfbbn_1  _2055_
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  _2056_
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2057_
timestamp 1688980957
transform 1 0 19872 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__ebufn_1  _2078_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2079_
timestamp 1688980957
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2080_
timestamp 1688980957
transform 1 0 27232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2081_
timestamp 1688980957
transform 1 0 27876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2082_
timestamp 1688980957
transform 1 0 27048 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2083_
timestamp 1688980957
transform 1 0 25852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2084_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2085_
timestamp 1688980957
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2086_
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2087_
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2088_
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2089_
timestamp 1688980957
transform 1 0 24196 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2090_
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2091_
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2092_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2093_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2094_
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2095_
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2096_
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2097_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2098_
timestamp 1688980957
transform 1 0 22632 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2099_
timestamp 1688980957
transform 1 0 25484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2100_
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2101_
timestamp 1688980957
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2102_
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2103_
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2104_
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2105_
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2106_
timestamp 1688980957
transform 1 0 27140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2107_
timestamp 1688980957
transform 1 0 27324 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2108_
timestamp 1688980957
transform 1 0 27784 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2109_
timestamp 1688980957
transform 1 0 24288 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2110_
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2111_
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2112_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2113_
timestamp 1688980957
transform 1 0 25392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2114_
timestamp 1688980957
transform 1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2115_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2116_
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2117_
timestamp 1688980957
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2118_
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2119__48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2119_
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2120_
timestamp 1688980957
transform 1 0 27876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2121_
timestamp 1688980957
transform 1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2122_
timestamp 1688980957
transform 1 0 27784 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2123_
timestamp 1688980957
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2124_
timestamp 1688980957
transform 1 0 21804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2125_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2126_
timestamp 1688980957
transform 1 0 20148 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2127_
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2128_
timestamp 1688980957
transform 1 0 20700 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2129_
timestamp 1688980957
transform 1 0 22448 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2130_
timestamp 1688980957
transform 1 0 21620 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2131_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2132_
timestamp 1688980957
transform 1 0 21620 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2133_
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2134_
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2135_
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2136_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24932 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2137_
timestamp 1688980957
transform 1 0 20240 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2138_
timestamp 1688980957
transform 1 0 21068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2139_
timestamp 1688980957
transform 1 0 20792 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2140_
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2141_
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2142_
timestamp 1688980957
transform 1 0 20516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2143_
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2144_
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2145_
timestamp 1688980957
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2146_
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2147__49
timestamp 1688980957
transform 1 0 23920 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2147_
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2148_
timestamp 1688980957
transform 1 0 22632 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2149_
timestamp 1688980957
transform 1 0 23644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2150_
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2151_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2152_
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2153_
timestamp 1688980957
transform 1 0 15456 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2154_
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2155_
timestamp 1688980957
transform 1 0 14168 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2156_
timestamp 1688980957
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2157_
timestamp 1688980957
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2158_
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2159_
timestamp 1688980957
transform 1 0 16652 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2160_
timestamp 1688980957
transform 1 0 15180 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2161_
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2162_
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2163_
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1688980957
transform 1 0 18124 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2165_
timestamp 1688980957
transform 1 0 16836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2166_
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2167_
timestamp 1688980957
transform 1 0 15364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2168_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2169_
timestamp 1688980957
transform 1 0 14168 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2170_
timestamp 1688980957
transform 1 0 14260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2171_
timestamp 1688980957
transform 1 0 15456 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2172_
timestamp 1688980957
transform 1 0 16744 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2173_
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2174_
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2175_
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2175__50
timestamp 1688980957
transform 1 0 17020 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2176_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2177_
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2178_
timestamp 1688980957
transform 1 0 18032 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _2179_
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2180_
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2181_
timestamp 1688980957
transform 1 0 9568 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2182_
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2183_
timestamp 1688980957
transform 1 0 8740 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2184_
timestamp 1688980957
transform 1 0 9016 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2185_
timestamp 1688980957
transform 1 0 9936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2186_
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2187_
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2188_
timestamp 1688980957
transform 1 0 9752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2189_
timestamp 1688980957
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2190_
timestamp 1688980957
transform 1 0 11684 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2191_
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2192_
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _2193_
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2194_
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2195_
timestamp 1688980957
transform 1 0 9476 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2196_
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2197_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2198_
timestamp 1688980957
transform 1 0 8280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2199_
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2200_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _2201_
timestamp 1688980957
transform 1 0 10212 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2202_
timestamp 1688980957
transform 1 0 9752 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2203_
timestamp 1688980957
transform 1 0 12328 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2203__51
timestamp 1688980957
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2204_
timestamp 1688980957
transform 1 0 10856 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _2205_
timestamp 1688980957
transform 1 0 11776 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2206_
timestamp 1688980957
transform 1 0 12420 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2207_
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2208_
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2209_
timestamp 1688980957
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2210_
timestamp 1688980957
transform 1 0 7084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2211_
timestamp 1688980957
transform 1 0 7268 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2212_
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2213_
timestamp 1688980957
transform 1 0 3312 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2214_
timestamp 1688980957
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2215_
timestamp 1688980957
transform 1 0 7360 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2216_
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2217_
timestamp 1688980957
transform 1 0 4048 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2218_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2219_
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2220_
timestamp 1688980957
transform 1 0 6440 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2221_
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2222_
timestamp 1688980957
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2223_
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2224_
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2225_
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2226_
timestamp 1688980957
transform 1 0 2668 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2227_
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2228_
timestamp 1688980957
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2229_
timestamp 1688980957
transform 1 0 7360 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2230_
timestamp 1688980957
transform 1 0 4324 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2231__52
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2231_
timestamp 1688980957
transform 1 0 4876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2232_
timestamp 1688980957
transform 1 0 6164 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2233_
timestamp 1688980957
transform 1 0 5428 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2234_
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2235_
timestamp 1688980957
transform 1 0 8740 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2236_
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2237_
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2238_
timestamp 1688980957
transform 1 0 9200 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2239_
timestamp 1688980957
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2240_
timestamp 1688980957
transform 1 0 12144 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2241_
timestamp 1688980957
transform 1 0 11868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2242_
timestamp 1688980957
transform 1 0 9108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2243_
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2244_
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2245_
timestamp 1688980957
transform 1 0 12328 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2246_
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2247_
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2248_
timestamp 1688980957
transform 1 0 10212 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2249_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2250_
timestamp 1688980957
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2251_
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2252_
timestamp 1688980957
transform 1 0 9936 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2253_
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2254_
timestamp 1688980957
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2255_
timestamp 1688980957
transform 1 0 11868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2256_
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2257_
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2258_
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2259__53
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2259_
timestamp 1688980957
transform 1 0 11592 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2260_
timestamp 1688980957
transform 1 0 9568 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2261_
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2262_
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2263_
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2264_
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2265_
timestamp 1688980957
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2266_
timestamp 1688980957
transform 1 0 11684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2267_
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2268_
timestamp 1688980957
transform 1 0 15364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2269_
timestamp 1688980957
transform 1 0 14628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2270_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2271_
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2272_
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2273_
timestamp 1688980957
transform 1 0 15364 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2274_
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2275_
timestamp 1688980957
transform 1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2276_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2277_
timestamp 1688980957
transform 1 0 10764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2278_
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2279_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2280_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2281_
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2282_
timestamp 1688980957
transform 1 0 16100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2283_
timestamp 1688980957
transform 1 0 14628 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2284_
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2285_
timestamp 1688980957
transform 1 0 12420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2286_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2287__54
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2287_
timestamp 1688980957
transform 1 0 15456 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2288_
timestamp 1688980957
transform 1 0 12512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2289_
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2290_
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2291_
timestamp 1688980957
transform 1 0 4508 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2292_
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2293_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2294_
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2295_
timestamp 1688980957
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2296_
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2297_
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2298_
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2299_
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2300_
timestamp 1688980957
transform 1 0 7544 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2301_
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2302_
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2303_
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2304_
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2305_
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2306_
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2307_
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2308_
timestamp 1688980957
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2309_
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2310_
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2311_
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2312_
timestamp 1688980957
transform 1 0 5060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2313_
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2314_
timestamp 1688980957
transform 1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2315_
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2315__55
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2316_
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2317_
timestamp 1688980957
transform 1 0 6716 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2318_
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2319_
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2320_
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2321_
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2322_
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2323_
timestamp 1688980957
transform 1 0 9752 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2324_
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2325_
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2326_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2327_
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2328_
timestamp 1688980957
transform 1 0 4324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2329_
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2330_
timestamp 1688980957
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2331_
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2332_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2333_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2334_
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2335_
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2336_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2337_
timestamp 1688980957
transform 1 0 9016 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2338_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2339_
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2340_
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2341_
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2342_
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2343__56
timestamp 1688980957
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2343_
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2344_
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2345_
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2346_
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2347_
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2348_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2349_
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2350_
timestamp 1688980957
transform 1 0 12512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2351_
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2352_
timestamp 1688980957
transform 1 0 11776 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2353_
timestamp 1688980957
transform 1 0 9108 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2354_
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2355_
timestamp 1688980957
transform 1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2356_
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2357_
timestamp 1688980957
transform 1 0 10212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2358_
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2359_
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2360_
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2361_
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2362_
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2363_
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2364_
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2365_
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2366_
timestamp 1688980957
transform 1 0 12512 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2367_
timestamp 1688980957
transform 1 0 9384 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2368_
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2369_
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2370_
timestamp 1688980957
transform 1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2371__57
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2371_
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2372_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2373_
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2374_
timestamp 1688980957
transform 1 0 9568 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2375_
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2376_
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2377_
timestamp 1688980957
transform 1 0 15364 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2378_
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2379_
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2380_
timestamp 1688980957
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2381_
timestamp 1688980957
transform 1 0 12972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2382_
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2383_
timestamp 1688980957
transform 1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2384_
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2385_
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2386_
timestamp 1688980957
transform 1 0 16836 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2387_
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2388_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2389_
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2390_
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2391_
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2392_
timestamp 1688980957
transform 1 0 14628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2393_
timestamp 1688980957
transform 1 0 14352 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2394_
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2395_
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2396_
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2397_
timestamp 1688980957
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2398_
timestamp 1688980957
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2399__58
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2399_
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2400_
timestamp 1688980957
transform 1 0 16100 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2401_
timestamp 1688980957
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2402_
timestamp 1688980957
transform 1 0 13248 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2403_
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2404_
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2405_
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2406_
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2407_
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2408_
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2409_
timestamp 1688980957
transform 1 0 17848 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2410_
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2411_
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2412_
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2413_
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2414_
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2415_
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2416_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2417_
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2418_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2419_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2420_
timestamp 1688980957
transform 1 0 17940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2421_
timestamp 1688980957
transform 1 0 17480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2422_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2423_
timestamp 1688980957
transform 1 0 17112 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2424_
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2425_
timestamp 1688980957
transform 1 0 18676 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2426_
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2427__59
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2427_
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2428_
timestamp 1688980957
transform 1 0 19688 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _2429_
timestamp 1688980957
transform 1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _2430_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2431_
timestamp 1688980957
transform 1 0 21620 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2432_
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2433_
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2434_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2435_
timestamp 1688980957
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2436_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2437_
timestamp 1688980957
transform 1 0 22816 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2438_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2439_
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2440_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2441_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2442_
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2443_
timestamp 1688980957
transform 1 0 25116 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _2444_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2445_
timestamp 1688980957
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2446_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2447_
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2448_
timestamp 1688980957
transform 1 0 21804 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2449_
timestamp 1688980957
transform 1 0 23460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2450_
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2451_
timestamp 1688980957
transform 1 0 22448 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2452_
timestamp 1688980957
transform 1 0 22080 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2453_
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2454_
timestamp 1688980957
transform 1 0 24380 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2455_
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2455__60
timestamp 1688980957
transform 1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2456_
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2457_
timestamp 1688980957
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2458_
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2459_
timestamp 1688980957
transform 1 0 20056 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2460_
timestamp 1688980957
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2461_
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2462_
timestamp 1688980957
transform 1 0 20148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2463_
timestamp 1688980957
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2464_
timestamp 1688980957
transform 1 0 17480 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2465_
timestamp 1688980957
transform 1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2466_
timestamp 1688980957
transform 1 0 20332 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2467_
timestamp 1688980957
transform 1 0 18952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2468_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2469_
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2470_
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2471_
timestamp 1688980957
transform 1 0 20700 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2472_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2473_
timestamp 1688980957
transform 1 0 19320 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2474_
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2475_
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2476_
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2477_
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2478_
timestamp 1688980957
transform 1 0 17296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2479_
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2480_
timestamp 1688980957
transform 1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2481_
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2482_
timestamp 1688980957
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2483_
timestamp 1688980957
transform 1 0 20516 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2483__61
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2484_
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2485_
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2486_
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2487_
timestamp 1688980957
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2488_
timestamp 1688980957
transform 1 0 22356 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2489_
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2490_
timestamp 1688980957
transform 1 0 23000 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2491_
timestamp 1688980957
transform 1 0 26220 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2492_
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2493_
timestamp 1688980957
transform 1 0 26680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2494_
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2495_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2496_
timestamp 1688980957
transform 1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2497_
timestamp 1688980957
transform 1 0 27324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2498_
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2499_
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2500_
timestamp 1688980957
transform 1 0 25576 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2501_
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2502_
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2503_
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2504_
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2505_
timestamp 1688980957
transform 1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2506_
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2507_
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2508_
timestamp 1688980957
transform 1 0 24932 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2509_
timestamp 1688980957
transform 1 0 23920 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2510_
timestamp 1688980957
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2511__62
timestamp 1688980957
transform 1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2511_
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2512_
timestamp 1688980957
transform 1 0 24380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2513_
timestamp 1688980957
transform 1 0 27508 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2514_
timestamp 1688980957
transform 1 0 26680 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2515_
timestamp 1688980957
transform 1 0 23184 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2516_
timestamp 1688980957
transform 1 0 22908 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2517_
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2518_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2519_
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2520_
timestamp 1688980957
transform 1 0 25576 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2521_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2522_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2523_
timestamp 1688980957
transform 1 0 25852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2524_
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2525_
timestamp 1688980957
transform 1 0 27416 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2526_
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2527_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2528_
timestamp 1688980957
transform 1 0 25024 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2529_
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2530_
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2531_
timestamp 1688980957
transform 1 0 24196 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2532_
timestamp 1688980957
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2533_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2534_
timestamp 1688980957
transform 1 0 24840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2535_
timestamp 1688980957
transform 1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2536_
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2537_
timestamp 1688980957
transform 1 0 25668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2538_
timestamp 1688980957
transform 1 0 25944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2539__63
timestamp 1688980957
transform 1 0 28336 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2539_
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2540_
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2541_
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2542_
timestamp 1688980957
transform 1 0 26404 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _2543_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2544__64
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2544_
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2545_
timestamp 1688980957
transform 1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2546_
timestamp 1688980957
transform 1 0 14260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2547_
timestamp 1688980957
transform 1 0 15088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2548_
timestamp 1688980957
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2549_
timestamp 1688980957
transform 1 0 16376 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2550_
timestamp 1688980957
transform 1 0 17848 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2551_
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2552_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2553_
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2554_
timestamp 1688980957
transform 1 0 15364 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2555_
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2556_
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2557_
timestamp 1688980957
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2558_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2559_
timestamp 1688980957
transform 1 0 18952 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2560_
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2561_
timestamp 1688980957
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2562_
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2563_
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2564_
timestamp 1688980957
transform 1 0 17112 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2565_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2566_
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2567_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2568_
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2569_
timestamp 1688980957
transform 1 0 16100 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2570_
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2571_
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2572_
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2573_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _2574_
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  _2575_
timestamp 1688980957
transform 1 0 6440 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2576_
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _2577_
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2578__65
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2578_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2579_
timestamp 1688980957
transform 1 0 2024 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2580_
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2581_
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2582_
timestamp 1688980957
transform 1 0 2944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2583_
timestamp 1688980957
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2584_
timestamp 1688980957
transform 1 0 2576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2585_
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2586_
timestamp 1688980957
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2587_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2588_
timestamp 1688980957
transform 1 0 4140 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2589_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2590_
timestamp 1688980957
transform 1 0 3956 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2591_
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2592_
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2593_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2594_
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2595_
timestamp 1688980957
transform 1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2596_
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2597_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2598_
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2599_
timestamp 1688980957
transform 1 0 3312 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2600_
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2601_
timestamp 1688980957
transform 1 0 3772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2602_
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2603_
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2604_
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2605_
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2606_
timestamp 1688980957
transform 1 0 5520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2607_
timestamp 1688980957
transform 1 0 4876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2608_
timestamp 1688980957
transform 1 0 4784 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2609_
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2610_
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _2611_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2612__66
timestamp 1688980957
transform 1 0 1564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2612_
timestamp 1688980957
transform 1 0 1840 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2613_
timestamp 1688980957
transform 1 0 11408 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2614_
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2615_
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2616_
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2617_
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2618_
timestamp 1688980957
transform 1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2619_
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2620_
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2621_
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2622_
timestamp 1688980957
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2623_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2624_
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2625_
timestamp 1688980957
transform 1 0 9016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2626_
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2627_
timestamp 1688980957
transform 1 0 7268 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2628_
timestamp 1688980957
transform 1 0 10672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2629_
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2630_
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2631_
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2632_
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2633_
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2634_
timestamp 1688980957
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2635_
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2636_
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2637_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2638_
timestamp 1688980957
transform 1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2639_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2640_
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2641_
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2642_
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2643_
timestamp 1688980957
transform 1 0 20240 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  _2644_
timestamp 1688980957
transform 1 0 20976 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _2645_
timestamp 1688980957
transform 1 0 20424 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _2646__67
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2646_
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _2647_
timestamp 1688980957
transform 1 0 27784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2648_
timestamp 1688980957
transform 1 0 26312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2649_
timestamp 1688980957
transform 1 0 26496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2650_
timestamp 1688980957
transform 1 0 27048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2651_
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2652_
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2653_
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2654_
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2655_
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2656_
timestamp 1688980957
transform 1 0 27416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2657_
timestamp 1688980957
transform 1 0 25392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2658_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2659_
timestamp 1688980957
transform 1 0 27048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2660_
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2661_
timestamp 1688980957
transform 1 0 25024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 27968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1688980957
transform 1 0 9844 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1688980957
transform 1 0 10396 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1688980957
transform 1 0 10120 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1688980957
transform 1 0 23644 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1688980957
transform 1 0 24656 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1688980957
transform 1 0 20056 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1688980957
transform 1 0 23184 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1688980957
transform 1 0 23000 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout21
timestamp 1688980957
transform 1 0 15272 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout22
timestamp 1688980957
transform 1 0 11040 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout24
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1688980957
transform 1 0 16928 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout26
timestamp 1688980957
transform 1 0 15272 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1688980957
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1688980957
transform 1 0 27324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1688980957
transform 1 0 6532 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1688980957
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1688980957
transform 1 0 19964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1688980957
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1688980957
transform 1 0 4968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1688980957
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1688980957
transform 1 0 20424 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1688980957
transform 1 0 5244 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1688980957
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_47
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_51
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_152
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_159
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1688980957
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_256
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_260
timestamp 1688980957
transform 1 0 25024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_267
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 1688980957
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_297
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_24
timestamp 1688980957
transform 1 0 3312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_191
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_10
timestamp 1688980957
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_43
timestamp 1688980957
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp 1688980957
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_180
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_202
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_290
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_297
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_32
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_44
timestamp 1688980957
transform 1 0 5152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_63
timestamp 1688980957
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_127
timestamp 1688980957
transform 1 0 12788 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_162
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_219
timestamp 1688980957
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_232
timestamp 1688980957
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_48
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_66
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_172
timestamp 1688980957
transform 1 0 16928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_192
timestamp 1688980957
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_234
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_259
timestamp 1688980957
transform 1 0 24932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 1688980957
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_57
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_105
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_173
timestamp 1688980957
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_237
timestamp 1688980957
transform 1 0 22908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_7
timestamp 1688980957
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_16
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_124
timestamp 1688980957
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_129
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_148
timestamp 1688980957
transform 1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_233
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_297
timestamp 1688980957
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_17
timestamp 1688980957
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_43
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_63
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_72
timestamp 1688980957
transform 1 0 7728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 1688980957
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_100
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_160
timestamp 1688980957
transform 1 0 15824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_182
timestamp 1688980957
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_208
timestamp 1688980957
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_242
timestamp 1688980957
transform 1 0 23368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_259
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_275
timestamp 1688980957
transform 1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_280
timestamp 1688980957
transform 1 0 26864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_298
timestamp 1688980957
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_106
timestamp 1688980957
transform 1 0 10856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_284
timestamp 1688980957
transform 1 0 27232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_297
timestamp 1688980957
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_20
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_116
timestamp 1688980957
transform 1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_186
timestamp 1688980957
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_219
timestamp 1688980957
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_227
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_239
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_275
timestamp 1688980957
transform 1 0 26404 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_292
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_28
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_44
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_52
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_108
timestamp 1688980957
transform 1 0 11040 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_119
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_132 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_144
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_151
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_187
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_236
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_252
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_298
timestamp 1688980957
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_122
timestamp 1688980957
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_152
timestamp 1688980957
transform 1 0 15088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_156
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_188
timestamp 1688980957
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_280
timestamp 1688980957
transform 1 0 26864 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_297
timestamp 1688980957
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_90
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_148
timestamp 1688980957
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_244
timestamp 1688980957
transform 1 0 23552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_270
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_284
timestamp 1688980957
transform 1 0 27232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_297
timestamp 1688980957
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_7
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_42
timestamp 1688980957
transform 1 0 4968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1688980957
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_112
timestamp 1688980957
transform 1 0 11408 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_130
timestamp 1688980957
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_134
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_166
timestamp 1688980957
transform 1 0 16376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_174
timestamp 1688980957
transform 1 0 17112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_181
timestamp 1688980957
transform 1 0 17756 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_205
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_215
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_243
timestamp 1688980957
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_298
timestamp 1688980957
transform 1 0 28520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_102
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_135
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_156
timestamp 1688980957
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1688980957
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_228
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_232
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_262
timestamp 1688980957
transform 1 0 25208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_298
timestamp 1688980957
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_7
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_43
timestamp 1688980957
transform 1 0 5060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_76
timestamp 1688980957
transform 1 0 8096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_98
timestamp 1688980957
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_103
timestamp 1688980957
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_122
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_152
timestamp 1688980957
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_163
timestamp 1688980957
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_175
timestamp 1688980957
transform 1 0 17204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_236
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_241
timestamp 1688980957
transform 1 0 23276 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_278
timestamp 1688980957
transform 1 0 26680 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_68
timestamp 1688980957
transform 1 0 7360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_75
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_85
timestamp 1688980957
transform 1 0 8924 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_91
timestamp 1688980957
transform 1 0 9476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_101
timestamp 1688980957
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 1688980957
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_129
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_133
timestamp 1688980957
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_138
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_157
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_192
timestamp 1688980957
transform 1 0 18768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_204
timestamp 1688980957
transform 1 0 19872 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_241
timestamp 1688980957
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_251
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_298
timestamp 1688980957
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_57
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_69
timestamp 1688980957
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_113
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_131
timestamp 1688980957
transform 1 0 13156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_171
timestamp 1688980957
transform 1 0 16836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_179
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_184
timestamp 1688980957
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_190
timestamp 1688980957
transform 1 0 18584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_213
timestamp 1688980957
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_222
timestamp 1688980957
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_239
timestamp 1688980957
transform 1 0 23092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_287
timestamp 1688980957
transform 1 0 27508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_29
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_86
timestamp 1688980957
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_108
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_139
timestamp 1688980957
transform 1 0 13892 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_155
timestamp 1688980957
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_159
timestamp 1688980957
transform 1 0 15732 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1688980957
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_177
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_184
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_219
timestamp 1688980957
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_259
timestamp 1688980957
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_297
timestamp 1688980957
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_32
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_113
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_166
timestamp 1688980957
transform 1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_175
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_208
timestamp 1688980957
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_212
timestamp 1688980957
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_229
timestamp 1688980957
transform 1 0 22172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_74
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_186
timestamp 1688980957
transform 1 0 18216 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_230
timestamp 1688980957
transform 1 0 22264 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 1688980957
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_40
timestamp 1688980957
transform 1 0 4784 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_44
timestamp 1688980957
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_117
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_192
timestamp 1688980957
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_200
timestamp 1688980957
transform 1 0 19504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_238
timestamp 1688980957
transform 1 0 23000 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_246
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_297
timestamp 1688980957
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_48
timestamp 1688980957
transform 1 0 5520 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_67
timestamp 1688980957
transform 1 0 7268 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_74
timestamp 1688980957
transform 1 0 7912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_99
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_135
timestamp 1688980957
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1688980957
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_184
timestamp 1688980957
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_202
timestamp 1688980957
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_250
timestamp 1688980957
transform 1 0 24104 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_270
timestamp 1688980957
transform 1 0 25944 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_21
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_92
timestamp 1688980957
transform 1 0 9568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_102
timestamp 1688980957
transform 1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_108
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_120
timestamp 1688980957
transform 1 0 12144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_182
timestamp 1688980957
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1688980957
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_257
timestamp 1688980957
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_272
timestamp 1688980957
transform 1 0 26128 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_298
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_34
timestamp 1688980957
transform 1 0 4232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_46
timestamp 1688980957
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_65
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_136
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_178
timestamp 1688980957
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_188
timestamp 1688980957
transform 1 0 18400 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_194
timestamp 1688980957
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_198
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_202
timestamp 1688980957
transform 1 0 19688 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_208
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_251
timestamp 1688980957
transform 1 0 24196 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_269
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_284
timestamp 1688980957
transform 1 0 27232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_297
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_40
timestamp 1688980957
transform 1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_48
timestamp 1688980957
transform 1 0 5520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_61
timestamp 1688980957
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_88
timestamp 1688980957
transform 1 0 9200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_92
timestamp 1688980957
transform 1 0 9568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_101
timestamp 1688980957
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_117
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_127
timestamp 1688980957
transform 1 0 12788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_158
timestamp 1688980957
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_167
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_225
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_258
timestamp 1688980957
transform 1 0 24840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_284
timestamp 1688980957
transform 1 0 27232 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_68
timestamp 1688980957
transform 1 0 7360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_102
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_136
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_143
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_152
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_156
timestamp 1688980957
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_184
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_192
timestamp 1688980957
transform 1 0 18768 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_236
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_248
timestamp 1688980957
transform 1 0 23920 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_258
timestamp 1688980957
transform 1 0 24840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_297
timestamp 1688980957
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_44
timestamp 1688980957
transform 1 0 5152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_56
timestamp 1688980957
transform 1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_99
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_117
timestamp 1688980957
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_124
timestamp 1688980957
transform 1 0 12512 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_132
timestamp 1688980957
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_157
timestamp 1688980957
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_200
timestamp 1688980957
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_218
timestamp 1688980957
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_45
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_94
timestamp 1688980957
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_107
timestamp 1688980957
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_129
timestamp 1688980957
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_133
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_145
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_233
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_238
timestamp 1688980957
transform 1 0 23000 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_263
timestamp 1688980957
transform 1 0 25300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_297
timestamp 1688980957
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_13
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_56
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_144
timestamp 1688980957
transform 1 0 14352 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_152
timestamp 1688980957
transform 1 0 15088 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_163
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_285
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_294
timestamp 1688980957
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_66
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_98
timestamp 1688980957
transform 1 0 10120 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_130
timestamp 1688980957
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_239
timestamp 1688980957
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1688980957
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_297
timestamp 1688980957
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_71
timestamp 1688980957
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_150
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_164
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_170
timestamp 1688980957
transform 1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_268
timestamp 1688980957
transform 1 0 25760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_297
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_25
timestamp 1688980957
transform 1 0 3404 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_78
timestamp 1688980957
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_108
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_129
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_140
timestamp 1688980957
transform 1 0 13984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_180
timestamp 1688980957
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_297
timestamp 1688980957
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_59
timestamp 1688980957
transform 1 0 6532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_164
timestamp 1688980957
transform 1 0 16192 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_184
timestamp 1688980957
transform 1 0 18032 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1688980957
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_216
timestamp 1688980957
transform 1 0 20976 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_262
timestamp 1688980957
transform 1 0 25208 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_274
timestamp 1688980957
transform 1 0 26312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_294
timestamp 1688980957
transform 1 0 28152 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_32
timestamp 1688980957
transform 1 0 4048 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_83
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_140
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_146
timestamp 1688980957
transform 1 0 14536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_179
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_198
timestamp 1688980957
transform 1 0 19320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_207
timestamp 1688980957
transform 1 0 20148 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_242
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_251
timestamp 1688980957
transform 1 0 24196 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_69
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_74
timestamp 1688980957
transform 1 0 7912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_152
timestamp 1688980957
transform 1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_163
timestamp 1688980957
transform 1 0 16100 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_192
timestamp 1688980957
transform 1 0 18768 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_28
timestamp 1688980957
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_122
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_128
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_184
timestamp 1688980957
transform 1 0 18032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_255
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_157
timestamp 1688980957
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_186
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_285
timestamp 1688980957
transform 1 0 27324 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_28
timestamp 1688980957
transform 1 0 3680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_41
timestamp 1688980957
transform 1 0 4876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_46
timestamp 1688980957
transform 1 0 5336 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_76
timestamp 1688980957
transform 1 0 8096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_89
timestamp 1688980957
transform 1 0 9292 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_124
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_141
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_151
timestamp 1688980957
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_175
timestamp 1688980957
transform 1 0 17204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_233
timestamp 1688980957
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_242
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_297
timestamp 1688980957
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_43
timestamp 1688980957
transform 1 0 5060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_63
timestamp 1688980957
transform 1 0 6900 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_90
timestamp 1688980957
transform 1 0 9384 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_136
timestamp 1688980957
transform 1 0 13616 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_152
timestamp 1688980957
transform 1 0 15088 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_161
timestamp 1688980957
transform 1 0 15916 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_166
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_170
timestamp 1688980957
transform 1 0 16744 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_180
timestamp 1688980957
transform 1 0 17664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_192
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_212
timestamp 1688980957
transform 1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_235
timestamp 1688980957
transform 1 0 22724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_242
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 1688980957
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_16
timestamp 1688980957
transform 1 0 2576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_67
timestamp 1688980957
transform 1 0 7268 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_71
timestamp 1688980957
transform 1 0 7636 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_76
timestamp 1688980957
transform 1 0 8096 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_174
timestamp 1688980957
transform 1 0 17112 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_179
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_194
timestamp 1688980957
transform 1 0 18952 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_203
timestamp 1688980957
transform 1 0 19780 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_276
timestamp 1688980957
transform 1 0 26496 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_284
timestamp 1688980957
transform 1 0 27232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_8
timestamp 1688980957
transform 1 0 1840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_171
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_175
timestamp 1688980957
transform 1 0 17204 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_205
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_236
timestamp 1688980957
transform 1 0 22816 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_241
timestamp 1688980957
transform 1 0 23276 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_6
timestamp 1688980957
transform 1 0 1656 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_13
timestamp 1688980957
transform 1 0 2300 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_33
timestamp 1688980957
transform 1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_43
timestamp 1688980957
transform 1 0 5060 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_77
timestamp 1688980957
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_102
timestamp 1688980957
transform 1 0 10488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_178
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_187
timestamp 1688980957
transform 1 0 18308 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_197
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_236
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_256
timestamp 1688980957
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_263
timestamp 1688980957
transform 1 0 25300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_297
timestamp 1688980957
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_22
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_56
timestamp 1688980957
transform 1 0 6256 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_122
timestamp 1688980957
transform 1 0 12328 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_161
timestamp 1688980957
transform 1 0 15916 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_211
timestamp 1688980957
transform 1 0 20516 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_220
timestamp 1688980957
transform 1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_234
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_259
timestamp 1688980957
transform 1 0 24932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_263
timestamp 1688980957
transform 1 0 25300 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_272
timestamp 1688980957
transform 1 0 26128 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_276
timestamp 1688980957
transform 1 0 26496 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_8
timestamp 1688980957
transform 1 0 1840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_49
timestamp 1688980957
transform 1 0 5612 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_65
timestamp 1688980957
transform 1 0 7084 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_91
timestamp 1688980957
transform 1 0 9476 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_131
timestamp 1688980957
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_151
timestamp 1688980957
transform 1 0 14996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_231
timestamp 1688980957
transform 1 0 22356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_267
timestamp 1688980957
transform 1 0 25668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_295
timestamp 1688980957
transform 1 0 28244 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_21
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 1688980957
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_40
timestamp 1688980957
transform 1 0 4784 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_44
timestamp 1688980957
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_73
timestamp 1688980957
transform 1 0 7820 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_96
timestamp 1688980957
transform 1 0 9936 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_111
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_138
timestamp 1688980957
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_156
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_166
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_184
timestamp 1688980957
transform 1 0 18032 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_206
timestamp 1688980957
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_223
timestamp 1688980957
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_225
timestamp 1688980957
transform 1 0 21804 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_232
timestamp 1688980957
transform 1 0 22448 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_240
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_272
timestamp 1688980957
transform 1 0 26128 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_279
timestamp 1688980957
transform 1 0 26772 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 1688980957
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_293
timestamp 1688980957
transform 1 0 28060 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 20148 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 21804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 16744 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 27048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 17020 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 15640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 2668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 1564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 14720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 27508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 1564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 2300 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 1840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 2576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 9936 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 27876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 1472 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 1472 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 7360 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 11684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 6624 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 24748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 12604 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 24104 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 27876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 5336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 22724 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 21620 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 4048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 18032 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform 1 0 27324 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform 1 0 6900 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 4232 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 17020 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 11776 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 24932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 19412 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 20516 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 5428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 26496 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1688980957
transform 1 0 2392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 28336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 3864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 19780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 27324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 26220 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0_subtile_0__pin_I_2_
port 0 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0_subtile_0__pin_I_6_
port 1 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0_subtile_0__pin_O_0_
port 2 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0_subtile_0__pin_clk_0_
port 3 nsew signal input
flabel metal3 s 29200 22040 30000 22160 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 29200 26936 30000 27056 0 FreeSans 480 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 clk
port 6 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 left_width_0_height_0_subtile_0__pin_I_3_
port 7 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 left_width_0_height_0_subtile_0__pin_I_7_
port 8 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 left_width_0_height_0_subtile_0__pin_O_1_
port 9 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 prog_clk
port 10 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 reset
port 11 nsew signal input
flabel metal3 s 29200 2456 30000 2576 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_I_1_
port 12 nsew signal input
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_I_5_
port 13 nsew signal input
flabel metal3 s 29200 12248 30000 12368 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_I_9_
port 14 nsew signal input
flabel metal3 s 29200 17144 30000 17264 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_O_3_
port 15 nsew signal tristate
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 set
port 16 nsew signal input
flabel metal2 s 3790 29200 3846 30000 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_I_0_
port 17 nsew signal input
flabel metal2 s 11242 29200 11298 30000 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_I_4_
port 18 nsew signal input
flabel metal2 s 18694 29200 18750 30000 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_I_8_
port 19 nsew signal input
flabel metal2 s 26146 29200 26202 30000 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_O_2_
port 20 nsew signal tristate
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 1920 90 0 0 vdd
port 21 nsew power bidirectional
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 1920 90 0 0 vdd
port 21 nsew power bidirectional
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 1920 90 0 0 vdd
port 21 nsew power bidirectional
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 1920 90 0 0 vdd
port 21 nsew power bidirectional
flabel metal4 s 7890 2128 8210 27792 0 FreeSans 1920 90 0 0 vss
port 22 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 27792 0 FreeSans 1920 90 0 0 vss
port 22 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 27792 0 FreeSans 1920 90 0 0 vss
port 22 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 27792 0 FreeSans 1920 90 0 0 vss
port 22 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vdd
rlabel via1 15076 27200 15076 27200 0 vss
rlabel metal1 19826 18292 19826 18292 0 _0000_
rlabel metal2 19366 18088 19366 18088 0 _0001_
rlabel metal1 17940 17306 17940 17306 0 _0002_
rlabel metal1 6808 17850 6808 17850 0 _0003_
rlabel metal1 6624 17850 6624 17850 0 _0004_
rlabel metal1 5980 18190 5980 18190 0 _0005_
rlabel metal2 7590 11322 7590 11322 0 _0006_
rlabel metal1 7551 11050 7551 11050 0 _0007_
rlabel metal1 5612 10234 5612 10234 0 _0008_
rlabel metal1 19458 16966 19458 16966 0 _0009_
rlabel metal1 18676 11526 18676 11526 0 _0010_
rlabel metal1 18032 10642 18032 10642 0 _0011_
rlabel metal1 28290 14960 28290 14960 0 _0012_
rlabel metal1 28198 13906 28198 13906 0 _0013_
rlabel metal1 28014 14960 28014 14960 0 _0014_
rlabel metal1 24840 15470 24840 15470 0 _0015_
rlabel metal1 27324 14382 27324 14382 0 _0016_
rlabel metal1 25714 12410 25714 12410 0 _0017_
rlabel metal1 24610 12818 24610 12818 0 _0018_
rlabel metal2 22586 13260 22586 13260 0 _0019_
rlabel metal1 23460 12614 23460 12614 0 _0020_
rlabel metal1 24610 14518 24610 14518 0 _0021_
rlabel metal1 22678 14348 22678 14348 0 _0022_
rlabel metal1 23598 16634 23598 16634 0 _0023_
rlabel metal2 16238 8857 16238 8857 0 _0024_
rlabel metal1 27554 15606 27554 15606 0 _0025_
rlabel metal1 27278 14892 27278 14892 0 _0026_
rlabel metal1 28520 14994 28520 14994 0 _0027_
rlabel metal1 23966 17612 23966 17612 0 _0028_
rlabel metal1 27324 20026 27324 20026 0 _0029_
rlabel metal1 26634 20026 26634 20026 0 _0030_
rlabel metal1 24886 20876 24886 20876 0 _0031_
rlabel metal1 6854 9146 6854 9146 0 _0032_
rlabel metal1 10718 2414 10718 2414 0 _0033_
rlabel metal1 4968 5202 4968 5202 0 _0034_
rlabel metal1 6210 5236 6210 5236 0 _0035_
rlabel metal1 1978 5644 1978 5644 0 _0036_
rlabel metal1 7774 5202 7774 5202 0 _0037_
rlabel metal2 5474 4726 5474 4726 0 _0038_
rlabel metal1 6026 4114 6026 4114 0 _0039_
rlabel metal1 1518 2414 1518 2414 0 _0040_
rlabel metal1 4186 10098 4186 10098 0 _0041_
rlabel metal1 3128 10030 3128 10030 0 _0042_
rlabel metal1 1978 8466 1978 8466 0 _0043_
rlabel metal1 2576 11118 2576 11118 0 _0044_
rlabel metal1 1886 9520 1886 9520 0 _0045_
rlabel metal2 2898 10676 2898 10676 0 _0046_
rlabel metal1 1886 10608 1886 10608 0 _0047_
rlabel metal1 8786 11152 8786 11152 0 _0048_
rlabel metal1 5106 8500 5106 8500 0 _0049_
rlabel metal1 6486 7378 6486 7378 0 _0050_
rlabel metal1 6210 6222 6210 6222 0 _0051_
rlabel metal1 8648 6630 8648 6630 0 _0052_
rlabel metal1 2622 8500 2622 8500 0 _0053_
rlabel metal1 2346 7276 2346 7276 0 _0054_
rlabel metal2 5382 7242 5382 7242 0 _0055_
rlabel metal1 8234 8500 8234 8500 0 _0056_
rlabel metal2 5658 3570 5658 3570 0 _0057_
rlabel metal1 8188 5202 8188 5202 0 _0058_
rlabel metal1 6486 3468 6486 3468 0 _0059_
rlabel metal1 9522 6732 9522 6732 0 _0060_
rlabel metal1 11362 8500 11362 8500 0 _0061_
rlabel metal1 12006 9554 12006 9554 0 _0062_
rlabel metal2 13018 9554 13018 9554 0 _0063_
rlabel metal1 8832 9146 8832 9146 0 _0064_
rlabel metal1 12604 9554 12604 9554 0 _0065_
rlabel viali 11730 10641 11730 10641 0 _0066_
rlabel metal1 10534 11152 10534 11152 0 _0067_
rlabel metal1 11224 7378 11224 7378 0 _0068_
rlabel metal1 12328 6426 12328 6426 0 _0069_
rlabel metal1 12926 6324 12926 6324 0 _0070_
rlabel metal1 11454 5882 11454 5882 0 _0071_
rlabel metal1 10902 5678 10902 5678 0 _0072_
rlabel metal2 8786 6596 8786 6596 0 _0073_
rlabel metal1 9614 5236 9614 5236 0 _0074_
rlabel metal1 9982 4556 9982 4556 0 _0075_
rlabel metal1 9384 4114 9384 4114 0 _0076_
rlabel metal1 13340 5202 13340 5202 0 _0077_
rlabel metal1 14306 3536 14306 3536 0 _0078_
rlabel metal1 13800 5678 13800 5678 0 _0079_
rlabel metal1 14214 10608 14214 10608 0 _0080_
rlabel metal1 14398 9554 14398 9554 0 _0081_
rlabel metal1 15916 8942 15916 8942 0 _0082_
rlabel metal1 15640 10778 15640 10778 0 _0083_
rlabel metal1 14122 10676 14122 10676 0 _0084_
rlabel metal1 18584 4250 18584 4250 0 _0085_
rlabel metal2 15594 7174 15594 7174 0 _0086_
rlabel metal2 14122 7990 14122 7990 0 _0087_
rlabel metal1 15180 7174 15180 7174 0 _0088_
rlabel metal1 16606 5202 16606 5202 0 _0089_
rlabel metal1 16100 6290 16100 6290 0 _0090_
rlabel metal1 14996 5610 14996 5610 0 _0091_
rlabel metal1 11592 4114 11592 4114 0 _0092_
rlabel metal2 23368 2516 23368 2516 0 _0093_
rlabel metal1 17986 2958 17986 2958 0 _0094_
rlabel metal1 18078 2414 18078 2414 0 _0095_
rlabel metal1 20148 8466 20148 8466 0 _0096_
rlabel metal1 17066 8942 17066 8942 0 _0097_
rlabel metal2 4738 21726 4738 21726 0 _0098_
rlabel metal1 2484 22610 2484 22610 0 _0099_
rlabel metal1 2346 24684 2346 24684 0 _0100_
rlabel metal1 3496 21862 3496 21862 0 _0101_
rlabel metal1 2530 25296 2530 25296 0 _0102_
rlabel metal1 4462 20026 4462 20026 0 _0103_
rlabel metal1 2116 22610 2116 22610 0 _0104_
rlabel metal1 4094 19380 4094 19380 0 _0105_
rlabel metal1 3450 20570 3450 20570 0 _0106_
rlabel metal1 5014 25194 5014 25194 0 _0107_
rlabel metal1 6578 26418 6578 26418 0 _0108_
rlabel metal1 4876 26554 4876 26554 0 _0109_
rlabel metal1 2070 25874 2070 25874 0 _0110_
rlabel metal1 2254 26452 2254 26452 0 _0111_
rlabel metal1 4278 25262 4278 25262 0 _0112_
rlabel metal1 2622 25908 2622 25908 0 _0113_
rlabel metal1 5842 26962 5842 26962 0 _0114_
rlabel metal2 4554 25024 4554 25024 0 _0115_
rlabel metal2 6762 25874 6762 25874 0 _0116_
rlabel metal1 4968 21114 4968 21114 0 _0117_
rlabel metal1 7682 24208 7682 24208 0 _0118_
rlabel metal1 4508 24174 4508 24174 0 _0119_
rlabel metal2 5566 21556 5566 21556 0 _0120_
rlabel metal1 3542 22202 3542 22202 0 _0121_
rlabel metal1 5934 19380 5934 19380 0 _0122_
rlabel metal1 3404 17646 3404 17646 0 _0123_
rlabel metal1 5106 17612 5106 17612 0 _0124_
rlabel metal1 3680 16082 3680 16082 0 _0125_
rlabel metal1 9338 20026 9338 20026 0 _0126_
rlabel metal1 13892 19822 13892 19822 0 _0127_
rlabel metal1 13110 20468 13110 20468 0 _0128_
rlabel metal1 7314 17612 7314 17612 0 _0129_
rlabel metal1 11822 18224 11822 18224 0 _0130_
rlabel metal1 12995 17170 12995 17170 0 _0131_
rlabel metal1 11822 16048 11822 16048 0 _0132_
rlabel metal1 10948 15470 10948 15470 0 _0133_
rlabel metal2 10074 19788 10074 19788 0 _0134_
rlabel metal1 9936 17646 9936 17646 0 _0135_
rlabel metal1 9108 15470 9108 15470 0 _0136_
rlabel metal1 8050 17612 8050 17612 0 _0137_
rlabel metal1 9062 18734 9062 18734 0 _0138_
rlabel metal1 7176 17850 7176 17850 0 _0139_
rlabel metal1 8188 17034 8188 17034 0 _0140_
rlabel metal1 4738 18700 4738 18700 0 _0141_
rlabel metal1 3312 14586 3312 14586 0 _0142_
rlabel metal1 13386 14586 13386 14586 0 _0143_
rlabel metal1 14478 16082 14478 16082 0 _0144_
rlabel metal1 16422 13872 16422 13872 0 _0145_
rlabel metal1 9154 13260 9154 13260 0 _0146_
rlabel metal2 13662 13124 13662 13124 0 _0147_
rlabel metal1 16054 12852 16054 12852 0 _0148_
rlabel metal1 16284 11730 16284 11730 0 _0149_
rlabel metal1 13754 11764 13754 11764 0 _0150_
rlabel metal1 12466 12852 12466 12852 0 _0151_
rlabel metal2 12604 12070 12604 12070 0 _0152_
rlabel metal2 10718 12036 10718 12036 0 _0153_
rlabel metal1 11362 12852 11362 12852 0 _0154_
rlabel metal1 11454 13872 11454 13872 0 _0155_
rlabel metal1 10902 15028 10902 15028 0 _0156_
rlabel metal1 9016 12818 9016 12818 0 _0157_
rlabel metal1 4462 14382 4462 14382 0 _0158_
rlabel metal1 8234 14586 8234 14586 0 _0159_
rlabel metal1 7866 15028 7866 15028 0 _0160_
rlabel metal1 6210 14960 6210 14960 0 _0161_
rlabel metal1 6210 17136 6210 17136 0 _0162_
rlabel metal1 5382 17204 5382 17204 0 _0163_
rlabel metal1 23184 19346 23184 19346 0 _0164_
rlabel metal1 15916 22066 15916 22066 0 _0165_
rlabel metal1 16928 21862 16928 21862 0 _0166_
rlabel metal1 18906 23120 18906 23120 0 _0167_
rlabel metal1 16698 24208 16698 24208 0 _0168_
rlabel metal1 18906 24922 18906 24922 0 _0169_
rlabel metal1 17388 24786 17388 24786 0 _0170_
rlabel metal1 17756 25262 17756 25262 0 _0171_
rlabel metal2 16698 26010 16698 26010 0 _0172_
rlabel metal1 28474 25466 28474 25466 0 _0173_
rlabel metal1 28336 24582 28336 24582 0 _0174_
rlabel metal1 28014 25466 28014 25466 0 _0175_
rlabel metal1 23966 21998 23966 21998 0 _0176_
rlabel metal1 25760 27098 25760 27098 0 _0177_
rlabel metal1 25944 24038 25944 24038 0 _0178_
rlabel metal1 25346 24140 25346 24140 0 _0179_
rlabel metal1 25116 25874 25116 25874 0 _0180_
rlabel metal1 27048 23086 27048 23086 0 _0181_
rlabel metal1 27186 22406 27186 22406 0 _0182_
rlabel metal1 24242 22746 24242 22746 0 _0183_
rlabel metal1 25530 21488 25530 21488 0 _0184_
rlabel metal1 26450 21522 26450 21522 0 _0185_
rlabel metal1 24564 20434 24564 20434 0 _0186_
rlabel metal1 25484 20910 25484 20910 0 _0187_
rlabel metal1 19228 24174 19228 24174 0 _0188_
rlabel metal2 12926 27234 12926 27234 0 _0189_
rlabel metal1 15916 24922 15916 24922 0 _0190_
rlabel metal1 14582 25908 14582 25908 0 _0191_
rlabel metal1 24196 24378 24196 24378 0 _0192_
rlabel metal1 23782 26384 23782 26384 0 _0193_
rlabel metal1 24058 26418 24058 26418 0 _0194_
rlabel metal1 22816 22610 22816 22610 0 _0195_
rlabel metal1 22126 27098 22126 27098 0 _0196_
rlabel metal1 22678 25262 22678 25262 0 _0197_
rlabel metal1 20286 25840 20286 25840 0 _0198_
rlabel metal1 20470 26384 20470 26384 0 _0199_
rlabel metal1 24150 23290 24150 23290 0 _0200_
rlabel metal1 23690 22746 23690 22746 0 _0201_
rlabel metal1 21850 21522 21850 21522 0 _0202_
rlabel metal2 23690 23698 23690 23698 0 _0203_
rlabel metal1 23690 22576 23690 22576 0 _0204_
rlabel metal1 22678 21080 22678 21080 0 _0205_
rlabel metal1 20838 21930 20838 21930 0 _0206_
rlabel metal1 18722 24208 18722 24208 0 _0207_
rlabel via1 13570 24162 13570 24162 0 _0208_
rlabel metal1 18170 20944 18170 20944 0 _0209_
rlabel metal1 18216 19958 18216 19958 0 _0210_
rlabel metal1 16698 19856 16698 19856 0 _0211_
rlabel metal1 13800 18734 13800 18734 0 _0212_
rlabel metal1 15134 21488 15134 21488 0 _0213_
rlabel metal1 16008 19346 16008 19346 0 _0214_
rlabel metal1 14306 18700 14306 18700 0 _0215_
rlabel metal1 13662 20468 13662 20468 0 _0216_
rlabel metal1 17434 18258 17434 18258 0 _0217_
rlabel metal1 16882 17204 16882 17204 0 _0218_
rlabel metal1 14214 17204 14214 17204 0 _0219_
rlabel metal1 15134 18224 15134 18224 0 _0220_
rlabel metal1 17710 17204 17710 17204 0 _0221_
rlabel metal1 15318 16082 15318 16082 0 _0222_
rlabel metal1 15134 16116 15134 16116 0 _0223_
rlabel metal1 15456 22610 15456 22610 0 _0224_
rlabel metal1 11224 24582 11224 24582 0 _0225_
rlabel metal1 11408 26962 11408 26962 0 _0226_
rlabel metal2 9706 27710 9706 27710 0 _0227_
rlabel metal1 10258 20774 10258 20774 0 _0228_
rlabel metal1 7038 27472 7038 27472 0 _0229_
rlabel metal1 9292 25398 9292 25398 0 _0230_
rlabel metal1 8786 26316 8786 26316 0 _0231_
rlabel metal1 7406 27098 7406 27098 0 _0232_
rlabel metal1 10810 24854 10810 24854 0 _0233_
rlabel metal1 10074 23290 10074 23290 0 _0234_
rlabel metal1 8326 21896 8326 21896 0 _0235_
rlabel metal1 8970 23698 8970 23698 0 _0236_
rlabel metal2 11868 21998 11868 21998 0 _0237_
rlabel metal1 8602 21896 8602 21896 0 _0238_
rlabel metal1 9384 23086 9384 23086 0 _0239_
rlabel metal2 13938 23018 13938 23018 0 _0240_
rlabel metal2 22218 19958 22218 19958 0 _0241_
rlabel metal1 9062 20468 9062 20468 0 _0242_
rlabel metal1 5474 15028 5474 15028 0 _0243_
rlabel metal1 4554 16116 4554 16116 0 _0244_
rlabel metal1 7314 17204 7314 17204 0 _0245_
rlabel metal1 8234 13498 8234 13498 0 _0246_
rlabel metal1 6486 12410 6486 12410 0 _0247_
rlabel metal1 6072 11322 6072 11322 0 _0248_
rlabel metal1 7452 11866 7452 11866 0 _0249_
rlabel metal1 6210 12852 6210 12852 0 _0250_
rlabel metal1 3910 11118 3910 11118 0 _0251_
rlabel metal1 5704 10642 5704 10642 0 _0252_
rlabel metal1 1978 13260 1978 13260 0 _0253_
rlabel metal1 19090 8908 19090 8908 0 _0254_
rlabel metal1 18354 9996 18354 9996 0 _0255_
rlabel metal1 2024 11118 2024 11118 0 _0256_
rlabel metal1 17112 10030 17112 10030 0 _0257_
rlabel viali 19458 2415 19458 2415 0 _0258_
rlabel metal1 18170 7888 18170 7888 0 _0259_
rlabel metal1 17572 6766 17572 6766 0 _0260_
rlabel metal1 19412 6970 19412 6970 0 _0261_
rlabel metal1 20056 3910 20056 3910 0 _0262_
rlabel metal1 19918 5678 19918 5678 0 _0263_
rlabel metal1 19458 4658 19458 4658 0 _0264_
rlabel metal1 15502 1972 15502 1972 0 _0265_
rlabel metal2 18814 2247 18814 2247 0 _0266_
rlabel metal1 27094 20570 27094 20570 0 _0267_
rlabel metal1 27784 16218 27784 16218 0 _0268_
rlabel metal2 26542 17697 26542 17697 0 _0269_
rlabel metal1 24150 18292 24150 18292 0 _0270_
rlabel metal1 24426 18292 24426 18292 0 _0271_
rlabel metal1 25392 17850 25392 17850 0 _0272_
rlabel metal1 21666 17748 21666 17748 0 _0273_
rlabel metal1 23690 17646 23690 17646 0 _0274_
rlabel metal1 28060 9554 28060 9554 0 _0275_
rlabel metal1 25024 4454 25024 4454 0 _0276_
rlabel metal1 24794 12240 24794 12240 0 _0277_
rlabel metal1 25392 3978 25392 3978 0 _0278_
rlabel metal1 14398 8058 14398 8058 0 _0279_
rlabel metal2 2162 2244 2162 2244 0 _0280_
rlabel metal1 17020 3502 17020 3502 0 _0281_
rlabel metal1 17388 6902 17388 6902 0 _0282_
rlabel metal1 17066 3706 17066 3706 0 _0283_
rlabel metal1 19596 8942 19596 8942 0 _0284_
rlabel metal1 27186 7412 27186 7412 0 _0285_
rlabel metal1 24932 8330 24932 8330 0 _0286_
rlabel metal1 24610 7820 24610 7820 0 _0287_
rlabel metal2 20700 9554 20700 9554 0 _0288_
rlabel metal1 21942 10030 21942 10030 0 _0289_
rlabel metal1 25898 9622 25898 9622 0 _0290_
rlabel metal1 22862 10608 22862 10608 0 _0291_
rlabel metal1 23138 11118 23138 11118 0 _0292_
rlabel metal1 23690 7786 23690 7786 0 _0293_
rlabel metal1 21689 8602 21689 8602 0 _0294_
rlabel metal1 21206 8432 21206 8432 0 _0295_
rlabel metal1 20470 8466 20470 8466 0 _0296_
rlabel metal1 24242 4556 24242 4556 0 _0297_
rlabel metal1 20746 7378 20746 7378 0 _0298_
rlabel metal1 21206 7888 21206 7888 0 _0299_
rlabel metal1 26818 3570 26818 3570 0 _0300_
rlabel metal1 15180 6902 15180 6902 0 _0301_
rlabel metal1 17894 8976 17894 8976 0 _0302_
rlabel metal1 4922 3162 4922 3162 0 _0303_
rlabel metal1 21666 10506 21666 10506 0 _0304_
rlabel metal2 21850 12750 21850 12750 0 _0305_
rlabel metal1 20286 12172 20286 12172 0 _0306_
rlabel metal1 19044 15470 19044 15470 0 _0307_
rlabel metal1 17894 12614 17894 12614 0 _0308_
rlabel metal1 19550 13940 19550 13940 0 _0309_
rlabel metal1 16974 15130 16974 15130 0 _0310_
rlabel metal1 17158 13328 17158 13328 0 _0311_
rlabel metal1 21022 14042 21022 14042 0 _0312_
rlabel metal1 20654 14416 20654 14416 0 _0313_
rlabel metal1 20102 14416 20102 14416 0 _0314_
rlabel metal1 18722 14348 18722 14348 0 _0315_
rlabel metal1 21114 16218 21114 16218 0 _0316_
rlabel metal2 21390 16150 21390 16150 0 _0317_
rlabel metal1 19182 16218 19182 16218 0 _0318_
rlabel metal2 23782 10676 23782 10676 0 _0319_
rlabel metal1 24334 9690 24334 9690 0 _0320_
rlabel metal1 28152 7854 28152 7854 0 _0321_
rlabel metal1 27370 10642 27370 10642 0 _0322_
rlabel metal1 26266 11322 26266 11322 0 _0323_
rlabel metal1 27186 3706 27186 3706 0 _0324_
rlabel metal1 28014 4046 28014 4046 0 _0325_
rlabel metal2 17894 8126 17894 8126 0 _0326_
rlabel metal1 24012 12070 24012 12070 0 _0327_
rlabel metal1 27140 4114 27140 4114 0 _0328_
rlabel metal2 17434 5593 17434 5593 0 _0329_
rlabel metal1 24564 2618 24564 2618 0 _0330_
rlabel metal1 23828 4590 23828 4590 0 _0331_
rlabel metal1 21528 5202 21528 5202 0 _0332_
rlabel metal1 20654 6120 20654 6120 0 _0333_
rlabel metal2 21298 8857 21298 8857 0 _0334_
rlabel metal2 14122 5933 14122 5933 0 _0335_
rlabel via2 16606 6715 16606 6715 0 _0336_
rlabel metal1 25576 2618 25576 2618 0 _0337_
rlabel metal1 24656 6358 24656 6358 0 _0338_
rlabel metal1 19642 18870 19642 18870 0 _0339_
rlabel metal1 20700 18258 20700 18258 0 _0340_
rlabel metal1 23920 21114 23920 21114 0 _0341_
rlabel metal1 23828 20978 23828 20978 0 _0342_
rlabel metal1 24702 22066 24702 22066 0 _0343_
rlabel metal1 23138 21522 23138 21522 0 _0344_
rlabel metal1 25990 25806 25990 25806 0 _0345_
rlabel metal1 25622 24378 25622 24378 0 _0346_
rlabel metal1 26174 26962 26174 26962 0 _0347_
rlabel metal1 26266 22066 26266 22066 0 _0348_
rlabel metal1 26772 21658 26772 21658 0 _0349_
rlabel metal1 26450 24922 26450 24922 0 _0350_
rlabel metal2 27094 25568 27094 25568 0 _0351_
rlabel metal1 27370 22644 27370 22644 0 _0352_
rlabel metal2 27554 24820 27554 24820 0 _0353_
rlabel metal1 28106 23018 28106 23018 0 _0354_
rlabel metal1 24748 21114 24748 21114 0 _0355_
rlabel metal2 24334 20808 24334 20808 0 _0356_
rlabel metal2 25346 21828 25346 21828 0 _0357_
rlabel metal1 23644 23222 23644 23222 0 _0358_
rlabel metal1 25346 26010 25346 26010 0 _0359_
rlabel metal1 25576 24310 25576 24310 0 _0360_
rlabel metal1 26864 26962 26864 26962 0 _0361_
rlabel metal1 25806 21420 25806 21420 0 _0362_
rlabel metal2 27554 22508 27554 22508 0 _0363_
rlabel metal1 26726 24922 26726 24922 0 _0364_
rlabel metal1 27646 26418 27646 26418 0 _0365_
rlabel metal1 27784 22610 27784 22610 0 _0366_
rlabel metal1 28152 25874 28152 25874 0 _0367_
rlabel metal1 28060 24106 28060 24106 0 _0368_
rlabel metal1 21068 21522 21068 21522 0 _0369_
rlabel metal1 22678 20944 22678 20944 0 _0370_
rlabel metal2 22126 23375 22126 23375 0 _0371_
rlabel metal1 20378 22644 20378 22644 0 _0372_
rlabel metal1 21206 26418 21206 26418 0 _0373_
rlabel metal1 21160 25330 21160 25330 0 _0374_
rlabel metal1 22448 26962 22448 26962 0 _0375_
rlabel metal1 21712 22066 21712 22066 0 _0376_
rlabel metal2 22586 23868 22586 23868 0 _0377_
rlabel metal1 22172 26418 22172 26418 0 _0378_
rlabel metal1 24104 26894 24104 26894 0 _0379_
rlabel metal1 22862 23732 22862 23732 0 _0380_
rlabel metal2 23138 25636 23138 25636 0 _0381_
rlabel metal1 25162 23800 25162 23800 0 _0382_
rlabel metal2 20654 21692 20654 21692 0 _0383_
rlabel metal1 21298 20842 21298 20842 0 _0384_
rlabel metal2 21022 24004 21022 24004 0 _0385_
rlabel metal1 21482 21386 21482 21386 0 _0386_
rlabel metal1 20700 26554 20700 26554 0 _0387_
rlabel metal1 20746 25772 20746 25772 0 _0388_
rlabel metal1 23092 26962 23092 26962 0 _0389_
rlabel metal1 23368 21998 23368 21998 0 _0390_
rlabel metal1 21988 23086 21988 23086 0 _0391_
rlabel metal1 22586 25160 22586 25160 0 _0392_
rlabel metal1 24380 26554 24380 26554 0 _0393_
rlabel metal2 22862 23596 22862 23596 0 _0394_
rlabel metal1 23736 25874 23736 25874 0 _0395_
rlabel metal2 24610 25432 24610 25432 0 _0396_
rlabel metal1 15778 16082 15778 16082 0 _0397_
rlabel metal1 16192 16626 16192 16626 0 _0398_
rlabel metal1 15502 18258 15502 18258 0 _0399_
rlabel metal1 14444 17714 14444 17714 0 _0400_
rlabel metal1 14720 20366 14720 20366 0 _0401_
rlabel metal1 15226 19244 15226 19244 0 _0402_
rlabel metal1 15548 21114 15548 21114 0 _0403_
rlabel metal1 17112 16626 17112 16626 0 _0404_
rlabel metal1 16698 17714 16698 17714 0 _0405_
rlabel metal1 15732 20026 15732 20026 0 _0406_
rlabel metal1 16284 20570 16284 20570 0 _0407_
rlabel metal1 17710 17578 17710 17578 0 _0408_
rlabel metal1 17342 19890 17342 19890 0 _0409_
rlabel metal2 18354 19329 18354 19329 0 _0410_
rlabel metal1 16008 15538 16008 15538 0 _0411_
rlabel metal1 15456 15946 15456 15946 0 _0412_
rlabel metal1 15272 18394 15272 18394 0 _0413_
rlabel metal1 14168 17306 14168 17306 0 _0414_
rlabel metal1 14398 19958 14398 19958 0 _0415_
rlabel metal1 14306 18938 14306 18938 0 _0416_
rlabel metal1 15318 20978 15318 20978 0 _0417_
rlabel metal1 17250 16082 17250 16082 0 _0418_
rlabel metal1 16422 17306 16422 17306 0 _0419_
rlabel metal1 15594 19482 15594 19482 0 _0420_
rlabel metal1 16698 20026 16698 20026 0 _0421_
rlabel metal1 18446 17544 18446 17544 0 _0422_
rlabel metal1 17480 20570 17480 20570 0 _0423_
rlabel metal1 18262 20536 18262 20536 0 _0424_
rlabel metal1 10028 21862 10028 21862 0 _0425_
rlabel metal1 10810 20366 10810 20366 0 _0426_
rlabel metal1 9246 24242 9246 24242 0 _0427_
rlabel metal2 8142 22151 8142 22151 0 _0428_
rlabel metal1 8970 26996 8970 26996 0 _0429_
rlabel metal1 8832 25466 8832 25466 0 _0430_
rlabel metal1 10166 27030 10166 27030 0 _0431_
rlabel metal1 10258 22984 10258 22984 0 _0432_
rlabel metal1 10534 23800 10534 23800 0 _0433_
rlabel metal1 9982 26452 9982 26452 0 _0434_
rlabel metal1 10488 26894 10488 26894 0 _0435_
rlabel metal1 11914 23800 11914 23800 0 _0436_
rlabel metal1 10810 25466 10810 25466 0 _0437_
rlabel metal1 12052 23018 12052 23018 0 _0438_
rlabel metal1 10718 21862 10718 21862 0 _0439_
rlabel metal2 8970 21726 8970 21726 0 _0440_
rlabel metal1 9706 23800 9706 23800 0 _0441_
rlabel metal1 6992 21658 6992 21658 0 _0442_
rlabel metal1 8832 26418 8832 26418 0 _0443_
rlabel metal1 8556 25874 8556 25874 0 _0444_
rlabel metal1 10488 27438 10488 27438 0 _0445_
rlabel metal2 11730 22440 11730 22440 0 _0446_
rlabel metal1 10672 22678 10672 22678 0 _0447_
rlabel metal1 9844 25874 9844 25874 0 _0448_
rlabel metal1 12558 27370 12558 27370 0 _0449_
rlabel metal2 11086 23800 11086 23800 0 _0450_
rlabel metal1 11776 27030 11776 27030 0 _0451_
rlabel metal1 12696 25806 12696 25806 0 _0452_
rlabel metal1 4968 22610 4968 22610 0 _0453_
rlabel metal1 4278 21930 4278 21930 0 _0454_
rlabel metal2 8326 23868 8326 23868 0 _0455_
rlabel metal1 7314 22644 7314 22644 0 _0456_
rlabel metal1 6808 26962 6808 26962 0 _0457_
rlabel metal1 3588 25466 3588 25466 0 _0458_
rlabel metal1 3450 26554 3450 26554 0 _0459_
rlabel metal1 5658 23732 5658 23732 0 _0460_
rlabel metal1 7544 23154 7544 23154 0 _0461_
rlabel metal1 7774 26418 7774 26418 0 _0462_
rlabel metal1 4278 27064 4278 27064 0 _0463_
rlabel metal1 6578 23732 6578 23732 0 _0464_
rlabel metal1 5612 26010 5612 26010 0 _0465_
rlabel metal1 6992 24854 6992 24854 0 _0466_
rlabel viali 6210 21999 6210 21999 0 _0467_
rlabel metal1 5382 21862 5382 21862 0 _0468_
rlabel metal1 8510 23596 8510 23596 0 _0469_
rlabel metal1 7912 22610 7912 22610 0 _0470_
rlabel metal1 5750 26860 5750 26860 0 _0471_
rlabel metal1 2599 25738 2599 25738 0 _0472_
rlabel metal2 2714 26792 2714 26792 0 _0473_
rlabel metal1 5152 24378 5152 24378 0 _0474_
rlabel metal1 7406 23698 7406 23698 0 _0475_
rlabel metal2 4002 25602 4002 25602 0 _0476_
rlabel metal1 5290 26962 5290 26962 0 _0477_
rlabel metal1 6624 24242 6624 24242 0 _0478_
rlabel metal1 5888 26282 5888 26282 0 _0479_
rlabel metal1 5704 25466 5704 25466 0 _0480_
rlabel metal1 8188 17850 8188 17850 0 _0481_
rlabel metal1 6302 18122 6302 18122 0 _0482_
rlabel metal1 9016 16762 9016 16762 0 _0483_
rlabel metal1 9246 16082 9246 16082 0 _0484_
rlabel metal1 10948 16762 10948 16762 0 _0485_
rlabel metal1 12190 16014 12190 16014 0 _0486_
rlabel metal1 12098 18292 12098 18292 0 _0487_
rlabel metal1 9476 18394 9476 18394 0 _0488_
rlabel metal1 10028 17102 10028 17102 0 _0489_
rlabel metal1 11914 17170 11914 17170 0 _0490_
rlabel metal2 13202 18836 13202 18836 0 _0491_
rlabel metal1 10488 18190 10488 18190 0 _0492_
rlabel metal1 13156 18802 13156 18802 0 _0493_
rlabel metal1 10074 19414 10074 19414 0 _0494_
rlabel metal1 8786 17714 8786 17714 0 _0495_
rlabel metal2 8326 18428 8326 18428 0 _0496_
rlabel metal1 8234 17204 8234 17204 0 _0497_
rlabel metal1 9752 15674 9752 15674 0 _0498_
rlabel metal1 11040 15334 11040 15334 0 _0499_
rlabel metal1 13110 15946 13110 15946 0 _0500_
rlabel metal1 11868 18394 11868 18394 0 _0501_
rlabel metal1 9062 18904 9062 18904 0 _0502_
rlabel metal1 9844 16626 9844 16626 0 _0503_
rlabel metal1 12834 17068 12834 17068 0 _0504_
rlabel metal2 13754 19720 13754 19720 0 _0505_
rlabel metal1 9844 18802 9844 18802 0 _0506_
rlabel metal1 13478 19890 13478 19890 0 _0507_
rlabel metal2 10994 19992 10994 19992 0 _0508_
rlabel metal1 10258 12716 10258 12716 0 _0509_
rlabel metal1 9798 13430 9798 13430 0 _0510_
rlabel metal2 12926 13158 12926 13158 0 _0511_
rlabel metal2 12834 12070 12834 12070 0 _0512_
rlabel metal1 14260 11730 14260 11730 0 _0513_
rlabel metal1 15732 11866 15732 11866 0 _0514_
rlabel metal1 14674 13362 14674 13362 0 _0515_
rlabel metal1 10856 12614 10856 12614 0 _0516_
rlabel metal2 13478 13090 13478 13090 0 _0517_
rlabel metal1 14674 12274 14674 12274 0 _0518_
rlabel metal1 15916 13362 15916 13362 0 _0519_
rlabel metal1 12420 14450 12420 14450 0 _0520_
rlabel metal1 15502 14042 15502 14042 0 _0521_
rlabel metal1 14306 14280 14306 14280 0 _0522_
rlabel metal1 9614 12954 9614 12954 0 _0523_
rlabel metal1 10672 14450 10672 14450 0 _0524_
rlabel metal1 11730 12716 11730 12716 0 _0525_
rlabel metal1 11500 11730 11500 11730 0 _0526_
rlabel metal1 13524 11866 13524 11866 0 _0527_
rlabel metal1 16146 11866 16146 11866 0 _0528_
rlabel metal1 14490 12818 14490 12818 0 _0529_
rlabel metal2 12282 14144 12282 14144 0 _0530_
rlabel metal2 12466 11968 12466 11968 0 _0531_
rlabel metal1 16882 12716 16882 12716 0 _0532_
rlabel metal1 15962 13906 15962 13906 0 _0533_
rlabel metal2 12742 13396 12742 13396 0 _0534_
rlabel metal1 15778 14450 15778 14450 0 _0535_
rlabel metal1 14214 14892 14214 14892 0 _0536_
rlabel metal1 4554 12818 4554 12818 0 _0537_
rlabel metal1 4094 12954 4094 12954 0 _0538_
rlabel metal1 9154 12172 9154 12172 0 _0539_
rlabel metal2 6946 13396 6946 13396 0 _0540_
rlabel metal1 8096 16626 8096 16626 0 _0541_
rlabel metal1 4784 15130 4784 15130 0 _0542_
rlabel metal1 6256 16626 6256 16626 0 _0543_
rlabel metal1 5980 13362 5980 13362 0 _0544_
rlabel metal1 8464 12818 8464 12818 0 _0545_
rlabel metal1 8142 15674 8142 15674 0 _0546_
rlabel metal1 6670 15130 6670 15130 0 _0547_
rlabel metal1 6624 12954 6624 12954 0 _0548_
rlabel metal1 7636 15130 7636 15130 0 _0549_
rlabel metal1 7958 13430 7958 13430 0 _0550_
rlabel metal1 5566 12750 5566 12750 0 _0551_
rlabel metal1 4002 10982 4002 10982 0 _0552_
rlabel metal1 7958 12274 7958 12274 0 _0553_
rlabel metal1 6716 12274 6716 12274 0 _0554_
rlabel metal1 7314 16626 7314 16626 0 _0555_
rlabel metal1 4830 15980 4830 15980 0 _0556_
rlabel metal1 6578 17068 6578 17068 0 _0557_
rlabel metal1 5842 12954 5842 12954 0 _0558_
rlabel metal1 7452 12818 7452 12818 0 _0559_
rlabel metal1 5382 15130 5382 15130 0 _0560_
rlabel metal1 6118 15130 6118 15130 0 _0561_
rlabel metal1 7728 13362 7728 13362 0 _0562_
rlabel metal1 7314 14858 7314 14858 0 _0563_
rlabel metal1 8510 14892 8510 14892 0 _0564_
rlabel metal2 4186 7174 4186 7174 0 _0565_
rlabel metal1 3864 6970 3864 6970 0 _0566_
rlabel metal1 8832 8398 8832 8398 0 _0567_
rlabel metal1 7084 6834 7084 6834 0 _0568_
rlabel metal1 9936 10642 9936 10642 0 _0569_
rlabel metal1 2576 11322 2576 11322 0 _0570_
rlabel metal1 1748 8602 1748 8602 0 _0571_
rlabel metal1 4968 7922 4968 7922 0 _0572_
rlabel metal1 6394 8466 6394 8466 0 _0573_
rlabel metal1 4370 11186 4370 11186 0 _0574_
rlabel metal1 2944 8262 2944 8262 0 _0575_
rlabel metal1 4462 8602 4462 8602 0 _0576_
rlabel metal1 4600 9554 4600 9554 0 _0577_
rlabel metal1 6578 9656 6578 9656 0 _0578_
rlabel metal1 5244 6970 5244 6970 0 _0579_
rlabel metal1 3082 7276 3082 7276 0 _0580_
rlabel metal1 8832 7922 8832 7922 0 _0581_
rlabel metal2 6026 7174 6026 7174 0 _0582_
rlabel metal1 9246 11220 9246 11220 0 _0583_
rlabel metal1 2162 10540 2162 10540 0 _0584_
rlabel metal1 2300 8942 2300 8942 0 _0585_
rlabel metal1 2599 8602 2599 8602 0 _0586_
rlabel metal1 6256 7514 6256 7514 0 _0587_
rlabel metal1 2944 11186 2944 11186 0 _0588_
rlabel metal1 3036 8466 3036 8466 0 _0589_
rlabel metal2 4922 8772 4922 8772 0 _0590_
rlabel metal1 3910 9656 3910 9656 0 _0591_
rlabel metal1 5704 8874 5704 8874 0 _0592_
rlabel metal1 10028 5338 10028 5338 0 _0593_
rlabel metal1 8878 5746 8878 5746 0 _0594_
rlabel metal1 12788 8398 12788 8398 0 _0595_
rlabel metal1 12742 6732 12742 6732 0 _0596_
rlabel metal2 10994 10948 10994 10948 0 _0597_
rlabel metal1 12006 10676 12006 10676 0 _0598_
rlabel metal1 9292 9010 9292 9010 0 _0599_
rlabel metal2 13110 6052 13110 6052 0 _0600_
rlabel metal1 13340 7922 13340 7922 0 _0601_
rlabel metal1 11776 9690 11776 9690 0 _0602_
rlabel metal2 10902 9044 10902 9044 0 _0603_
rlabel metal2 10994 7378 10994 7378 0 _0604_
rlabel metal1 11684 8602 11684 8602 0 _0605_
rlabel metal2 9890 7208 9890 7208 0 _0606_
rlabel metal1 10166 5100 10166 5100 0 _0607_
rlabel metal1 9246 6358 9246 6358 0 _0608_
rlabel metal1 11914 6970 11914 6970 0 _0609_
rlabel metal1 12650 6426 12650 6426 0 _0610_
rlabel metal1 11822 11220 11822 11220 0 _0611_
rlabel metal1 12788 10574 12788 10574 0 _0612_
rlabel metal1 9246 9690 9246 9690 0 _0613_
rlabel metal1 10442 5882 10442 5882 0 _0614_
rlabel metal1 13294 7276 13294 7276 0 _0615_
rlabel metal2 12558 9860 12558 9860 0 _0616_
rlabel metal1 9706 9452 9706 9452 0 _0617_
rlabel metal1 11730 7276 11730 7276 0 _0618_
rlabel metal1 11132 8602 11132 8602 0 _0619_
rlabel metal2 9706 7582 9706 7582 0 _0620_
rlabel metal1 15180 5746 15180 5746 0 _0621_
rlabel metal1 15778 6188 15778 6188 0 _0622_
rlabel metal1 15916 8398 15916 8398 0 _0623_
rlabel metal1 14674 6970 14674 6970 0 _0624_
rlabel metal1 14490 10642 14490 10642 0 _0625_
rlabel metal1 15916 10098 15916 10098 0 _0626_
rlabel metal1 13524 9146 13524 9146 0 _0627_
rlabel metal1 15778 5100 15778 5100 0 _0628_
rlabel metal1 16468 7922 16468 7922 0 _0629_
rlabel metal1 15226 9146 15226 9146 0 _0630_
rlabel metal1 14628 9010 14628 9010 0 _0631_
rlabel metal2 16238 4454 16238 4454 0 _0632_
rlabel metal1 14030 5270 14030 5270 0 _0633_
rlabel metal1 14122 4658 14122 4658 0 _0634_
rlabel metal1 15042 5236 15042 5236 0 _0635_
rlabel metal1 15916 5746 15916 5746 0 _0636_
rlabel metal1 15410 7820 15410 7820 0 _0637_
rlabel metal1 14766 7378 14766 7378 0 _0638_
rlabel metal1 14260 10778 14260 10778 0 _0639_
rlabel metal2 15870 10812 15870 10812 0 _0640_
rlabel metal1 14214 9486 14214 9486 0 _0641_
rlabel metal1 16422 5338 16422 5338 0 _0642_
rlabel metal1 15870 7276 15870 7276 0 _0643_
rlabel metal1 15778 9146 15778 9146 0 _0644_
rlabel metal1 13340 5882 13340 5882 0 _0645_
rlabel metal1 16330 4556 16330 4556 0 _0646_
rlabel metal2 14122 4080 14122 4080 0 _0647_
rlabel metal1 13478 4216 13478 4216 0 _0648_
rlabel metal1 17848 5746 17848 5746 0 _0649_
rlabel metal1 18998 6290 18998 6290 0 _0650_
rlabel metal1 19458 8398 19458 8398 0 _0651_
rlabel metal1 17250 7378 17250 7378 0 _0652_
rlabel metal1 17434 10234 17434 10234 0 _0653_
rlabel metal1 18308 10098 18308 10098 0 _0654_
rlabel metal1 17756 9146 17756 9146 0 _0655_
rlabel metal2 19366 5117 19366 5117 0 _0656_
rlabel metal1 19090 7514 19090 7514 0 _0657_
rlabel metal1 18538 9146 18538 9146 0 _0658_
rlabel metal1 17848 8398 17848 8398 0 _0659_
rlabel metal2 17986 3332 17986 3332 0 _0660_
rlabel metal1 21390 2312 21390 2312 0 _0661_
rlabel metal1 21022 3162 21022 3162 0 _0662_
rlabel metal1 18630 4794 18630 4794 0 _0663_
rlabel metal1 19458 5780 19458 5780 0 _0664_
rlabel metal2 19734 7684 19734 7684 0 _0665_
rlabel metal1 17756 6970 17756 6970 0 _0666_
rlabel metal1 17480 9894 17480 9894 0 _0667_
rlabel metal1 19389 10030 19389 10030 0 _0668_
rlabel metal1 17204 9146 17204 9146 0 _0669_
rlabel metal1 22034 5032 22034 5032 0 _0670_
rlabel metal1 18676 7378 18676 7378 0 _0671_
rlabel metal1 19228 9146 19228 9146 0 _0672_
rlabel metal1 17572 2618 17572 2618 0 _0673_
rlabel metal1 19596 2618 19596 2618 0 _0674_
rlabel metal1 17986 2822 17986 2822 0 _0675_
rlabel metal1 19044 2958 19044 2958 0 _0676_
rlabel metal1 21666 6834 21666 6834 0 _0677_
rlabel metal1 22770 6834 22770 6834 0 _0678_
rlabel metal1 21022 9010 21022 9010 0 _0679_
rlabel metal1 21804 8058 21804 8058 0 _0680_
rlabel metal1 23644 11118 23644 11118 0 _0681_
rlabel metal1 23874 10098 23874 10098 0 _0682_
rlabel metal1 23138 9554 23138 9554 0 _0683_
rlabel metal1 23966 6902 23966 6902 0 _0684_
rlabel metal1 23092 8602 23092 8602 0 _0685_
rlabel metal1 24380 10778 24380 10778 0 _0686_
rlabel metal1 24242 8602 24242 8602 0 _0687_
rlabel metal1 23736 5746 23736 5746 0 _0688_
rlabel metal1 25208 9146 25208 9146 0 _0689_
rlabel metal1 24288 6698 24288 6698 0 _0690_
rlabel metal2 21022 7004 21022 7004 0 _0691_
rlabel metal1 22034 7276 22034 7276 0 _0692_
rlabel metal1 20516 8602 20516 8602 0 _0693_
rlabel metal2 21022 8738 21022 8738 0 _0694_
rlabel metal1 23368 11322 23368 11322 0 _0695_
rlabel metal1 23460 10574 23460 10574 0 _0696_
rlabel metal1 22678 10132 22678 10132 0 _0697_
rlabel metal1 23966 4726 23966 4726 0 _0698_
rlabel via2 24058 9163 24058 9163 0 _0699_
rlabel metal1 25392 9350 25392 9350 0 _0700_
rlabel metal1 24518 8058 24518 8058 0 _0701_
rlabel metal1 23368 8058 23368 8058 0 _0702_
rlabel metal1 26312 8466 26312 8466 0 _0703_
rlabel metal1 23782 7276 23782 7276 0 _0704_
rlabel metal1 19918 16218 19918 16218 0 _0705_
rlabel metal1 20286 16014 20286 16014 0 _0706_
rlabel metal1 18676 15538 18676 15538 0 _0707_
rlabel metal1 20608 15538 20608 15538 0 _0708_
rlabel metal1 17986 12954 17986 12954 0 _0709_
rlabel metal1 17894 14042 17894 14042 0 _0710_
rlabel metal1 19044 12410 19044 12410 0 _0711_
rlabel metal1 20562 16116 20562 16116 0 _0712_
rlabel metal1 19274 14586 19274 14586 0 _0713_
rlabel metal1 19228 13362 19228 13362 0 _0714_
rlabel metal1 19826 12410 19826 12410 0 _0715_
rlabel metal2 21482 14178 21482 14178 0 _0716_
rlabel metal1 21252 12954 21252 12954 0 _0717_
rlabel metal2 22034 11560 22034 11560 0 _0718_
rlabel metal1 19642 16626 19642 16626 0 _0719_
rlabel metal1 20930 17068 20930 17068 0 _0720_
rlabel metal1 18400 14586 18400 14586 0 _0721_
rlabel metal1 20010 14586 20010 14586 0 _0722_
rlabel metal1 17618 13396 17618 13396 0 _0723_
rlabel metal1 17572 14994 17572 14994 0 _0724_
rlabel metal1 18354 12682 18354 12682 0 _0725_
rlabel metal2 21114 16422 21114 16422 0 _0726_
rlabel metal1 20654 14586 20654 14586 0 _0727_
rlabel metal1 19090 13906 19090 13906 0 _0728_
rlabel metal1 20424 12410 20424 12410 0 _0729_
rlabel metal1 20976 14450 20976 14450 0 _0730_
rlabel metal1 21022 12342 21022 12342 0 _0731_
rlabel metal1 21965 12138 21965 12138 0 _0732_
rlabel metal1 23598 15436 23598 15436 0 _0733_
rlabel metal1 22724 14586 22724 14586 0 _0734_
rlabel metal1 23322 13906 23322 13906 0 _0735_
rlabel metal1 23000 12954 23000 12954 0 _0736_
rlabel metal1 26450 15606 26450 15606 0 _0737_
rlabel metal1 25668 15538 25668 15538 0 _0738_
rlabel metal1 27692 14314 27692 14314 0 _0739_
rlabel metal1 24748 14586 24748 14586 0 _0740_
rlabel metal1 24380 13362 24380 13362 0 _0741_
rlabel metal1 28428 14042 28428 14042 0 _0742_
rlabel metal1 27370 13906 27370 13906 0 _0743_
rlabel metal1 25668 13362 25668 13362 0 _0744_
rlabel metal1 27922 12852 27922 12852 0 _0745_
rlabel metal1 26266 12274 26266 12274 0 _0746_
rlabel metal1 23552 16082 23552 16082 0 _0747_
rlabel metal2 22034 14756 22034 14756 0 _0748_
rlabel metal1 23598 12818 23598 12818 0 _0749_
rlabel metal1 22448 12954 22448 12954 0 _0750_
rlabel metal2 27462 15334 27462 15334 0 _0751_
rlabel metal2 24886 15810 24886 15810 0 _0752_
rlabel metal1 28106 13804 28106 13804 0 _0753_
rlabel metal1 25438 14926 25438 14926 0 _0754_
rlabel metal1 24150 12716 24150 12716 0 _0755_
rlabel metal1 26680 14926 26680 14926 0 _0756_
rlabel metal1 27922 12308 27922 12308 0 _0757_
rlabel metal2 24610 13855 24610 13855 0 _0758_
rlabel metal1 27324 10778 27324 10778 0 _0759_
rlabel metal1 27416 13226 27416 13226 0 _0760_
rlabel metal1 23920 17850 23920 17850 0 _0761_
rlabel metal1 22908 17306 22908 17306 0 _0762_
rlabel metal1 25254 18394 25254 18394 0 _0763_
rlabel metal1 24748 18394 24748 18394 0 _0764_
rlabel metal1 27324 20434 27324 20434 0 _0765_
rlabel metal1 25714 20026 25714 20026 0 _0766_
rlabel metal1 27140 19346 27140 19346 0 _0767_
rlabel metal1 25438 17714 25438 17714 0 _0768_
rlabel metal1 26312 18802 26312 18802 0 _0769_
rlabel metal1 27416 20978 27416 20978 0 _0770_
rlabel metal1 27830 18802 27830 18802 0 _0771_
rlabel metal1 26680 16762 26680 16762 0 _0772_
rlabel metal1 27370 17170 27370 17170 0 _0773_
rlabel metal2 27830 15980 27830 15980 0 _0774_
rlabel metal1 23552 17170 23552 17170 0 _0775_
rlabel metal1 22402 17748 22402 17748 0 _0776_
rlabel metal1 24334 18394 24334 18394 0 _0777_
rlabel metal1 23874 18394 23874 18394 0 _0778_
rlabel metal1 27784 20434 27784 20434 0 _0779_
rlabel metal1 24978 20434 24978 20434 0 _0780_
rlabel metal2 28106 20570 28106 20570 0 _0781_
rlabel metal1 24564 16082 24564 16082 0 _0782_
rlabel metal1 25576 19346 25576 19346 0 _0783_
rlabel metal1 26266 19890 26266 19890 0 _0784_
rlabel metal1 28152 15130 28152 15130 0 _0785_
rlabel metal1 26818 18836 26818 18836 0 _0786_
rlabel metal1 28152 17170 28152 17170 0 _0787_
rlabel metal1 26450 16218 26450 16218 0 _0788_
rlabel metal2 22862 19856 22862 19856 0 _0789_
rlabel metal2 21482 20536 21482 20536 0 _0790_
rlabel metal1 14536 23154 14536 23154 0 _0791_
rlabel metal1 14214 23630 14214 23630 0 _0792_
rlabel metal2 15318 25228 15318 25228 0 _0793_
rlabel metal1 15686 25874 15686 25874 0 _0794_
rlabel metal1 16606 26452 16606 26452 0 _0795_
rlabel metal1 17480 24650 17480 24650 0 _0796_
rlabel metal1 17015 24174 17015 24174 0 _0797_
rlabel metal1 17802 21658 17802 21658 0 _0798_
rlabel metal1 15318 22508 15318 22508 0 _0799_
rlabel metal1 15594 25364 15594 25364 0 _0800_
rlabel metal1 17710 25466 17710 25466 0 _0801_
rlabel metal1 18400 23290 18400 23290 0 _0802_
rlabel metal1 17986 24276 17986 24276 0 _0803_
rlabel metal1 19458 25364 19458 25364 0 _0804_
rlabel metal1 19044 23766 19044 23766 0 _0805_
rlabel metal1 14628 22066 14628 22066 0 _0806_
rlabel metal1 15870 22746 15870 22746 0 _0807_
rlabel metal1 14720 24718 14720 24718 0 _0808_
rlabel metal1 15272 25874 15272 25874 0 _0809_
rlabel metal2 17066 25908 17066 25908 0 _0810_
rlabel metal1 19090 26418 19090 26418 0 _0811_
rlabel metal1 17250 23154 17250 23154 0 _0812_
rlabel metal1 19688 21998 19688 21998 0 _0813_
rlabel metal1 15778 23834 15778 23834 0 _0814_
rlabel metal1 16836 25330 16836 25330 0 _0815_
rlabel metal2 18722 25636 18722 25636 0 _0816_
rlabel metal1 18814 22678 18814 22678 0 _0817_
rlabel metal1 18216 24718 18216 24718 0 _0818_
rlabel metal1 19550 23018 19550 23018 0 _0819_
rlabel metal2 20010 23630 20010 23630 0 _0820_
rlabel metal1 6624 18802 6624 18802 0 _0821_
rlabel metal1 7820 19414 7820 19414 0 _0822_
rlabel metal1 7498 18666 7498 18666 0 _0823_
rlabel metal1 9200 20230 9200 20230 0 _0824_
rlabel metal1 2024 13362 2024 13362 0 _0825_
rlabel metal2 3082 14892 3082 14892 0 _0826_
rlabel metal1 3956 15946 3956 15946 0 _0827_
rlabel metal1 3082 17850 3082 17850 0 _0828_
rlabel metal1 3128 19822 3128 19822 0 _0829_
rlabel metal1 2346 22406 2346 22406 0 _0830_
rlabel metal2 2806 24990 2806 24990 0 _0831_
rlabel metal1 2990 23154 2990 23154 0 _0832_
rlabel metal1 4002 14484 4002 14484 0 _0833_
rlabel metal1 4370 17748 4370 17748 0 _0834_
rlabel metal1 3956 19482 3956 19482 0 _0835_
rlabel metal1 4462 21114 4462 21114 0 _0836_
rlabel metal1 5014 18836 5014 18836 0 _0837_
rlabel metal1 4876 19346 4876 19346 0 _0838_
rlabel metal1 6578 19448 6578 19448 0 _0839_
rlabel metal1 3404 13838 3404 13838 0 _0840_
rlabel metal1 3588 14994 3588 14994 0 _0841_
rlabel metal1 3266 17170 3266 17170 0 _0842_
rlabel metal1 3910 18394 3910 18394 0 _0843_
rlabel metal1 3634 19278 3634 19278 0 _0844_
rlabel metal1 2622 22576 2622 22576 0 _0845_
rlabel metal1 3634 24242 3634 24242 0 _0846_
rlabel metal1 4002 22508 4002 22508 0 _0847_
rlabel metal1 4232 14926 4232 14926 0 _0848_
rlabel metal1 4508 18190 4508 18190 0 _0849_
rlabel metal1 3634 20978 3634 20978 0 _0850_
rlabel metal1 3726 21114 3726 21114 0 _0851_
rlabel metal1 5428 18394 5428 18394 0 _0852_
rlabel metal1 5106 20332 5106 20332 0 _0853_
rlabel metal1 5014 19720 5014 19720 0 _0854_
rlabel metal1 7682 9996 7682 9996 0 _0855_
rlabel metal1 8188 10234 8188 10234 0 _0856_
rlabel metal1 7452 9622 7452 9622 0 _0857_
rlabel metal2 2070 11560 2070 11560 0 _0858_
rlabel metal1 11408 3434 11408 3434 0 _0859_
rlabel metal1 9568 3570 9568 3570 0 _0860_
rlabel metal1 8142 3604 8142 3604 0 _0861_
rlabel metal1 6394 3706 6394 3706 0 _0862_
rlabel metal1 4922 2380 4922 2380 0 _0863_
rlabel metal1 4830 4658 4830 4658 0 _0864_
rlabel metal2 3082 5372 3082 5372 0 _0865_
rlabel metal1 4922 5338 4922 5338 0 _0866_
rlabel metal2 12558 4522 12558 4522 0 _0867_
rlabel metal1 8372 4114 8372 4114 0 _0868_
rlabel metal1 6578 4012 6578 4012 0 _0869_
rlabel metal1 6394 5338 6394 5338 0 _0870_
rlabel metal1 9522 4658 9522 4658 0 _0871_
rlabel metal1 7728 5066 7728 5066 0 _0872_
rlabel metal1 7774 8602 7774 8602 0 _0873_
rlabel metal1 10948 2618 10948 2618 0 _0874_
rlabel metal1 10258 4046 10258 4046 0 _0875_
rlabel metal2 6624 3434 6624 3434 0 _0876_
rlabel metal1 6578 2516 6578 2516 0 _0877_
rlabel metal1 2622 2856 2622 2856 0 _0878_
rlabel metal1 4784 4114 4784 4114 0 _0879_
rlabel metal2 3174 4420 3174 4420 0 _0880_
rlabel metal1 5842 5814 5842 5814 0 _0881_
rlabel metal1 10626 4658 10626 4658 0 _0882_
rlabel metal1 7590 4522 7590 4522 0 _0883_
rlabel metal1 6072 4658 6072 4658 0 _0884_
rlabel metal1 6946 4794 6946 4794 0 _0885_
rlabel metal1 8372 4658 8372 4658 0 _0886_
rlabel metal2 7498 5508 7498 5508 0 _0887_
rlabel metal1 7222 8534 7222 8534 0 _0888_
rlabel metal2 20470 5474 20470 5474 0 _0889_
rlabel metal1 22770 5644 22770 5644 0 _0890_
rlabel metal2 21390 6290 21390 6290 0 _0891_
rlabel metal1 19550 1938 19550 1938 0 _0892_
rlabel metal1 28106 9690 28106 9690 0 _0893_
rlabel metal1 26404 10030 26404 10030 0 _0894_
rlabel metal2 24794 4726 24794 4726 0 _0895_
rlabel metal3 19780 8092 19780 8092 0 _0896_
rlabel metal2 19642 7973 19642 7973 0 _0897_
rlabel metal2 23506 9486 23506 9486 0 _0898_
rlabel metal1 2070 2040 2070 2040 0 _0899_
rlabel metal1 22632 4590 22632 4590 0 _0900_
rlabel metal2 28014 8908 28014 8908 0 _0901_
rlabel metal2 21574 7072 21574 7072 0 _0902_
rlabel metal2 19182 4862 19182 4862 0 _0903_
rlabel metal1 21206 11560 21206 11560 0 _0904_
rlabel metal1 27140 8398 27140 8398 0 _0905_
rlabel metal1 17572 3366 17572 3366 0 _0906_
rlabel metal2 26634 5066 26634 5066 0 _0907_
rlabel metal2 2530 3417 2530 3417 0 bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal2 13662 2142 13662 2142 0 bottom_width_0_height_0_subtile_0__pin_I_6_
rlabel metal2 21022 2516 21022 2516 0 bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 26726 23120 26726 23120 0 ccff_head
rlabel metal2 28474 27149 28474 27149 0 ccff_tail
rlabel metal3 1050 9588 1050 9588 0 clk
rlabel metal1 18722 8534 18722 8534 0 clknet_0_prog_clk
rlabel metal1 2208 2482 2208 2482 0 clknet_4_0_0_prog_clk
rlabel metal1 21850 3978 21850 3978 0 clknet_4_10_0_prog_clk
rlabel metal1 20838 11152 20838 11152 0 clknet_4_11_0_prog_clk
rlabel metal1 19688 17646 19688 17646 0 clknet_4_12_0_prog_clk
rlabel metal1 19550 20910 19550 20910 0 clknet_4_13_0_prog_clk
rlabel metal1 24012 19346 24012 19346 0 clknet_4_14_0_prog_clk
rlabel metal1 21252 24786 21252 24786 0 clknet_4_15_0_prog_clk
rlabel metal1 1518 12750 1518 12750 0 clknet_4_1_0_prog_clk
rlabel metal1 11500 2482 11500 2482 0 clknet_4_2_0_prog_clk
rlabel metal1 13294 13940 13294 13940 0 clknet_4_3_0_prog_clk
rlabel metal2 1426 19584 1426 19584 0 clknet_4_4_0_prog_clk
rlabel metal1 2254 23732 2254 23732 0 clknet_4_5_0_prog_clk
rlabel metal2 12742 20060 12742 20060 0 clknet_4_6_0_prog_clk
rlabel metal1 8878 20944 8878 20944 0 clknet_4_7_0_prog_clk
rlabel metal1 16974 6324 16974 6324 0 clknet_4_8_0_prog_clk
rlabel metal2 16698 2621 16698 2621 0 clknet_4_9_0_prog_clk
rlabel metal1 2714 24616 2714 24616 0 left_width_0_height_0_subtile_0__pin_I_3_
rlabel metal3 1142 23732 1142 23732 0 left_width_0_height_0_subtile_0__pin_I_7_
rlabel metal3 820 27268 820 27268 0 left_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 23272 3502 23272 3502 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
rlabel metal2 22034 6817 22034 6817 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
rlabel metal2 23552 2550 23552 2550 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
rlabel metal1 16974 6732 16974 6732 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
rlabel metal1 21390 9554 21390 9554 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
rlabel metal1 16652 8942 16652 8942 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
rlabel metal2 24242 7038 24242 7038 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
rlabel metal1 28336 16626 28336 16626 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
rlabel metal1 24748 6630 24748 6630 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
rlabel metal2 27094 3519 27094 3519 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
rlabel metal2 22126 10336 22126 10336 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
rlabel metal3 21436 3332 21436 3332 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
rlabel metal3 21252 3468 21252 3468 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
rlabel metal3 17204 7548 17204 7548 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
rlabel metal2 15778 3604 15778 3604 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
rlabel metal1 14398 2584 14398 2584 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
rlabel via2 4370 2907 4370 2907 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
rlabel metal1 23506 4046 23506 4046 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
rlabel metal2 23782 3910 23782 3910 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
rlabel metal1 24472 2278 24472 2278 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
rlabel metal1 23138 6732 23138 6732 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
rlabel via2 27554 10557 27554 10557 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
rlabel metal1 27278 9554 27278 9554 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
rlabel metal1 26818 11254 26818 11254 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
rlabel metal1 26358 10132 26358 10132 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
rlabel metal1 26910 10098 26910 10098 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
rlabel metal1 27048 9010 27048 9010 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
rlabel metal1 20746 11288 20746 11288 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
rlabel via2 19458 11203 19458 11203 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
rlabel metal2 26174 7548 26174 7548 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
rlabel metal1 26542 5882 26542 5882 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
rlabel metal2 17434 7905 17434 7905 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
rlabel metal1 26680 6970 26680 6970 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
rlabel metal1 28198 5882 28198 5882 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
rlabel metal1 27784 4658 27784 4658 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
rlabel metal2 28566 5559 28566 5559 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
rlabel metal4 20700 6664 20700 6664 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
rlabel metal2 15870 6137 15870 6137 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
rlabel metal2 16330 5100 16330 5100 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
rlabel metal1 28290 9622 28290 9622 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
rlabel metal2 25806 4930 25806 4930 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
rlabel metal1 25024 5338 25024 5338 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
rlabel metal1 26588 6902 26588 6902 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
rlabel metal1 25346 5882 25346 5882 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
rlabel metal2 27646 9520 27646 9520 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
rlabel metal1 27416 7990 27416 7990 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
rlabel metal1 27784 6222 27784 6222 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
rlabel metal1 26634 4522 26634 4522 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
rlabel metal1 26312 3978 26312 3978 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
rlabel metal1 24564 4250 24564 4250 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
rlabel metal1 23460 4726 23460 4726 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
rlabel metal1 28428 8602 28428 8602 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
rlabel metal1 27876 6766 27876 6766 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
rlabel metal1 22452 5202 22452 5202 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
rlabel metal1 20102 5746 20102 5746 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
rlabel metal2 20930 6358 20930 6358 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 19090 14926 19090 14926 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2530 12308 2530 12308 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
rlabel metal1 8372 9146 8372 9146 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
rlabel metal1 6394 6324 6394 6324 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
rlabel metal1 19182 4080 19182 4080 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
rlabel metal2 13846 3876 13846 3876 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
rlabel metal1 10764 7446 10764 7446 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
rlabel metal1 6992 9418 6992 9418 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
rlabel metal2 16790 3825 16790 3825 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
rlabel metal1 11638 3162 11638 3162 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
rlabel metal1 4094 4114 4094 4114 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
rlabel metal1 5014 4250 5014 4250 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
rlabel metal1 2024 3502 2024 3502 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
rlabel metal1 4370 3672 4370 3672 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
rlabel metal1 2369 6222 2369 6222 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
rlabel metal2 2898 5916 2898 5916 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
rlabel metal2 3450 6324 3450 6324 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
rlabel metal1 3680 5202 3680 5202 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
rlabel metal2 4186 5882 4186 5882 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
rlabel metal1 4830 5678 4830 5678 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
rlabel metal1 6072 5678 6072 5678 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
rlabel metal1 7636 9010 7636 9010 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
rlabel metal2 13202 2346 13202 2346 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
rlabel metal1 9614 2618 9614 2618 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
rlabel metal1 13616 2550 13616 2550 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
rlabel metal1 9154 3502 9154 3502 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
rlabel metal1 10534 2618 10534 2618 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
rlabel metal1 10212 4114 10212 4114 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
rlabel metal1 7314 2958 7314 2958 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
rlabel metal1 7452 3570 7452 3570 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
rlabel metal1 7314 3026 7314 3026 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
rlabel metal2 6486 3536 6486 3536 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
rlabel metal1 7038 3502 7038 3502 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
rlabel metal1 5106 3570 5106 3570 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
rlabel metal1 4140 2482 4140 2482 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
rlabel metal1 6118 2482 6118 2482 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
rlabel metal1 2070 3060 2070 3060 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
rlabel metal1 2208 2822 2208 2822 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
rlabel metal1 2070 3570 2070 3570 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
rlabel metal1 3772 3502 3772 3502 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
rlabel metal2 12466 4420 12466 4420 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
rlabel metal1 7222 4726 7222 4726 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
rlabel metal1 7176 5542 7176 5542 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
rlabel metal2 8510 6936 8510 6936 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
rlabel metal1 7636 5882 7636 5882 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
rlabel metal1 10258 3910 10258 3910 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
rlabel metal1 8970 3706 8970 3706 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
rlabel metal1 7268 3978 7268 3978 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
rlabel metal1 4968 3706 4968 3706 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
rlabel metal2 4830 4216 4830 4216 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
rlabel metal1 4784 4998 4784 4998 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
rlabel metal1 5934 5542 5934 5542 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
rlabel metal2 12834 4896 12834 4896 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
rlabel metal1 8096 4590 8096 4590 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
rlabel metal1 6762 8942 6762 8942 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
rlabel metal1 7544 10030 7544 10030 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
rlabel metal2 7866 10404 7866 10404 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 12558 11152 12558 11152 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7866 21556 7866 21556 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
rlabel metal1 6440 18258 6440 18258 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
rlabel metal1 5106 23290 5106 23290 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
rlabel metal1 2346 22644 2346 22644 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
rlabel metal1 4554 14994 4554 14994 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
rlabel metal2 11362 19584 11362 19584 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
rlabel metal1 6026 20400 6026 20400 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
rlabel metal1 1702 14450 1702 14450 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
rlabel metal2 2070 13770 2070 13770 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
rlabel metal2 1702 23392 1702 23392 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
rlabel metal1 2346 21454 2346 21454 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
rlabel metal2 2714 22372 2714 22372 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
rlabel metal1 2599 21386 2599 21386 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
rlabel metal2 2622 24276 2622 24276 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
rlabel metal2 3082 24990 3082 24990 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
rlabel metal1 2852 24378 2852 24378 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
rlabel metal1 3404 24174 3404 24174 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
rlabel metal1 3726 23834 3726 23834 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
rlabel metal1 3220 23086 3220 23086 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
rlabel metal1 4094 22610 4094 22610 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
rlabel metal1 6670 19210 6670 19210 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
rlabel metal1 3358 13294 3358 13294 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
rlabel metal1 3404 13498 3404 13498 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
rlabel metal1 1978 14348 1978 14348 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
rlabel metal1 2300 14450 2300 14450 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
rlabel metal2 2254 15300 2254 15300 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
rlabel metal2 2898 14756 2898 14756 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
rlabel metal1 3588 16626 3588 16626 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
rlabel metal1 4508 16762 4508 16762 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
rlabel metal1 2990 16762 2990 16762 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
rlabel metal2 3266 16932 3266 16932 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
rlabel metal1 2576 18734 2576 18734 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
rlabel metal1 2530 18326 2530 18326 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
rlabel metal1 3450 18768 3450 18768 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
rlabel metal1 3680 18734 3680 18734 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
rlabel metal1 2231 20434 2231 20434 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
rlabel metal1 2277 20298 2277 20298 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
rlabel metal2 2070 20196 2070 20196 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
rlabel metal1 1518 19448 1518 19448 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
rlabel metal2 3266 13532 3266 13532 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
rlabel metal2 4278 20400 4278 20400 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
rlabel metal1 4738 21658 4738 21658 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
rlabel metal1 6348 18938 6348 18938 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
rlabel metal2 4922 19992 4922 19992 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
rlabel metal1 3220 14790 3220 14790 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
rlabel metal1 4140 17034 4140 17034 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
rlabel metal1 4232 18258 4232 18258 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
rlabel metal1 3588 19686 3588 19686 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
rlabel metal1 3496 21318 3496 21318 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
rlabel metal1 3864 22066 3864 22066 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
rlabel metal1 4324 22746 4324 22746 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
rlabel metal1 4646 14790 4646 14790 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
rlabel metal1 4922 18326 4922 18326 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
rlabel metal2 6486 21250 6486 21250 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
rlabel metal1 7958 18394 7958 18394 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
rlabel metal1 7360 18802 7360 18802 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9614 19278 9614 19278 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 21758 18258 21758 18258 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
rlabel metal1 18170 18258 18170 18258 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in
rlabel metal1 19780 21522 19780 21522 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail
rlabel metal1 12466 24820 12466 24820 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out
rlabel metal1 18584 23086 18584 23086 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out
rlabel metal1 19596 24174 19596 24174 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out
rlabel metal1 19734 24718 19734 24718 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out
rlabel metal1 13248 20978 13248 20978 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in
rlabel metal1 14076 21658 14076 21658 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out
rlabel metal1 18814 27438 18814 27438 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in
rlabel metal1 17940 26350 17940 26350 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out
rlabel metal1 19654 27438 19654 27438 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in
rlabel metal1 19458 26350 19458 26350 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out
rlabel metal2 17894 25585 17894 25585 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in
rlabel metal1 16974 24310 16974 24310 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out
rlabel metal1 17158 22678 17158 22678 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in
rlabel metal1 17572 22746 17572 22746 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out
rlabel metal1 18538 21998 18538 21998 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in
rlabel metal1 18584 22202 18584 22202 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out
rlabel metal1 19688 22066 19688 22066 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out
rlabel metal1 20010 23630 20010 23630 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in
rlabel metal1 13800 22066 13800 22066 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in
rlabel metal1 13984 21998 13984 21998 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out
rlabel metal1 14076 24174 14076 24174 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in
rlabel metal1 14260 23698 14260 23698 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out
rlabel metal1 14076 23834 14076 23834 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in
rlabel metal1 14490 22746 14490 22746 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out
rlabel metal1 14214 26282 14214 26282 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in
rlabel metal1 15042 24718 15042 24718 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out
rlabel metal2 13938 25602 13938 25602 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in
rlabel metal1 14398 24684 14398 24684 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out
rlabel metal1 13570 27438 13570 27438 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in
rlabel metal1 13294 27540 13294 27540 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out
rlabel metal1 14628 27438 14628 27438 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in
rlabel metal1 14904 25806 14904 25806 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out
rlabel metal1 16652 27438 16652 27438 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in
rlabel metal1 16468 26418 16468 26418 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out
rlabel metal1 17342 27506 17342 27506 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in
rlabel metal1 17434 26418 17434 26418 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out
rlabel metal1 15180 22542 15180 22542 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out
rlabel metal1 18584 25670 18584 25670 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out
rlabel metal2 19366 23290 19366 23290 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out
rlabel metal2 18262 24480 18262 24480 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out
rlabel metal1 19780 23698 19780 23698 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out
rlabel metal2 14766 24072 14766 24072 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out
rlabel metal1 15272 24582 15272 24582 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out
rlabel metal1 15916 25670 15916 25670 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out
rlabel metal1 17296 26486 17296 26486 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out
rlabel metal1 19228 26282 19228 26282 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out
rlabel metal1 17756 23698 17756 23698 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out
rlabel metal1 19228 22406 19228 22406 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out
rlabel metal1 15824 24038 15824 24038 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out
rlabel metal1 16422 25126 16422 25126 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out
rlabel metal1 21068 19346 21068 19346 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q
rlabel metal1 20378 18156 20378 18156 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out
rlabel metal1 22264 20366 22264 20366 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out
rlabel via1 20930 19958 20930 19958 0 logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 21942 17646 21942 17646 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q
rlabel metal1 28244 20910 28244 20910 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q
rlabel metal1 27692 19890 27692 19890 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q
rlabel metal1 25760 16966 25760 16966 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q
rlabel metal1 22586 13906 22586 13906 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q
rlabel metal2 27094 13583 27094 13583 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q
rlabel metal1 27002 12682 27002 12682 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q
rlabel metal1 26864 12818 26864 12818 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q
rlabel metal1 18492 16082 18492 16082 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q
rlabel metal1 20378 14348 20378 14348 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q
rlabel metal1 21758 12818 21758 12818 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q
rlabel metal1 21758 11118 21758 11118 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q
rlabel metal1 20056 10030 20056 10030 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q
rlabel metal1 21528 10438 21528 10438 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q
rlabel metal1 24518 8466 24518 8466 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q
rlabel metal1 24058 5338 24058 5338 0 logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q
rlabel metal2 19366 6596 19366 6596 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q
rlabel metal1 19642 4080 19642 4080 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q
rlabel metal1 18446 2346 18446 2346 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q
rlabel metal1 15962 2380 15962 2380 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q
rlabel metal1 15180 2414 15180 2414 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q
rlabel metal1 16882 5168 16882 5168 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q
rlabel metal1 13202 3468 13202 3468 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q
rlabel metal1 12926 4658 12926 4658 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q
rlabel metal1 9200 5202 9200 5202 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q
rlabel metal1 12834 9588 12834 9588 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q
rlabel metal1 10580 7718 10580 7718 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q
rlabel metal1 9614 7310 9614 7310 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q
rlabel metal1 2070 7378 2070 7378 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q
rlabel metal1 2576 10030 2576 10030 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q
rlabel metal1 4646 8432 4646 8432 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q
rlabel metal1 6256 10642 6256 10642 0 logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q
rlabel metal1 3726 11730 3726 11730 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q
rlabel via2 8050 13923 8050 13923 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q
rlabel metal1 7452 13838 7452 13838 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q
rlabel metal1 8464 14246 8464 14246 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q
rlabel metal1 10948 12818 10948 12818 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q
rlabel metal2 11086 12546 11086 12546 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q
rlabel metal1 14490 14042 14490 14042 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q
rlabel metal2 13478 14654 13478 14654 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q
rlabel metal1 13938 15538 13938 15538 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q
rlabel metal2 8970 20944 8970 20944 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q
rlabel metal1 10672 18258 10672 18258 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q
rlabel metal1 9614 19414 9614 19414 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q
rlabel metal1 6808 21522 6808 21522 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q
rlabel metal1 8188 26350 8188 26350 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q
rlabel metal1 5336 24582 5336 24582 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q
rlabel metal1 6854 25806 6854 25806 0 logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q
rlabel metal1 8648 21998 8648 21998 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q
rlabel metal2 10442 24106 10442 24106 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q
rlabel metal1 11730 25160 11730 25160 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q
rlabel metal1 11500 24786 11500 24786 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q
rlabel metal1 14260 18258 14260 18258 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q
rlabel metal1 15870 17612 15870 17612 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q
rlabel metal1 17434 18836 17434 18836 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q
rlabel metal2 18906 19074 18906 19074 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q
rlabel metal1 20884 20910 20884 20910 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q
rlabel metal1 23644 27438 23644 27438 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q
rlabel metal2 23138 23596 23138 23596 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q
rlabel metal1 24702 24684 24702 24684 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q
rlabel metal1 25070 21522 25070 21522 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q
rlabel metal1 27002 24820 27002 24820 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q
rlabel metal1 27232 23086 27232 23086 0 logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q
rlabel metal1 20378 21896 20378 21896 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out
rlabel metal1 20562 7752 20562 7752 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out
rlabel metal1 13754 6120 13754 6120 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out
rlabel metal1 2714 24242 2714 24242 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out
rlabel metal1 19734 24174 19734 24174 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out
rlabel metal2 20102 8993 20102 8993 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out
rlabel metal1 13524 6766 13524 6766 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out
rlabel metal2 1978 25041 1978 25041 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out
rlabel metal1 19274 26860 19274 26860 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out
rlabel metal1 20838 14008 20838 14008 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out
rlabel metal2 23874 17680 23874 17680 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 23092 17782 23092 17782 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 25208 18938 25208 18938 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 25070 19074 25070 19074 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 27692 20570 27692 20570 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 25760 20230 25760 20230 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 28014 19346 28014 19346 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out
rlabel metal2 25070 16864 25070 16864 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 26358 19040 26358 19040 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 26818 19958 26818 19958 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 28244 18394 28244 18394 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 26542 17782 26542 17782 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 27048 17306 27048 17306 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 24058 15776 24058 15776 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 23000 14790 23000 14790 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 23690 13192 23690 13192 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 23184 13430 23184 13430 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 27508 15674 27508 15674 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out
rlabel metal2 25806 15776 25806 15776 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 27738 14518 27738 14518 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 25116 14790 25116 14790 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 24610 13498 24610 13498 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 27692 15334 27692 15334 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 27784 11730 27784 11730 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 25300 13498 25300 13498 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 28244 12954 28244 12954 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out
rlabel via1 20378 16422 20378 16422 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 21206 16422 21206 16422 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 18538 15062 18538 15062 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 20700 15130 20700 15130 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 18308 13430 18308 13430 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out
rlabel metal2 17986 14688 17986 14688 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 19228 12682 19228 12682 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 21114 15674 21114 15674 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 20332 14790 20332 14790 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 19642 13600 19642 13600 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 20700 12614 20700 12614 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 21804 11798 21804 11798 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 21574 12274 21574 12274 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 22310 7106 22310 7106 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 22356 7514 22356 7514 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 21252 9078 21252 9078 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 22172 9146 22172 9146 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out
rlabel metal2 24150 11424 24150 11424 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 24242 10574 24242 10574 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 23184 9418 23184 9418 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 23000 7514 23000 7514 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 23230 9146 23230 9146 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 25116 10710 25116 10710 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out
rlabel metal2 25070 8670 25070 8670 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 23598 7582 23598 7582 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 26312 8262 26312 8262 0 logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 18538 5338 18538 5338 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 19458 5882 19458 5882 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 19090 8160 19090 8160 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 18124 7242 18124 7242 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 17940 10778 17940 10778 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 19366 10166 19366 10166 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 18032 9350 18032 9350 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 18170 4454 18170 4454 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 19458 7242 19458 7242 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 20194 2482 20194 2482 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out
rlabel via1 18446 4539 18446 4539 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 19274 3434 19274 3434 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 18078 3094 18078 3094 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 15502 5440 15502 5440 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 16238 5984 16238 5984 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 15870 8160 15870 8160 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 15272 7514 15272 7514 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 14904 10778 14904 10778 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out
rlabel metal2 16054 10336 16054 10336 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 13892 9350 13892 9350 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 16422 5270 16422 5270 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 16146 5916 16146 5916 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 15502 7565 15502 7565 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 14030 6426 14030 6426 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 16330 4454 16330 4454 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 14122 4726 14122 4726 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 10672 5542 10672 5542 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 9614 5984 9614 5984 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 12742 8160 12742 8160 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 13064 7310 13064 7310 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 11776 11322 11776 11322 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out
rlabel metal2 12374 10268 12374 10268 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 10166 9486 10166 9486 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 10672 6154 10672 6154 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13432 7446 13432 7446 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 12052 9894 12052 9894 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 10396 9350 10396 9350 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 11178 7072 11178 7072 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 11040 8806 11040 8806 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 4876 7514 4876 7514 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3772 7242 3772 7242 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 7590 8330 7590 8330 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 6486 7990 6486 7990 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 8786 11322 8786 11322 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 3220 11118 3220 11118 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 2898 9486 2898 9486 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 4416 8534 4416 8534 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6486 7854 6486 7854 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 4186 11254 4186 11254 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 3588 9418 3588 9418 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 5382 9316 5382 9316 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 4646 9418 4646 9418 0 logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 5428 12614 5428 12614 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 4830 13600 4830 13600 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 8464 12682 8464 12682 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 7452 12750 7452 12750 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 8326 16422 8326 16422 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out
rlabel metal2 5198 15776 5198 15776 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 6670 16490 6670 16490 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 5888 13498 5888 13498 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7866 12954 7866 12954 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 7682 15368 7682 15368 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 6716 15674 6716 15674 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 7544 13498 7544 13498 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 7728 15538 7728 15538 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 11132 13158 11132 13158 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 10994 14246 10994 14246 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 12236 13158 12236 13158 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 12282 12070 12282 12070 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 14674 12172 14674 12172 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 16284 12342 16284 12342 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 15364 13294 15364 13294 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out
rlabel via1 12190 14382 12190 14382 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 12650 13498 12650 13498 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 17066 12954 17066 12954 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 16100 14042 16100 14042 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 13064 14042 13064 14042 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 15318 14586 15318 14586 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 9292 18190 9292 18190 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 8786 18734 8786 18734 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 8924 17034 8924 17034 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 9798 16218 9798 16218 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 11638 17102 11638 17102 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 12742 16218 12742 16218 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out
rlabel metal2 12466 19142 12466 19142 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 10028 19958 10028 19958 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10028 17306 10028 17306 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 12604 17306 12604 17306 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out
rlabel metal2 13018 19652 13018 19652 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 10304 18938 10304 18938 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 12282 19686 12282 19686 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 5704 22746 5704 22746 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5750 21998 5750 21998 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 8694 23392 8694 23392 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 7590 22746 7590 22746 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 7314 26826 7314 26826 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 3588 25738 3588 25738 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 3450 26826 3450 26826 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out
rlabel metal2 6118 24208 6118 24208 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7590 23494 7590 23494 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 6394 26452 6394 26452 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 5014 26826 5014 26826 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out
rlabel metal2 6578 24548 6578 24548 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 6210 26588 6210 26588 0 logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 10304 22066 10304 22066 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 11178 21386 11178 21386 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 10258 23766 10258 23766 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 9798 22508 9798 22508 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out
rlabel metal2 9430 26656 9430 26656 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 9200 25738 9200 25738 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 10810 27098 10810 27098 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 11546 23630 11546 23630 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 10994 22780 10994 22780 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 10442 26112 10442 26112 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 12742 26962 12742 26962 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 12052 23154 12052 23154 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 12328 26486 12328 26486 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 16836 15878 16836 15878 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 16238 16864 16238 16864 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 16100 18394 16100 18394 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 14996 17782 14996 17782 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 15226 20332 15226 20332 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 15502 19346 15502 19346 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out
rlabel metal2 16146 21216 16146 21216 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out
rlabel metal2 17250 17170 17250 17170 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 16836 17782 16836 17782 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 15870 20094 15870 20094 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 17158 20910 17158 20910 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 18124 17782 18124 17782 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 18032 20434 18032 20434 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out
rlabel metal1 21160 21318 21160 21318 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 22310 21556 22310 21556 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 21666 23698 21666 23698 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 21068 22202 21068 22202 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out
rlabel metal2 21298 26928 21298 26928 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 21528 25806 21528 25806 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 23368 26826 23368 26826 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out
rlabel via1 22678 21862 22678 21862 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 22218 23392 22218 23392 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 22402 26010 22402 26010 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out
rlabel metal2 24334 26282 24334 26282 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 23920 23494 23920 23494 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 23828 25670 23828 25670 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 24978 21862 24978 21862 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 23966 21114 23966 21114 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 25300 22134 25300 22134 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 25576 22202 25576 22202 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out
rlabel metal1 26128 26010 26128 26010 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out
rlabel metal1 26404 25126 26404 25126 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out
rlabel metal1 27094 26758 27094 26758 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out
rlabel metal1 26404 21862 26404 21862 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 27646 21930 27646 21930 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 27324 25466 27324 25466 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out
rlabel metal1 27646 26282 27646 26282 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out
rlabel metal1 27876 22746 27876 22746 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 28014 25534 28014 25534 0 logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out
rlabel metal2 2346 3978 2346 3978 0 net1
rlabel metal1 27140 2414 27140 2414 0 net10
rlabel metal1 24697 3026 24697 3026 0 net100
rlabel metal1 14025 22678 14025 22678 0 net101
rlabel metal2 2254 21794 2254 21794 0 net102
rlabel metal1 4140 5882 4140 5882 0 net103
rlabel metal1 14991 26350 14991 26350 0 net104
rlabel metal1 12921 2346 12921 2346 0 net105
rlabel metal1 27554 10710 27554 10710 0 net106
rlabel metal1 27048 2618 27048 2618 0 net107
rlabel metal2 2254 19142 2254 19142 0 net108
rlabel metal1 13657 27030 13657 27030 0 net109
rlabel metal2 19182 17646 19182 17646 0 net11
rlabel metal1 2801 12818 2801 12818 0 net110
rlabel metal1 27503 5270 27503 5270 0 net111
rlabel metal1 3128 13430 3128 13430 0 net112
rlabel metal2 2990 15198 2990 15198 0 net113
rlabel via1 2341 5678 2341 5678 0 net114
rlabel metal2 3266 3910 3266 3910 0 net115
rlabel metal1 27186 2550 27186 2550 0 net116
rlabel metal1 2806 2992 2806 2992 0 net117
rlabel metal1 10345 3026 10345 3026 0 net118
rlabel metal1 28290 2618 28290 2618 0 net119
rlabel metal1 4278 27472 4278 27472 0 net12
rlabel metal1 8316 3026 8316 3026 0 net120
rlabel metal2 4278 4386 4278 4386 0 net121
rlabel metal2 2162 4998 2162 4998 0 net122
rlabel metal2 2162 23970 2162 23970 0 net123
rlabel metal1 7769 2346 7769 2346 0 net124
rlabel metal1 16279 23018 16279 23018 0 net125
rlabel metal1 13979 24786 13979 24786 0 net126
rlabel metal1 25893 6290 25893 6290 0 net127
rlabel metal1 12870 23698 12870 23698 0 net128
rlabel metal1 27462 12954 27462 12954 0 net129
rlabel metal1 10074 27404 10074 27404 0 net13
rlabel metal1 12594 25262 12594 25262 0 net130
rlabel metal1 13110 2448 13110 2448 0 net131
rlabel metal2 12650 26146 12650 26146 0 net132
rlabel metal1 11254 20842 11254 20842 0 net133
rlabel metal1 20093 4488 20093 4488 0 net134
rlabel metal1 2893 2346 2893 2346 0 net135
rlabel metal1 22765 3434 22765 3434 0 net136
rlabel metal2 7222 9860 7222 9860 0 net137
rlabel metal1 7217 20502 7217 20502 0 net138
rlabel metal1 20838 19720 20838 19720 0 net139
rlabel metal1 19044 26350 19044 26350 0 net14
rlabel metal1 13795 15402 13795 15402 0 net140
rlabel metal1 20787 3026 20787 3026 0 net141
rlabel metal1 24191 23698 24191 23698 0 net146
rlabel metal2 12834 4114 12834 4114 0 net147
rlabel metal2 9982 13906 9982 13906 0 net148
rlabel metal1 12737 21590 12737 21590 0 net149
rlabel metal1 21390 5338 21390 5338 0 net15
rlabel metal1 22811 16558 22811 16558 0 net150
rlabel metal1 28428 16422 28428 16422 0 net151
rlabel metal1 21344 22610 21344 22610 0 net152
rlabel metal2 23506 19346 23506 19346 0 net153
rlabel metal1 20930 6256 20930 6256 0 net154
rlabel metal1 15916 2618 15916 2618 0 net155
rlabel metal1 9471 24786 9471 24786 0 net156
rlabel metal1 2226 12138 2226 12138 0 net157
rlabel metal1 12645 4114 12645 4114 0 net158
rlabel metal2 13938 14858 13938 14858 0 net159
rlabel metal1 28566 25296 28566 25296 0 net16
rlabel metal1 20787 10710 20787 10710 0 net160
rlabel metal1 20925 11798 20925 11798 0 net161
rlabel metal1 2226 7786 2226 7786 0 net162
rlabel metal1 17981 6290 17981 6290 0 net163
rlabel metal1 22995 6358 22995 6358 0 net164
rlabel metal1 7452 22202 7452 22202 0 net165
rlabel metal1 10396 13158 10396 13158 0 net166
rlabel metal1 23133 14994 23133 14994 0 net167
rlabel metal2 22310 16048 22310 16048 0 net168
rlabel metal2 4738 12002 4738 12002 0 net169
rlabel metal1 1610 27098 1610 27098 0 net17
rlabel metal1 18257 18734 18257 18734 0 net170
rlabel metal1 8781 7378 8781 7378 0 net171
rlabel metal1 26123 17238 26123 17238 0 net172
rlabel metal1 14290 3434 14290 3434 0 net173
rlabel metal1 23823 24854 23823 24854 0 net174
rlabel metal1 27641 23766 27641 23766 0 net175
rlabel via1 24973 23086 24973 23086 0 net176
rlabel metal1 5745 25194 5745 25194 0 net177
rlabel metal2 7590 14178 7590 14178 0 net178
rlabel metal1 11454 5338 11454 5338 0 net179
rlabel metal2 28382 16082 28382 16082 0 net18
rlabel metal2 4922 10438 4922 10438 0 net180
rlabel metal1 18492 2550 18492 2550 0 net181
rlabel via1 22121 24786 22121 24786 0 net182
rlabel metal1 14296 16558 14296 16558 0 net183
rlabel metal2 26496 12988 26496 12988 0 net184
rlabel metal1 17337 2414 17337 2414 0 net185
rlabel metal2 12466 24616 12466 24616 0 net186
rlabel metal1 12328 16762 12328 16762 0 net187
rlabel metal1 25617 12886 25617 12886 0 net188
rlabel metal1 24053 5270 24053 5270 0 net189
rlabel metal1 28014 26554 28014 26554 0 net19
rlabel via1 9609 20434 9609 20434 0 net190
rlabel metal2 3542 9894 3542 9894 0 net191
rlabel metal2 17342 18870 17342 18870 0 net192
rlabel viali 25709 18326 25709 18326 0 net193
rlabel metal2 26818 23970 26818 23970 0 net194
rlabel metal1 19959 13974 19959 13974 0 net195
rlabel metal1 13662 13498 13662 13498 0 net196
rlabel metal1 11408 18938 11408 18938 0 net197
rlabel metal1 15911 3026 15911 3026 0 net198
rlabel metal1 14766 2618 14766 2618 0 net2
rlabel metal1 2714 25908 2714 25908 0 net20
rlabel metal1 10897 25262 10897 25262 0 net200
rlabel metal2 5566 13906 5566 13906 0 net201
rlabel metal2 12466 7378 12466 7378 0 net202
rlabel metal1 7493 25262 7493 25262 0 net203
rlabel metal1 20695 4114 20695 4114 0 net204
rlabel metal1 20281 17646 20281 17646 0 net205
rlabel metal1 6067 11730 6067 11730 0 net206
rlabel metal1 5980 24378 5980 24378 0 net207
rlabel metal1 16698 14926 16698 14926 0 net21
rlabel metal2 12558 12716 12558 12716 0 net22
rlabel metal1 16054 21522 16054 21522 0 net23
rlabel metal2 19274 4420 19274 4420 0 net24
rlabel metal1 25714 19414 25714 19414 0 net25
rlabel via2 2622 27013 2622 27013 0 net26
rlabel metal1 18032 9622 18032 9622 0 net27
rlabel metal1 14076 19890 14076 19890 0 net28
rlabel metal2 17526 11407 17526 11407 0 net29
rlabel metal1 27140 21658 27140 21658 0 net3
rlabel metal1 14306 11662 14306 11662 0 net30
rlabel metal1 18216 13294 18216 13294 0 net31
rlabel metal2 16146 14926 16146 14926 0 net32
rlabel metal1 18538 7752 18538 7752 0 net33
rlabel metal1 14812 17646 14812 17646 0 net34
rlabel metal1 17388 7718 17388 7718 0 net35
rlabel metal1 15042 18734 15042 18734 0 net36
rlabel metal2 21574 20995 21574 20995 0 net37
rlabel metal1 13110 18088 13110 18088 0 net38
rlabel metal2 21068 20876 21068 20876 0 net39
rlabel metal1 18032 11118 18032 11118 0 net4
rlabel metal1 21528 20978 21528 20978 0 net40
rlabel metal1 21850 15028 21850 15028 0 net41
rlabel metal1 15594 16626 15594 16626 0 net42
rlabel metal1 20838 16694 20838 16694 0 net43
rlabel metal2 20838 7038 20838 7038 0 net44
rlabel metal2 19366 15980 19366 15980 0 net45
rlabel metal2 21574 6273 21574 6273 0 net46
rlabel metal1 20102 16592 20102 16592 0 net47
rlabel metal1 27370 26452 27370 26452 0 net48
rlabel metal1 24472 26962 24472 26962 0 net49
rlabel metal1 1748 24786 1748 24786 0 net5
rlabel metal1 16882 20434 16882 20434 0 net50
rlabel metal1 11270 27540 11270 27540 0 net51
rlabel metal1 4922 27030 4922 27030 0 net52
rlabel metal2 12926 20128 12926 20128 0 net53
rlabel metal1 15502 13940 15502 13940 0 net54
rlabel metal2 6394 15334 6394 15334 0 net55
rlabel metal2 2990 9180 2990 9180 0 net56
rlabel metal1 10258 9554 10258 9554 0 net57
rlabel metal1 13386 5746 13386 5746 0 net58
rlabel metal1 16790 2992 16790 2992 0 net59
rlabel metal1 1518 25262 1518 25262 0 net6
rlabel metal1 25668 6834 25668 6834 0 net60
rlabel metal1 20424 12818 20424 12818 0 net61
rlabel metal1 25990 14042 25990 14042 0 net62
rlabel metal1 28060 18258 28060 18258 0 net63
rlabel metal2 22402 20672 22402 20672 0 net64
rlabel metal1 8648 20842 8648 20842 0 net65
rlabel metal1 1794 11662 1794 11662 0 net66
rlabel metal2 23874 2533 23874 2533 0 net67
rlabel metal1 22581 4114 22581 4114 0 net68
rlabel metal1 25617 7854 25617 7854 0 net69
rlabel metal1 19182 17102 19182 17102 0 net7
rlabel metal2 13294 21522 13294 21522 0 net70
rlabel metal2 2622 20706 2622 20706 0 net71
rlabel metal1 20373 27030 20373 27030 0 net72
rlabel metal1 6435 3094 6435 3094 0 net73
rlabel metal1 7263 7446 7263 7446 0 net74
rlabel metal2 17342 3689 17342 3689 0 net75
rlabel metal1 7907 20842 7907 20842 0 net76
rlabel metal1 21201 11050 21201 11050 0 net77
rlabel metal1 18671 27030 18671 27030 0 net78
rlabel metal1 19821 20842 19821 20842 0 net79
rlabel metal1 17296 7514 17296 7514 0 net8
rlabel metal1 17199 26962 17199 26962 0 net80
rlabel metal1 3358 19788 3358 19788 0 net81
rlabel metal2 2254 15878 2254 15878 0 net82
rlabel metal1 3215 16490 3215 16490 0 net83
rlabel metal1 5653 20910 5653 20910 0 net84
rlabel metal1 26767 8874 26767 8874 0 net85
rlabel metal1 2019 18326 2019 18326 0 net86
rlabel metal1 17291 21998 17291 21998 0 net87
rlabel metal2 3542 23868 3542 23868 0 net88
rlabel metal1 18441 21522 18441 21522 0 net89
rlabel metal2 6026 2329 6026 2329 0 net9
rlabel metal1 6716 6426 6716 6426 0 net90
rlabel metal1 26215 10710 26215 10710 0 net91
rlabel metal1 15865 26962 15865 26962 0 net92
rlabel metal1 4181 23018 4181 23018 0 net93
rlabel metal2 22494 18530 22494 18530 0 net94
rlabel metal2 2346 17442 2346 17442 0 net95
rlabel metal1 4779 6290 4779 6290 0 net96
rlabel metal2 3358 22882 3358 22882 0 net97
rlabel metal1 27181 5678 27181 5678 0 net98
rlabel metal1 22765 3026 22765 3026 0 net99
rlabel metal3 1717 6052 1717 6052 0 prog_clk
rlabel metal3 1004 16660 1004 16660 0 reset
rlabel metal3 17319 7004 17319 7004 0 right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal1 6256 2414 6256 2414 0 right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal1 28612 7854 28612 7854 0 right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal1 27784 16762 27784 16762 0 right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal3 820 13124 820 13124 0 set
rlabel metal1 3956 27438 3956 27438 0 top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal1 11730 27472 11730 27472 0 top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal1 20010 27472 20010 27472 0 top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal1 26404 27574 26404 27574 0 top_width_0_height_0_subtile_0__pin_O_2_
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
