magic
tech sky130A
magscale 1 2
timestamp 1708041521
<< viali >>
rect 13829 13481 13863 13515
rect 2329 13413 2363 13447
rect 5181 13413 5215 13447
rect 12173 13413 12207 13447
rect 14105 13413 14139 13447
rect 5365 13345 5399 13379
rect 1685 13277 1719 13311
rect 1777 13277 1811 13311
rect 2145 13277 2179 13311
rect 2513 13277 2547 13311
rect 2789 13277 2823 13311
rect 3065 13277 3099 13311
rect 3341 13277 3375 13311
rect 3985 13277 4019 13311
rect 4077 13277 4111 13311
rect 4353 13277 4387 13311
rect 4813 13277 4847 13311
rect 5273 13277 5307 13311
rect 5549 13277 5583 13311
rect 6552 13277 6586 13311
rect 6653 13277 6687 13311
rect 8033 13277 8067 13311
rect 9413 13277 9447 13311
rect 10977 13277 11011 13311
rect 12357 13277 12391 13311
rect 13185 13277 13219 13311
rect 14289 13277 14323 13311
rect 13553 13209 13587 13243
rect 1593 13141 1627 13175
rect 1869 13141 1903 13175
rect 2697 13141 2731 13175
rect 2973 13141 3007 13175
rect 3249 13141 3283 13175
rect 3433 13141 3467 13175
rect 3801 13141 3835 13175
rect 4169 13141 4203 13175
rect 4537 13141 4571 13175
rect 4997 13141 5031 13175
rect 6009 13141 6043 13175
rect 6377 13141 6411 13175
rect 6837 13141 6871 13175
rect 8217 13141 8251 13175
rect 9597 13141 9631 13175
rect 10793 13141 10827 13175
rect 13093 13141 13127 13175
rect 4537 12937 4571 12971
rect 6837 12937 6871 12971
rect 5457 12869 5491 12903
rect 6009 12869 6043 12903
rect 7481 12869 7515 12903
rect 1777 12801 1811 12835
rect 2053 12801 2087 12835
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 3709 12801 3743 12835
rect 3893 12801 3927 12835
rect 4169 12801 4203 12835
rect 4445 12801 4479 12835
rect 4721 12801 4755 12835
rect 6377 12801 6411 12835
rect 6653 12801 6687 12835
rect 11796 12801 11830 12835
rect 13185 12801 13219 12835
rect 14197 12801 14231 12835
rect 14473 12801 14507 12835
rect 2237 12733 2271 12767
rect 4905 12733 4939 12767
rect 5365 12733 5399 12767
rect 6101 12733 6135 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 11529 12733 11563 12767
rect 13369 12733 13403 12767
rect 4077 12665 4111 12699
rect 4353 12665 4387 12699
rect 6561 12665 6595 12699
rect 7021 12665 7055 12699
rect 14289 12665 14323 12699
rect 1501 12597 1535 12631
rect 2697 12597 2731 12631
rect 2789 12597 2823 12631
rect 3617 12597 3651 12631
rect 12909 12597 12943 12631
rect 13829 12597 13863 12631
rect 14013 12597 14047 12631
rect 1593 12393 1627 12427
rect 2421 12393 2455 12427
rect 6377 12393 6411 12427
rect 13093 12393 13127 12427
rect 4629 12325 4663 12359
rect 6193 12325 6227 12359
rect 2237 12257 2271 12291
rect 2973 12257 3007 12291
rect 3341 12257 3375 12291
rect 12909 12257 12943 12291
rect 1409 12189 1443 12223
rect 2605 12189 2639 12223
rect 4353 12189 4387 12223
rect 4721 12189 4755 12223
rect 4813 12189 4847 12223
rect 6469 12199 6503 12233
rect 6653 12189 6687 12223
rect 13001 12189 13035 12223
rect 13277 12189 13311 12223
rect 13737 12189 13771 12223
rect 14105 12189 14139 12223
rect 3249 12121 3283 12155
rect 5080 12121 5114 12155
rect 1685 12053 1719 12087
rect 3801 12053 3835 12087
rect 7941 12053 7975 12087
rect 12265 12053 12299 12087
rect 13369 12053 13403 12087
rect 13921 12053 13955 12087
rect 14197 12053 14231 12087
rect 2973 11849 3007 11883
rect 4445 11849 4479 11883
rect 5457 11849 5491 11883
rect 11529 11849 11563 11883
rect 3332 11781 3366 11815
rect 9536 11781 9570 11815
rect 10425 11781 10459 11815
rect 10517 11781 10551 11815
rect 12725 11781 12759 11815
rect 13461 11781 13495 11815
rect 1593 11713 1627 11747
rect 1849 11713 1883 11747
rect 4813 11713 4847 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 13921 11713 13955 11747
rect 14105 11713 14139 11747
rect 14197 11713 14231 11747
rect 3065 11645 3099 11679
rect 6193 11645 6227 11679
rect 7941 11645 7975 11679
rect 9781 11645 9815 11679
rect 13185 11645 13219 11679
rect 13369 11645 13403 11679
rect 8401 11577 8435 11611
rect 9965 11577 9999 11611
rect 14289 11577 14323 11611
rect 5549 11509 5583 11543
rect 12633 11509 12667 11543
rect 1409 11305 1443 11339
rect 3065 11305 3099 11339
rect 9597 11305 9631 11339
rect 13553 11305 13587 11339
rect 4445 11237 4479 11271
rect 7297 11237 7331 11271
rect 2789 11169 2823 11203
rect 7941 11169 7975 11203
rect 8309 11169 8343 11203
rect 11345 11169 11379 11203
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 9505 11101 9539 11135
rect 11612 11101 11646 11135
rect 13369 11101 13403 11135
rect 13737 11101 13771 11135
rect 14473 11101 14507 11135
rect 2544 11033 2578 11067
rect 3617 11033 3651 11067
rect 3893 11033 3927 11067
rect 3985 11033 4019 11067
rect 8033 11033 8067 11067
rect 3341 10965 3375 10999
rect 7757 10965 7791 10999
rect 12725 10965 12759 10999
rect 12817 10965 12851 10999
rect 14289 10965 14323 10999
rect 2881 10761 2915 10795
rect 14013 10761 14047 10795
rect 4353 10693 4387 10727
rect 7849 10693 7883 10727
rect 11796 10693 11830 10727
rect 1777 10625 1811 10659
rect 9597 10625 9631 10659
rect 11529 10625 11563 10659
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 1501 10421 1535 10455
rect 12909 10421 12943 10455
rect 13185 10421 13219 10455
rect 1777 10013 1811 10047
rect 3065 10013 3099 10047
rect 11529 10013 11563 10047
rect 11805 10013 11839 10047
rect 13737 10013 13771 10047
rect 14473 10013 14507 10047
rect 12173 9945 12207 9979
rect 12265 9945 12299 9979
rect 12817 9945 12851 9979
rect 12909 9945 12943 9979
rect 13461 9945 13495 9979
rect 13553 9945 13587 9979
rect 1593 9877 1627 9911
rect 2973 9877 3007 9911
rect 11713 9877 11747 9911
rect 11989 9877 12023 9911
rect 13921 9877 13955 9911
rect 14289 9877 14323 9911
rect 12265 9673 12299 9707
rect 12909 9673 12943 9707
rect 13737 9673 13771 9707
rect 1777 9537 1811 9571
rect 12817 9537 12851 9571
rect 13645 9537 13679 9571
rect 14197 9537 14231 9571
rect 14381 9469 14415 9503
rect 13461 9401 13495 9435
rect 1501 9333 1535 9367
rect 14197 9129 14231 9163
rect 14289 8925 14323 8959
rect 1961 8585 1995 8619
rect 1777 8449 1811 8483
rect 2145 8449 2179 8483
rect 14473 8449 14507 8483
rect 1501 8313 1535 8347
rect 14289 8245 14323 8279
rect 2053 7497 2087 7531
rect 2329 7497 2363 7531
rect 1777 7429 1811 7463
rect 2237 7361 2271 7395
rect 2513 7361 2547 7395
rect 1501 7157 1535 7191
rect 14289 6953 14323 6987
rect 14473 6749 14507 6783
rect 1777 6273 1811 6307
rect 14197 6273 14231 6307
rect 14013 6137 14047 6171
rect 1501 6069 1535 6103
rect 14473 5661 14507 5695
rect 14289 5525 14323 5559
rect 1777 5253 1811 5287
rect 1501 4981 1535 5015
rect 1777 4097 1811 4131
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 14473 4097 14507 4131
rect 1501 3893 1535 3927
rect 14289 3893 14323 3927
rect 13921 3145 13955 3179
rect 14105 3077 14139 3111
rect 1777 3009 1811 3043
rect 6929 3009 6963 3043
rect 13737 3009 13771 3043
rect 1501 2805 1535 2839
rect 7113 2805 7147 2839
rect 14381 2805 14415 2839
rect 1685 2601 1719 2635
rect 14289 2601 14323 2635
rect 9505 2533 9539 2567
rect 1777 2397 1811 2431
rect 2973 2397 3007 2431
rect 4721 2397 4755 2431
rect 6101 2397 6135 2431
rect 6377 2397 6411 2431
rect 7665 2397 7699 2431
rect 8217 2397 8251 2431
rect 9689 2397 9723 2431
rect 14473 2397 14507 2431
rect 2605 2329 2639 2363
rect 4169 2329 4203 2363
rect 4537 2329 4571 2363
rect 5733 2329 5767 2363
rect 7297 2329 7331 2363
rect 9045 2329 9079 2363
rect 10517 2329 10551 2363
rect 12081 2329 12115 2363
rect 13553 2329 13587 2363
rect 4905 2261 4939 2295
rect 6561 2261 6595 2295
rect 8401 2261 8435 2295
rect 9137 2261 9171 2295
rect 10609 2261 10643 2295
rect 12173 2261 12207 2295
rect 13829 2261 13863 2295
<< metal1 >>
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2096 13484 4016 13512
rect 2096 13472 2102 13484
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 2363 13416 3372 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 1302 13336 1308 13388
rect 1360 13376 1366 13388
rect 1360 13348 2636 13376
rect 1360 13336 1366 13348
rect 1026 13268 1032 13320
rect 1084 13268 1090 13320
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 2038 13308 2044 13320
rect 1811 13280 2044 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 1044 13240 1072 13268
rect 2148 13240 2176 13271
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2464 13280 2513 13308
rect 2464 13268 2470 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 2608 13308 2636 13348
rect 3344 13317 3372 13416
rect 3988 13317 4016 13484
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13780 13484 13829 13512
rect 13780 13472 13786 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13413 5227 13447
rect 12161 13447 12219 13453
rect 12161 13444 12173 13447
rect 5169 13407 5227 13413
rect 5460 13416 12173 13444
rect 5184 13376 5212 13407
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 5184 13348 5365 13376
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2608 13280 2789 13308
rect 2501 13271 2559 13277
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 3068 13240 3096 13271
rect 4080 13240 4108 13271
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4212 13280 4353 13308
rect 4212 13268 4218 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5166 13308 5172 13320
rect 4847 13280 5172 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5460 13308 5488 13416
rect 12161 13413 12173 13416
rect 12207 13413 12219 13447
rect 12161 13407 12219 13413
rect 14093 13447 14151 13453
rect 14093 13413 14105 13447
rect 14139 13413 14151 13447
rect 14093 13407 14151 13413
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6512 13348 6684 13376
rect 6512 13336 6518 13348
rect 5307 13280 5488 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 6656 13317 6684 13348
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 14108 13376 14136 13407
rect 6788 13348 11100 13376
rect 6788 13336 6794 13348
rect 6540 13311 6598 13317
rect 6540 13277 6552 13311
rect 6586 13277 6598 13311
rect 6540 13271 6598 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 1044 13212 2176 13240
rect 2700 13212 3096 13240
rect 3160 13212 4108 13240
rect 6564 13240 6592 13271
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 7984 13280 8033 13308
rect 7984 13268 7990 13280
rect 8021 13277 8033 13280
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 9401 13311 9459 13317
rect 9401 13308 9413 13311
rect 9364 13280 9413 13308
rect 9364 13268 9370 13280
rect 9401 13277 9413 13280
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10744 13280 10977 13308
rect 10744 13268 10750 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11072 13240 11100 13348
rect 13188 13348 14136 13376
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 13188 13317 13216 13348
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12124 13280 12357 13308
rect 12124 13268 12130 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13504 13280 14289 13308
rect 13504 13268 13510 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 6564 13212 10824 13240
rect 11072 13212 13553 13240
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 1854 13132 1860 13184
rect 1912 13132 1918 13184
rect 2700 13181 2728 13212
rect 2685 13175 2743 13181
rect 2685 13141 2697 13175
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3160 13172 3188 13212
rect 3007 13144 3188 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 3234 13132 3240 13184
rect 3292 13132 3298 13184
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 3786 13132 3792 13184
rect 3844 13132 3850 13184
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 4706 13172 4712 13184
rect 4571 13144 4712 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4985 13175 5043 13181
rect 4985 13141 4997 13175
rect 5031 13172 5043 13175
rect 5718 13172 5724 13184
rect 5031 13144 5724 13172
rect 5031 13141 5043 13144
rect 4985 13135 5043 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5868 13144 6009 13172
rect 5868 13132 5874 13144
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6144 13144 6377 13172
rect 6144 13132 6150 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 6822 13132 6828 13184
rect 6880 13132 6886 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7708 13144 8217 13172
rect 7708 13132 7714 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 8205 13135 8263 13141
rect 9585 13175 9643 13181
rect 9585 13141 9597 13175
rect 9631 13172 9643 13175
rect 9858 13172 9864 13184
rect 9631 13144 9864 13172
rect 9631 13141 9643 13144
rect 9585 13135 9643 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10796 13181 10824 13212
rect 13541 13209 13553 13212
rect 13587 13209 13599 13243
rect 13541 13203 13599 13209
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13141 10839 13175
rect 10781 13135 10839 13141
rect 13078 13132 13084 13184
rect 13136 13132 13142 13184
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1578 12928 1584 12980
rect 1636 12928 1642 12980
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 1912 12940 2774 12968
rect 1912 12928 1918 12940
rect 1596 12900 1624 12928
rect 1596 12872 2084 12900
rect 1762 12792 1768 12844
rect 1820 12792 1826 12844
rect 2056 12841 2084 12872
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2746 12832 2774 12940
rect 3418 12928 3424 12980
rect 3476 12928 3482 12980
rect 4154 12928 4160 12980
rect 4212 12928 4218 12980
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 5534 12968 5540 12980
rect 4571 12940 5540 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 3436 12841 3464 12928
rect 4172 12900 4200 12928
rect 5445 12903 5503 12909
rect 4172 12872 4752 12900
rect 4724 12841 4752 12872
rect 5445 12869 5457 12903
rect 5491 12900 5503 12903
rect 5626 12900 5632 12912
rect 5491 12872 5632 12900
rect 5491 12869 5503 12872
rect 5445 12863 5503 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 5994 12860 6000 12912
rect 6052 12860 6058 12912
rect 6730 12900 6736 12912
rect 6380 12872 6736 12900
rect 6380 12841 6408 12872
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 6840 12900 6868 12931
rect 13078 12928 13084 12980
rect 13136 12928 13142 12980
rect 14458 12928 14464 12980
rect 14516 12928 14522 12980
rect 14550 12928 14556 12980
rect 14608 12928 14614 12980
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 6840 12872 7481 12900
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 7469 12863 7527 12869
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 2746 12804 3249 12832
rect 2041 12795 2099 12801
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3927 12804 4016 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 2222 12724 2228 12776
rect 2280 12724 2286 12776
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3712 12764 3740 12795
rect 3108 12736 3740 12764
rect 3108 12724 3114 12736
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 2685 12631 2743 12637
rect 2685 12597 2697 12631
rect 2731 12628 2743 12631
rect 2777 12631 2835 12637
rect 2777 12628 2789 12631
rect 2731 12600 2789 12628
rect 2731 12597 2743 12600
rect 2685 12591 2743 12597
rect 2777 12597 2789 12600
rect 2823 12628 2835 12631
rect 3142 12628 3148 12640
rect 2823 12600 3148 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3234 12588 3240 12640
rect 3292 12628 3298 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3292 12600 3617 12628
rect 3292 12588 3298 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 3988 12628 4016 12804
rect 4080 12804 4169 12832
rect 4080 12705 4108 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4157 12795 4215 12801
rect 4264 12804 4445 12832
rect 4264 12708 4292 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6365 12795 6423 12801
rect 6564 12804 6653 12832
rect 4893 12767 4951 12773
rect 4893 12733 4905 12767
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12764 5411 12767
rect 5810 12764 5816 12776
rect 5399 12736 5816 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12665 4123 12699
rect 4065 12659 4123 12665
rect 4246 12656 4252 12708
rect 4304 12656 4310 12708
rect 4341 12699 4399 12705
rect 4341 12665 4353 12699
rect 4387 12696 4399 12699
rect 4908 12696 4936 12727
rect 5810 12724 5816 12736
rect 5868 12764 5874 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5868 12736 6101 12764
rect 5868 12724 5874 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 6564 12705 6592 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 11784 12835 11842 12841
rect 11784 12801 11796 12835
rect 11830 12832 11842 12835
rect 13096 12832 13124 12928
rect 14476 12900 14504 12928
rect 14200 12872 14504 12900
rect 14200 12841 14228 12872
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 11830 12804 13032 12832
rect 13096 12804 13185 12832
rect 11830 12801 11842 12804
rect 11784 12795 11842 12801
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7607 12736 7757 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 4387 12668 4936 12696
rect 6549 12699 6607 12705
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 6549 12665 6561 12699
rect 6595 12665 6607 12699
rect 6549 12659 6607 12665
rect 7009 12699 7067 12705
rect 7009 12665 7021 12699
rect 7055 12665 7067 12699
rect 13004 12696 13032 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14568 12832 14596 12928
rect 14507 12804 14596 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14277 12699 14335 12705
rect 14277 12696 14289 12699
rect 13004 12668 14289 12696
rect 7009 12659 7067 12665
rect 14277 12665 14289 12668
rect 14323 12665 14335 12699
rect 14277 12659 14335 12665
rect 4264 12628 4292 12656
rect 3988 12600 4292 12628
rect 3605 12591 3663 12597
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 7024 12628 7052 12659
rect 5684 12600 7052 12628
rect 5684 12588 5690 12600
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12768 12600 12909 12628
rect 12768 12588 12774 12600
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 12897 12591 12955 12597
rect 13814 12588 13820 12640
rect 13872 12588 13878 12640
rect 13998 12588 14004 12640
rect 14056 12588 14062 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1670 12424 1676 12436
rect 1627 12396 1676 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2280 12396 2421 12424
rect 2280 12384 2286 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 6052 12396 6377 12424
rect 6052 12384 6058 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 6730 12384 6736 12436
rect 6788 12384 6794 12436
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13354 12424 13360 12436
rect 13127 12396 13360 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 3786 12356 3792 12368
rect 2608 12328 3792 12356
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2225 12291 2283 12297
rect 2225 12288 2237 12291
rect 2096 12260 2237 12288
rect 2096 12248 2102 12260
rect 2225 12257 2237 12260
rect 2271 12257 2283 12291
rect 2225 12251 2283 12257
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 2608 12229 2636 12328
rect 3786 12316 3792 12328
rect 3844 12316 3850 12368
rect 4617 12359 4675 12365
rect 4617 12325 4629 12359
rect 4663 12356 4675 12359
rect 4798 12356 4804 12368
rect 4663 12328 4804 12356
rect 4663 12325 4675 12328
rect 4617 12319 4675 12325
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 6181 12359 6239 12365
rect 6181 12325 6193 12359
rect 6227 12356 6239 12359
rect 6748 12356 6776 12384
rect 6227 12328 6776 12356
rect 6227 12325 6239 12328
rect 6181 12319 6239 12325
rect 2958 12248 2964 12300
rect 3016 12248 3022 12300
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3329 12291 3387 12297
rect 3329 12288 3341 12291
rect 3200 12260 3341 12288
rect 3200 12248 3206 12260
rect 3329 12257 3341 12260
rect 3375 12257 3387 12291
rect 3329 12251 3387 12257
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4120 12260 4936 12288
rect 4120 12248 4126 12260
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 3568 12192 4353 12220
rect 3568 12180 3574 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4341 12183 4399 12189
rect 4540 12192 4721 12220
rect 3234 12112 3240 12164
rect 3292 12112 3298 12164
rect 1670 12044 1676 12096
rect 1728 12044 1734 12096
rect 3786 12044 3792 12096
rect 3844 12044 3850 12096
rect 4540 12084 4568 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4908 12220 4936 12260
rect 6472 12239 6500 12328
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 12768 12260 12909 12288
rect 12768 12248 12774 12260
rect 12897 12257 12909 12260
rect 12943 12288 12955 12291
rect 12943 12260 13032 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 6457 12233 6515 12239
rect 4908 12192 5212 12220
rect 6457 12199 6469 12233
rect 6503 12199 6515 12233
rect 13004 12229 13032 12260
rect 13740 12260 14596 12288
rect 6457 12193 6515 12199
rect 6641 12223 6699 12229
rect 4801 12183 4859 12189
rect 4816 12152 4844 12183
rect 4890 12152 4896 12164
rect 4816 12124 4896 12152
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5074 12161 5080 12164
rect 5068 12115 5080 12161
rect 5074 12112 5080 12115
rect 5132 12112 5138 12164
rect 5184 12152 5212 12192
rect 6641 12189 6653 12223
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 6656 12152 6684 12183
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13740 12229 13768 12260
rect 14568 12232 14596 12260
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 13136 12192 13277 12220
rect 13136 12180 13142 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 14056 12192 14105 12220
rect 14056 12180 14062 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 5184 12124 6684 12152
rect 5534 12084 5540 12096
rect 4540 12056 5540 12084
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7708 12056 7941 12084
rect 7708 12044 7714 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11940 12056 12265 12084
rect 11940 12044 11946 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 13906 12044 13912 12096
rect 13964 12044 13970 12096
rect 14182 12044 14188 12096
rect 14240 12044 14246 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3142 11880 3148 11892
rect 3007 11852 3148 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3142 11840 3148 11852
rect 3200 11880 3206 11892
rect 3510 11880 3516 11892
rect 3200 11852 3516 11880
rect 3200 11840 3206 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3786 11840 3792 11892
rect 3844 11840 3850 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4304 11852 4445 11880
rect 4304 11840 4310 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 3320 11815 3378 11821
rect 1596 11784 2774 11812
rect 1596 11753 1624 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1670 11704 1676 11756
rect 1728 11744 1734 11756
rect 1837 11747 1895 11753
rect 1837 11744 1849 11747
rect 1728 11716 1849 11744
rect 1728 11704 1734 11716
rect 1837 11713 1849 11716
rect 1883 11713 1895 11747
rect 2746 11744 2774 11784
rect 3320 11781 3332 11815
rect 3366 11812 3378 11815
rect 3804 11812 3832 11840
rect 3366 11784 3832 11812
rect 3366 11781 3378 11784
rect 3320 11775 3378 11781
rect 4448 11744 4476 11843
rect 4890 11840 4896 11892
rect 4948 11840 4954 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5132 11852 5457 11880
rect 5132 11840 5138 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 5445 11843 5503 11849
rect 10336 11852 11529 11880
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 2746 11716 4108 11744
rect 4448 11716 4813 11744
rect 1837 11707 1895 11713
rect 3068 11688 3096 11716
rect 3050 11636 3056 11688
rect 3108 11636 3114 11688
rect 4080 11676 4108 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4908 11676 4936 11840
rect 9524 11815 9582 11821
rect 9524 11781 9536 11815
rect 9570 11812 9582 11815
rect 10336 11812 10364 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13412 11852 13676 11880
rect 13412 11840 13418 11852
rect 9570 11784 10364 11812
rect 9570 11781 9582 11784
rect 9524 11775 9582 11781
rect 10410 11772 10416 11824
rect 10468 11772 10474 11824
rect 10505 11815 10563 11821
rect 10505 11781 10517 11815
rect 10551 11812 10563 11815
rect 12713 11815 12771 11821
rect 12713 11812 12725 11815
rect 10551 11784 12725 11812
rect 10551 11781 10563 11784
rect 10505 11775 10563 11781
rect 12713 11781 12725 11784
rect 12759 11812 12771 11815
rect 13449 11815 13507 11821
rect 13449 11812 13461 11815
rect 12759 11784 13461 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 13449 11781 13461 11784
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 12207 11716 12449 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 12437 11713 12449 11716
rect 12483 11744 12495 11747
rect 12802 11744 12808 11756
rect 12483 11716 12808 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 13078 11744 13084 11756
rect 12860 11716 13084 11744
rect 12860 11704 12866 11716
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13648 11744 13676 11852
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 13964 11852 14044 11880
rect 13964 11840 13970 11852
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13648 11716 13921 11744
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 4080 11648 4936 11676
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 7006 11676 7012 11688
rect 6227 11648 7012 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7926 11636 7932 11688
rect 7984 11636 7990 11688
rect 9769 11679 9827 11685
rect 9769 11645 9781 11679
rect 9815 11676 9827 11679
rect 9815 11648 10456 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 7024 11608 7052 11636
rect 8386 11608 8392 11620
rect 7024 11580 8392 11608
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11577 10011 11611
rect 10428 11608 10456 11648
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 13262 11676 13268 11688
rect 13219 11648 13268 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11645 13415 11679
rect 14016 11676 14044 11852
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 14200 11812 14228 11840
rect 14108 11784 14228 11812
rect 14108 11753 14136 11784
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14200 11676 14228 11707
rect 14016 11648 14228 11676
rect 13357 11639 13415 11645
rect 11624 11608 11652 11636
rect 10428 11580 11652 11608
rect 13372 11608 13400 11639
rect 14277 11611 14335 11617
rect 14277 11608 14289 11611
rect 13372 11580 14289 11608
rect 9953 11571 10011 11577
rect 14277 11577 14289 11580
rect 14323 11577 14335 11611
rect 14277 11571 14335 11577
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3418 11540 3424 11552
rect 3016 11512 3424 11540
rect 3016 11500 3022 11512
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 5534 11500 5540 11552
rect 5592 11500 5598 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9968 11540 9996 11571
rect 8168 11512 9996 11540
rect 8168 11500 8174 11512
rect 12618 11500 12624 11552
rect 12676 11500 12682 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 2038 11336 2044 11348
rect 1443 11308 2044 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2958 11296 2964 11348
rect 3016 11296 3022 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11305 3111 11339
rect 3053 11299 3111 11305
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2976 11200 3004 11296
rect 3068 11268 3096 11299
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 7006 11296 7012 11348
rect 7064 11296 7070 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 9585 11339 9643 11345
rect 9585 11305 9597 11339
rect 9631 11336 9643 11339
rect 10410 11336 10416 11348
rect 9631 11308 10416 11336
rect 9631 11305 9643 11308
rect 9585 11299 9643 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 11606 11336 11612 11348
rect 11348 11308 11612 11336
rect 3068 11240 3188 11268
rect 2832 11172 3004 11200
rect 2832 11160 2838 11172
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3160 11141 3188 11240
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 4433 11271 4491 11277
rect 4433 11268 4445 11271
rect 3476 11240 4445 11268
rect 3476 11228 3482 11240
rect 4433 11237 4445 11240
rect 4479 11237 4491 11271
rect 4433 11231 4491 11237
rect 5552 11200 5580 11296
rect 3528 11172 5580 11200
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11101 3203 11135
rect 3145 11095 3203 11101
rect 2532 11067 2590 11073
rect 2532 11033 2544 11067
rect 2578 11064 2590 11067
rect 3528 11064 3556 11172
rect 7024 11132 7052 11296
rect 7285 11271 7343 11277
rect 7285 11237 7297 11271
rect 7331 11237 7343 11271
rect 8110 11268 8116 11280
rect 7285 11231 7343 11237
rect 7392 11240 8116 11268
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 7024 11104 7113 11132
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7300 11132 7328 11231
rect 7392 11212 7420 11240
rect 8110 11228 8116 11240
rect 8168 11268 8174 11280
rect 8168 11240 8340 11268
rect 8168 11228 8174 11240
rect 7374 11160 7380 11212
rect 7432 11160 7438 11212
rect 7926 11160 7932 11212
rect 7984 11160 7990 11212
rect 8312 11209 8340 11240
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 8404 11200 8432 11296
rect 11348 11209 11376 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12618 11296 12624 11348
rect 12676 11296 12682 11348
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13320 11308 13553 11336
rect 13320 11296 13326 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 11333 11203 11391 11209
rect 8404 11172 9536 11200
rect 8297 11163 8355 11169
rect 9508 11141 9536 11172
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 12636 11200 12664 11296
rect 12636 11172 13768 11200
rect 11333 11163 11391 11169
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7300 11104 7573 11132
rect 7101 11095 7159 11101
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 11600 11135 11658 11141
rect 11600 11101 11612 11135
rect 11646 11132 11658 11135
rect 11882 11132 11888 11144
rect 11646 11104 11888 11132
rect 11646 11101 11658 11104
rect 11600 11095 11658 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 13740 11141 13768 11172
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14507 11104 14596 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 2578 11036 3556 11064
rect 3605 11067 3663 11073
rect 2578 11033 2590 11036
rect 2532 11027 2590 11033
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 3881 11067 3939 11073
rect 3881 11064 3893 11067
rect 3651 11036 3893 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 3881 11033 3893 11036
rect 3927 11033 3939 11067
rect 3881 11027 3939 11033
rect 3973 11067 4031 11073
rect 3973 11033 3985 11067
rect 4019 11033 4031 11067
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 3973 11027 4031 11033
rect 7760 11036 8033 11064
rect 3329 10999 3387 11005
rect 3329 10965 3341 10999
rect 3375 10996 3387 10999
rect 3988 10996 4016 11027
rect 7760 11005 7788 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 13372 11064 13400 11095
rect 14568 11076 14596 11104
rect 8021 11027 8079 11033
rect 12728 11036 13400 11064
rect 3375 10968 4016 10996
rect 7745 10999 7803 11005
rect 3375 10965 3387 10968
rect 3329 10959 3387 10965
rect 7745 10965 7757 10999
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 12728 11005 12756 11036
rect 14550 11024 14556 11076
rect 14608 11024 14614 11076
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12676 10968 12725 10996
rect 12676 10956 12682 10968
rect 12713 10965 12725 10968
rect 12759 10965 12771 10999
rect 12713 10959 12771 10965
rect 12802 10956 12808 11008
rect 12860 10956 12866 11008
rect 14274 10956 14280 11008
rect 14332 10956 14338 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 1762 10752 1768 10804
rect 1820 10752 1826 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2832 10764 2881 10792
rect 2832 10752 2838 10764
rect 2869 10761 2881 10764
rect 2915 10761 2927 10795
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 2869 10755 2927 10761
rect 4264 10764 14013 10792
rect 1780 10724 1808 10752
rect 4264 10724 4292 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 1780 10696 4292 10724
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 7650 10724 7656 10736
rect 4387 10696 7656 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 7650 10684 7656 10696
rect 7708 10724 7714 10736
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 7708 10696 7849 10724
rect 7708 10684 7714 10696
rect 7837 10693 7849 10696
rect 7883 10693 7895 10727
rect 7837 10687 7895 10693
rect 11784 10727 11842 10733
rect 11784 10693 11796 10727
rect 11830 10724 11842 10727
rect 12802 10724 12808 10736
rect 11830 10696 12808 10724
rect 11830 10693 11842 10696
rect 11784 10687 11842 10693
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 1762 10616 1768 10668
rect 1820 10616 1826 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 9631 10628 11529 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 11517 10625 11529 10628
rect 11563 10656 11575 10659
rect 11606 10656 11612 10668
rect 11563 10628 11612 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12768 10628 13001 10656
rect 12768 10616 12774 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 14182 10616 14188 10668
rect 14240 10616 14246 10668
rect 14274 10520 14280 10532
rect 12452 10492 14280 10520
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 992 10424 1501 10452
rect 992 10412 998 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 12452 10452 12480 10492
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 7616 10424 12480 10452
rect 7616 10412 7622 10424
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13446 10452 13452 10464
rect 13219 10424 13452 10452
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 12434 10248 12440 10260
rect 1820 10220 12440 10248
rect 1820 10208 1826 10220
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 7558 10180 7564 10192
rect 2746 10152 7564 10180
rect 2746 10112 2774 10152
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 13446 10140 13452 10192
rect 13504 10140 13510 10192
rect 3418 10112 3424 10124
rect 1780 10084 2774 10112
rect 3068 10084 3424 10112
rect 1780 10053 1808 10084
rect 3068 10053 3096 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 12618 10112 12624 10124
rect 11532 10084 12624 10112
rect 11532 10053 11560 10084
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13464 10112 13492 10140
rect 13464 10084 13768 10112
rect 13740 10053 13768 10084
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11517 10007 11575 10013
rect 11716 10016 11805 10044
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 2958 9868 2964 9920
rect 3016 9868 3022 9920
rect 11716 9917 11744 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13814 10004 13820 10056
rect 13872 10004 13878 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 14507 10016 14596 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 12158 9936 12164 9988
rect 12216 9936 12222 9988
rect 12253 9979 12311 9985
rect 12253 9945 12265 9979
rect 12299 9945 12311 9979
rect 12253 9939 12311 9945
rect 11701 9911 11759 9917
rect 11701 9877 11713 9911
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12268 9908 12296 9939
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12897 9979 12955 9985
rect 12897 9976 12909 9979
rect 12860 9948 12909 9976
rect 12860 9936 12866 9948
rect 12897 9945 12909 9948
rect 12943 9945 12955 9979
rect 12897 9939 12955 9945
rect 13446 9936 13452 9988
rect 13504 9936 13510 9988
rect 13541 9979 13599 9985
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13832 9976 13860 10004
rect 13587 9948 13860 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 14568 9920 14596 10016
rect 12023 9880 12296 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 13906 9868 13912 9920
rect 13964 9868 13970 9920
rect 14274 9868 14280 9920
rect 14332 9868 14338 9920
rect 14550 9868 14556 9920
rect 14608 9868 14614 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 12216 9676 12265 9704
rect 12216 9664 12222 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 12618 9664 12624 9716
rect 12676 9664 12682 9716
rect 12897 9707 12955 9713
rect 12897 9673 12909 9707
rect 12943 9704 12955 9707
rect 13446 9704 13452 9716
rect 12943 9676 13452 9704
rect 12943 9673 12955 9676
rect 12897 9667 12955 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13725 9707 13783 9713
rect 13725 9673 13737 9707
rect 13771 9704 13783 9707
rect 13814 9704 13820 9716
rect 13771 9676 13820 9704
rect 13771 9673 13783 9676
rect 13725 9667 13783 9673
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 12636 9568 12664 9664
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 12636 9540 12817 9568
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9568 13691 9571
rect 13814 9568 13820 9580
rect 13679 9540 13820 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13964 9540 14197 9568
rect 13964 9528 13970 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14415 9472 14872 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 12452 9432 12480 9460
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 12452 9404 13461 9432
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 1489 9367 1547 9373
rect 1489 9364 1501 9367
rect 992 9336 1501 9364
rect 992 9324 998 9336
rect 1489 9333 1501 9336
rect 1535 9333 1547 9367
rect 1489 9327 1547 9333
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14844 9160 14872 9472
rect 14231 9132 14872 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14274 8916 14280 8968
rect 14332 8916 14338 8968
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1820 8588 1961 8616
rect 1820 8576 1826 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 1949 8579 2007 8585
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2038 8480 2044 8492
rect 1811 8452 2044 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14507 8452 14964 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14936 8356 14964 8452
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 14918 8304 14924 8356
rect 14976 8304 14982 8356
rect 14274 8236 14280 8288
rect 14332 8236 14338 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 1765 7463 1823 7469
rect 1765 7429 1777 7463
rect 1811 7460 1823 7463
rect 2332 7460 2360 7491
rect 1811 7432 2360 7460
rect 1811 7429 1823 7432
rect 1765 7423 1823 7429
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 14274 7392 14280 7404
rect 2547 7364 14280 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2240 7256 2268 7355
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14274 7256 14280 7268
rect 2240 7228 14280 7256
rect 14274 7216 14280 7228
rect 14332 7216 14338 7268
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 14274 6944 14280 6996
rect 14332 6944 14338 6996
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14918 6780 14924 6792
rect 14507 6752 14924 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 1811 6276 2774 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 2746 6168 2774 6276
rect 14182 6264 14188 6316
rect 14240 6264 14246 6316
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 2746 6140 14013 6168
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14001 6131 14059 6137
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 992 6072 1501 6100
rect 992 6060 998 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1489 6063 1547 6069
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 14507 5664 14596 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 14568 5568 14596 5664
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 2188 5528 14289 5556
rect 2188 5516 2194 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14277 5519 14335 5525
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 1762 5244 1768 5296
rect 1820 5244 1826 5296
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1811 4100 2053 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 7374 4128 7380 4140
rect 2179 4100 7380 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 14507 4100 14964 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14936 4004 14964 4100
rect 14918 3952 14924 4004
rect 14976 3952 14982 4004
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 992 3896 1501 3924
rect 992 3884 998 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13872 3896 14289 3924
rect 13872 3884 13878 3896
rect 14277 3893 14289 3896
rect 14323 3893 14335 3927
rect 14277 3887 14335 3893
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 13906 3136 13912 3188
rect 13964 3136 13970 3188
rect 3694 3068 3700 3120
rect 3752 3108 3758 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 3752 3080 14105 3108
rect 3752 3068 3758 3080
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6880 3012 6929 3040
rect 6880 3000 6886 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 8846 2836 8852 2848
rect 7147 2808 8852 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 15010 2836 15016 2848
rect 14415 2808 15016 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1762 2632 1768 2644
rect 1719 2604 1768 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 14277 2635 14335 2641
rect 6886 2604 12848 2632
rect 6886 2564 6914 2604
rect 12820 2576 12848 2604
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14366 2632 14372 2644
rect 14323 2604 14372 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 1780 2536 6914 2564
rect 9493 2567 9551 2573
rect 1780 2437 1808 2536
rect 9493 2533 9505 2567
rect 9539 2533 9551 2567
rect 9493 2527 9551 2533
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 9508 2496 9536 2527
rect 12802 2524 12808 2576
rect 12860 2524 12866 2576
rect 5960 2468 6408 2496
rect 5960 2456 5966 2468
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3050 2428 3056 2440
rect 3007 2400 3056 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 4982 2388 4988 2440
rect 5040 2388 5046 2440
rect 6086 2388 6092 2440
rect 6144 2388 6150 2440
rect 6380 2437 6408 2468
rect 7668 2468 9536 2496
rect 7668 2437 7696 2468
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8846 2388 8852 2440
rect 8904 2428 8910 2440
rect 8904 2400 9168 2428
rect 8904 2388 8910 2400
rect 2590 2320 2596 2372
rect 2648 2320 2654 2372
rect 4154 2320 4160 2372
rect 4212 2320 4218 2372
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 5000 2360 5028 2388
rect 4571 2332 5028 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 5718 2320 5724 2372
rect 5776 2320 5782 2372
rect 7282 2320 7288 2372
rect 7340 2320 7346 2372
rect 9033 2363 9091 2369
rect 9033 2329 9045 2363
rect 9079 2329 9091 2363
rect 9140 2360 9168 2400
rect 9674 2388 9680 2440
rect 9732 2388 9738 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14507 2400 14596 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 10505 2363 10563 2369
rect 10505 2360 10517 2363
rect 9140 2332 10517 2360
rect 9033 2323 9091 2329
rect 10505 2329 10517 2332
rect 10551 2329 10563 2363
rect 10505 2323 10563 2329
rect 4890 2252 4896 2304
rect 4948 2252 4954 2304
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 9048 2292 9076 2323
rect 12066 2320 12072 2372
rect 12124 2320 12130 2372
rect 13538 2320 13544 2372
rect 13596 2320 13602 2372
rect 14568 2304 14596 2400
rect 8435 2264 9076 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 9122 2252 9128 2304
rect 9180 2252 9186 2304
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 11940 2264 12173 2292
rect 11940 2252 11946 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12161 2255 12219 2261
rect 13814 2252 13820 2304
rect 13872 2252 13878 2304
rect 14550 2252 14556 2304
rect 14608 2252 14614 2304
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 4890 2048 4896 2100
rect 4948 2048 4954 2100
rect 6546 2048 6552 2100
rect 6604 2088 6610 2100
rect 12066 2088 12072 2100
rect 6604 2060 12072 2088
rect 6604 2048 6610 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 13538 2048 13544 2100
rect 13596 2048 13602 2100
rect 4908 1952 4936 2048
rect 13556 1952 13584 2048
rect 4908 1924 13584 1952
<< via1 >>
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 2044 13472 2096 13524
rect 1308 13336 1360 13388
rect 1032 13268 1084 13320
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2044 13268 2096 13320
rect 2412 13268 2464 13320
rect 13728 13472 13780 13524
rect 4160 13268 4212 13320
rect 5172 13268 5224 13320
rect 6460 13336 6512 13388
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6736 13336 6788 13388
rect 7932 13268 7984 13320
rect 9312 13268 9364 13320
rect 10692 13268 10744 13320
rect 12072 13268 12124 13320
rect 13452 13268 13504 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4712 13132 4764 13184
rect 5724 13132 5776 13184
rect 5816 13132 5868 13184
rect 6092 13132 6144 13184
rect 6828 13175 6880 13184
rect 6828 13141 6837 13175
rect 6837 13141 6871 13175
rect 6871 13141 6880 13175
rect 6828 13132 6880 13141
rect 7656 13132 7708 13184
rect 9864 13132 9916 13184
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 1584 12928 1636 12980
rect 1860 12928 1912 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 3424 12928 3476 12980
rect 4160 12928 4212 12980
rect 5540 12928 5592 12980
rect 5632 12860 5684 12912
rect 6000 12903 6052 12912
rect 6000 12869 6009 12903
rect 6009 12869 6043 12903
rect 6043 12869 6052 12903
rect 6000 12860 6052 12869
rect 6736 12860 6788 12912
rect 13084 12928 13136 12980
rect 14464 12928 14516 12980
rect 14556 12928 14608 12980
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 3056 12724 3108 12776
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 3148 12588 3200 12640
rect 3240 12588 3292 12640
rect 4252 12656 4304 12708
rect 5816 12724 5868 12776
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 5632 12588 5684 12640
rect 12716 12588 12768 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 1676 12384 1728 12436
rect 2228 12384 2280 12436
rect 6000 12384 6052 12436
rect 6736 12384 6788 12436
rect 13360 12384 13412 12436
rect 2044 12248 2096 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3792 12316 3844 12368
rect 4804 12316 4856 12368
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 3148 12248 3200 12300
rect 4068 12248 4120 12300
rect 3516 12180 3568 12232
rect 3240 12155 3292 12164
rect 3240 12121 3249 12155
rect 3249 12121 3283 12155
rect 3283 12121 3292 12155
rect 3240 12112 3292 12121
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 12716 12248 12768 12300
rect 4896 12112 4948 12164
rect 5080 12155 5132 12164
rect 5080 12121 5114 12155
rect 5114 12121 5132 12155
rect 5080 12112 5132 12121
rect 13084 12180 13136 12232
rect 14004 12180 14056 12232
rect 14556 12180 14608 12232
rect 5540 12044 5592 12096
rect 7656 12044 7708 12096
rect 11888 12044 11940 12096
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 3148 11840 3200 11892
rect 3516 11840 3568 11892
rect 3792 11840 3844 11892
rect 4252 11840 4304 11892
rect 1676 11704 1728 11756
rect 4896 11840 4948 11892
rect 5080 11840 5132 11892
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 13360 11840 13412 11892
rect 10416 11815 10468 11824
rect 10416 11781 10425 11815
rect 10425 11781 10459 11815
rect 10459 11781 10468 11815
rect 10416 11772 10468 11781
rect 12808 11704 12860 11756
rect 13084 11704 13136 11756
rect 13912 11840 13964 11892
rect 7012 11636 7064 11688
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 8392 11611 8444 11620
rect 8392 11577 8401 11611
rect 8401 11577 8435 11611
rect 8435 11577 8444 11611
rect 8392 11568 8444 11577
rect 11612 11636 11664 11688
rect 13268 11636 13320 11688
rect 14188 11840 14240 11892
rect 2964 11500 3016 11552
rect 3424 11500 3476 11552
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 8116 11500 8168 11552
rect 12624 11543 12676 11552
rect 12624 11509 12633 11543
rect 12633 11509 12667 11543
rect 12667 11509 12676 11543
rect 12624 11500 12676 11509
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 2044 11296 2096 11348
rect 2964 11296 3016 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 5540 11296 5592 11348
rect 7012 11296 7064 11348
rect 8392 11296 8444 11348
rect 10416 11296 10468 11348
rect 2780 11160 2832 11169
rect 2964 11092 3016 11144
rect 3424 11228 3476 11280
rect 8116 11228 8168 11280
rect 7380 11160 7432 11212
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 11612 11296 11664 11348
rect 12624 11296 12676 11348
rect 13268 11296 13320 11348
rect 11888 11092 11940 11144
rect 12624 10956 12676 11008
rect 14556 11024 14608 11076
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 1768 10752 1820 10804
rect 2780 10752 2832 10804
rect 7656 10684 7708 10736
rect 12808 10684 12860 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 11612 10616 11664 10668
rect 12716 10616 12768 10668
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 940 10412 992 10464
rect 7564 10412 7616 10464
rect 14280 10480 14332 10532
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13452 10412 13504 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 1768 10208 1820 10260
rect 12440 10208 12492 10260
rect 7564 10140 7616 10192
rect 13452 10140 13504 10192
rect 3424 10072 3476 10124
rect 12624 10072 12676 10124
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 13820 10004 13872 10056
rect 12164 9979 12216 9988
rect 12164 9945 12173 9979
rect 12173 9945 12207 9979
rect 12207 9945 12216 9979
rect 12164 9936 12216 9945
rect 12808 9979 12860 9988
rect 12808 9945 12817 9979
rect 12817 9945 12851 9979
rect 12851 9945 12860 9979
rect 12808 9936 12860 9945
rect 13452 9979 13504 9988
rect 13452 9945 13461 9979
rect 13461 9945 13495 9979
rect 13495 9945 13504 9979
rect 13452 9936 13504 9945
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 14556 9868 14608 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 12164 9664 12216 9716
rect 12624 9664 12676 9716
rect 13452 9664 13504 9716
rect 13820 9664 13872 9716
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 13820 9528 13872 9580
rect 13912 9528 13964 9580
rect 12440 9460 12492 9512
rect 940 9324 992 9376
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 1768 8576 1820 8628
rect 2044 8440 2096 8492
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 14924 8304 14976 8356
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 14280 7352 14332 7404
rect 14280 7216 14332 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 14280 6987 14332 6996
rect 14280 6953 14289 6987
rect 14289 6953 14323 6987
rect 14323 6953 14332 6987
rect 14280 6944 14332 6953
rect 14924 6740 14976 6792
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 14188 6307 14240 6316
rect 14188 6273 14197 6307
rect 14197 6273 14231 6307
rect 14231 6273 14240 6307
rect 14188 6264 14240 6273
rect 940 6060 992 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 2136 5516 2188 5568
rect 14556 5516 14608 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 1768 5287 1820 5296
rect 1768 5253 1777 5287
rect 1777 5253 1811 5287
rect 1811 5253 1820 5287
rect 1768 5244 1820 5253
rect 940 4972 992 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 7380 4088 7432 4140
rect 14924 3952 14976 4004
rect 940 3884 992 3936
rect 13820 3884 13872 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 3700 3068 3752 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 6828 3000 6880 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 8852 2796 8904 2848
rect 15016 2796 15068 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 1768 2592 1820 2644
rect 14372 2592 14424 2644
rect 5908 2456 5960 2508
rect 12808 2524 12860 2576
rect 3056 2388 3108 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 4988 2388 5040 2440
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8852 2388 8904 2440
rect 2596 2363 2648 2372
rect 2596 2329 2605 2363
rect 2605 2329 2639 2363
rect 2639 2329 2648 2363
rect 2596 2320 2648 2329
rect 4160 2363 4212 2372
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 4160 2320 4212 2329
rect 5724 2363 5776 2372
rect 5724 2329 5733 2363
rect 5733 2329 5767 2363
rect 5767 2329 5776 2363
rect 5724 2320 5776 2329
rect 7288 2363 7340 2372
rect 7288 2329 7297 2363
rect 7297 2329 7331 2363
rect 7331 2329 7340 2363
rect 7288 2320 7340 2329
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 4896 2295 4948 2304
rect 4896 2261 4905 2295
rect 4905 2261 4939 2295
rect 4939 2261 4948 2295
rect 4896 2252 4948 2261
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 13544 2363 13596 2372
rect 13544 2329 13553 2363
rect 13553 2329 13587 2363
rect 13587 2329 13596 2363
rect 13544 2320 13596 2329
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 10324 2252 10376 2304
rect 11888 2252 11940 2304
rect 13820 2295 13872 2304
rect 13820 2261 13829 2295
rect 13829 2261 13863 2295
rect 13863 2261 13872 2295
rect 13820 2252 13872 2261
rect 14556 2252 14608 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 4896 2048 4948 2100
rect 6552 2048 6604 2100
rect 12072 2048 12124 2100
rect 13544 2048 13596 2100
<< metal2 >>
rect 1030 15200 1086 16000
rect 2410 15200 2466 16000
rect 3790 15314 3846 16000
rect 3790 15286 4108 15314
rect 3790 15200 3846 15286
rect 1044 13326 1072 15200
rect 1398 14376 1454 14385
rect 1398 14311 1454 14320
rect 1306 13424 1362 13433
rect 1306 13359 1308 13368
rect 1360 13359 1362 13368
rect 1308 13330 1360 13336
rect 1032 13320 1084 13326
rect 1032 13262 1084 13268
rect 1412 12238 1440 14311
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2056 13326 2084 13466
rect 2424 13326 2452 15200
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2412 13320 2464 13326
rect 4080 13308 4108 15286
rect 5170 15200 5226 16000
rect 6550 15200 6606 16000
rect 7930 15200 7986 16000
rect 9310 15200 9366 16000
rect 10690 15200 10746 16000
rect 12070 15200 12126 16000
rect 13450 15200 13506 16000
rect 14830 15314 14886 16000
rect 14476 15286 14886 15314
rect 5184 13326 5212 15200
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6564 13410 6592 15200
rect 6472 13394 6592 13410
rect 6460 13388 6592 13394
rect 6512 13382 6592 13388
rect 6736 13388 6788 13394
rect 6460 13330 6512 13336
rect 6736 13330 6788 13336
rect 4160 13320 4212 13326
rect 4080 13280 4160 13308
rect 2412 13262 2464 13268
rect 4160 13262 4212 13268
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12986 1624 13126
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1504 11665 1532 12582
rect 1688 12442 1716 13262
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12986 1900 13126
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11762 1716 12038
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1780 10810 1808 12786
rect 2056 12306 2084 13262
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 3252 12866 3280 13126
rect 3436 12986 3464 13126
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3252 12838 3740 12866
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2240 12442 2268 12718
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2056 11354 2084 12242
rect 2976 11558 3004 12242
rect 3068 12186 3096 12718
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3160 12306 3188 12582
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3068 12158 3188 12186
rect 3252 12170 3280 12582
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3160 11898 3188 12158
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3528 11898 3556 12174
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2964 11348 3016 11354
rect 3068 11336 3096 11630
rect 3016 11308 3096 11336
rect 2964 11290 3016 11296
rect 3160 11234 3188 11834
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 11286 3464 11494
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2976 11206 3188 11234
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 2792 10810 2820 11154
rect 2976 11150 3004 11206
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10169 980 10406
rect 1780 10266 1808 10610
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 938 10160 994 10169
rect 3436 10130 3464 11222
rect 938 10095 994 10104
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 952 9081 980 9318
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1596 6914 1624 9862
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 8634 1808 9522
rect 2976 9466 3004 9862
rect 2976 9438 3096 9466
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2056 7546 2084 8434
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1490 6896 1546 6905
rect 1596 6886 1808 6914
rect 1490 6831 1546 6840
rect 940 6112 992 6118
rect 940 6054 992 6060
rect 952 5817 980 6054
rect 938 5808 994 5817
rect 938 5743 994 5752
rect 1780 5302 1808 6886
rect 2148 5574 2176 8434
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4729 980 4966
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 3641 980 3878
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2689 1532 2790
rect 1490 2680 1546 2689
rect 1780 2650 1808 2994
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 1490 2615 1546 2624
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 3068 2446 3096 9438
rect 3712 3126 3740 12838
rect 3804 12374 3832 13126
rect 4172 12986 4200 13126
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 4066 12336 4122 12345
rect 4066 12271 4068 12280
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11898 3832 12038
rect 4264 11898 4292 12650
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 4724 2446 4752 13126
rect 5552 12986 5580 13262
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5644 12646 5672 12854
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 12458 5672 12582
rect 5552 12430 5672 12458
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4816 2774 4844 12310
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4908 11898 4936 12106
rect 5092 11898 5120 12106
rect 5552 12102 5580 12430
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5736 2774 5764 13126
rect 5828 12782 5856 13126
rect 6104 13002 6132 13126
rect 5920 12974 6132 13002
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5920 7562 5948 12974
rect 6748 12918 6776 13330
rect 7944 13326 7972 15200
rect 9324 13326 9352 15200
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 10704 13326 10732 15200
rect 12084 13326 12112 15200
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 13464 13326 13492 15200
rect 13726 14784 13782 14793
rect 13726 14719 13782 14728
rect 13740 13530 13768 14719
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6012 12442 6040 12854
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6748 12442 6776 12854
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 5920 7534 6040 7562
rect 4816 2746 5028 2774
rect 5736 2746 5948 2774
rect 5000 2446 5028 2746
rect 5920 2514 5948 2746
rect 6012 2530 6040 7534
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6840 3058 6868 13126
rect 7668 12434 7696 13126
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 7668 12406 8248 12434
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 11354 7052 11630
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 4146 7420 11154
rect 7668 10742 7696 12038
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7944 11218 7972 11630
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11286 8156 11494
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 10198 7604 10406
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 5908 2508 5960 2514
rect 6012 2502 6132 2530
rect 5908 2450 5960 2456
rect 6104 2446 6132 2502
rect 8220 2446 8248 12406
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 11354 8432 11562
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8864 2446 8892 2790
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 9876 2530 9904 13126
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 13096 12986 13124 13126
rect 14476 12986 14504 15286
rect 14830 15200 14886 15286
rect 14646 13424 14702 13433
rect 14568 13382 14646 13410
rect 14568 12986 14596 13382
rect 14646 13359 14702 13368
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 11532 12434 11560 12718
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 11532 12406 11652 12434
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10428 11354 10456 11766
rect 11624 11694 11652 12406
rect 12728 12306 12756 12582
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 13372 12442 13400 12718
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11624 11354 11652 11630
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11624 10674 11652 11290
rect 11900 11150 11928 12038
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 11354 12664 11494
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 12176 9722 12204 9930
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12452 9518 12480 10202
rect 12636 10130 12664 10950
rect 12728 10674 12756 12242
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11762 13124 12174
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11898 13400 12038
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12820 11234 12848 11698
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 13280 11354 13308 11630
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12820 11206 12940 11234
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10742 12848 10950
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12912 10470 12940 11206
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13464 10198 13492 10406
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12636 9722 12664 10066
rect 13832 10062 13860 12582
rect 14016 12238 14044 12582
rect 14004 12232 14056 12238
rect 14556 12232 14608 12238
rect 14004 12174 14056 12180
rect 14554 12200 14556 12209
rect 14608 12200 14610 12209
rect 14554 12135 14610 12144
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 13924 11898 13952 12038
rect 14200 11898 14228 12038
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 12820 2582 12848 9930
rect 13464 9722 13492 9930
rect 13832 9722 13860 9998
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 9586 13952 9862
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 13832 3942 13860 9522
rect 14200 9194 14228 10610
rect 14292 10538 14320 10950
rect 14568 10713 14596 11018
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14554 10704 14610 10713
rect 14554 10639 14610 10648
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 13924 9166 14228 9194
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 13924 3194 13952 9166
rect 14292 9058 14320 9862
rect 14568 9353 14596 9862
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14554 9344 14610 9353
rect 14554 9279 14610 9288
rect 14200 9030 14320 9058
rect 14200 6322 14228 9030
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8378 14320 8910
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14292 8350 14412 8378
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7410 14320 8230
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 7002 14320 7210
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 9692 2502 9904 2530
rect 12808 2576 12860 2582
rect 13740 2553 13768 2994
rect 14384 2650 14412 8350
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7993 14964 8298
rect 14922 7984 14978 7993
rect 14922 7919 14978 7928
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14924 6792 14976 6798
rect 14922 6760 14924 6769
rect 14976 6760 14978 6769
rect 14922 6695 14978 6704
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5273 14596 5510
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14554 5264 14610 5273
rect 14554 5199 14610 5208
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14936 3913 14964 3946
rect 14922 3904 14978 3913
rect 14922 3839 14978 3848
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 12808 2518 12860 2524
rect 13726 2544 13782 2553
rect 9692 2446 9720 2502
rect 13726 2479 13782 2488
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 2596 2372 2648 2378
rect 2516 2332 2596 2360
rect 2516 800 2544 2332
rect 4160 2372 4212 2378
rect 2596 2314 2648 2320
rect 4080 2332 4160 2360
rect 4080 800 4108 2332
rect 5724 2372 5776 2378
rect 4160 2314 4212 2320
rect 5644 2332 5724 2360
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 4908 2106 4936 2246
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5644 800 5672 2332
rect 5724 2314 5776 2320
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 2106 6592 2246
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 7300 1170 7328 2314
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 7208 1142 7328 1170
rect 7208 800 7236 1142
rect 8772 870 8892 898
rect 8772 800 8800 870
rect 2502 0 2558 800
rect 4066 0 4122 800
rect 5630 0 5686 800
rect 7194 0 7250 800
rect 8758 0 8814 800
rect 8864 762 8892 870
rect 9140 762 9168 2246
rect 10336 800 10364 2246
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 11900 800 11928 2246
rect 12084 2106 12112 2314
rect 13556 2106 13584 2314
rect 13820 2304 13872 2310
rect 13740 2264 13820 2292
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13464 870 13584 898
rect 13464 800 13492 870
rect 8864 734 9168 762
rect 10322 0 10378 800
rect 11886 0 11942 800
rect 13450 0 13506 800
rect 13556 762 13584 870
rect 13740 762 13768 2264
rect 13820 2246 13872 2252
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14568 1193 14596 2246
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 14554 1184 14610 1193
rect 14554 1119 14610 1128
rect 15028 800 15056 2790
rect 13556 734 13768 762
rect 15014 0 15070 800
<< via2 >>
rect 1398 14320 1454 14376
rect 1306 13388 1362 13424
rect 1306 13368 1308 13388
rect 1308 13368 1360 13388
rect 1360 13368 1362 13388
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 1490 11600 1546 11656
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 938 10104 994 10160
rect 938 9016 994 9072
rect 1490 8200 1546 8256
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 1490 6840 1546 6896
rect 938 5752 994 5808
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 938 4664 994 4720
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 938 3576 994 3632
rect 1490 2624 1546 2680
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 13726 14728 13782 14784
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 14646 13368 14702 13424
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 14554 12180 14556 12200
rect 14556 12180 14608 12200
rect 14608 12180 14610 12200
rect 14554 12144 14610 12180
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14554 10648 14610 10704
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14554 9288 14610 9344
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14922 7928 14978 7984
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14922 6740 14924 6760
rect 14924 6740 14976 6760
rect 14976 6740 14978 6760
rect 14922 6704 14978 6740
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14554 5208 14610 5264
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14922 3848 14978 3904
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 13726 2488 13782 2544
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 14554 1128 14610 1184
<< metal3 >>
rect 13721 14786 13787 14789
rect 15200 14786 16000 14816
rect 13721 14784 16000 14786
rect 13721 14728 13726 14784
rect 13782 14728 16000 14784
rect 13721 14726 16000 14728
rect 13721 14723 13787 14726
rect 15200 14696 16000 14726
rect 0 14514 800 14544
rect 0 14454 1042 14514
rect 0 14424 800 14454
rect 982 14378 1042 14454
rect 1393 14378 1459 14381
rect 982 14376 1459 14378
rect 982 14320 1398 14376
rect 1454 14320 1459 14376
rect 982 14318 1459 14320
rect 1393 14315 1459 14318
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 0 13426 800 13456
rect 1301 13426 1367 13429
rect 0 13424 1367 13426
rect 0 13368 1306 13424
rect 1362 13368 1367 13424
rect 0 13366 1367 13368
rect 0 13336 800 13366
rect 1301 13363 1367 13366
rect 14641 13426 14707 13429
rect 15200 13426 16000 13456
rect 14641 13424 16000 13426
rect 14641 13368 14646 13424
rect 14702 13368 16000 13424
rect 14641 13366 16000 13368
rect 14641 13363 14707 13366
rect 15200 13336 16000 13366
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 14549 12202 14615 12205
rect 14549 12200 15210 12202
rect 14549 12144 14554 12200
rect 14610 12144 15210 12200
rect 14549 12142 15210 12144
rect 14549 12139 14615 12142
rect 15150 12096 15210 12142
rect 15150 12006 16000 12096
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 15200 11976 16000 12006
rect 14653 11935 14969 11936
rect 1485 11656 1551 11661
rect 1485 11600 1490 11656
rect 1546 11600 1551 11656
rect 1485 11595 1551 11600
rect 0 11250 800 11280
rect 1488 11250 1548 11595
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 0 11190 1548 11250
rect 0 11160 800 11190
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 14549 10706 14615 10709
rect 15200 10706 16000 10736
rect 14549 10704 16000 10706
rect 14549 10648 14554 10704
rect 14610 10648 16000 10704
rect 14549 10646 16000 10648
rect 14549 10643 14615 10646
rect 15200 10616 16000 10646
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 14549 9346 14615 9349
rect 15200 9346 16000 9376
rect 14549 9344 16000 9346
rect 14549 9288 14554 9344
rect 14610 9288 16000 9344
rect 14549 9286 16000 9288
rect 14549 9283 14615 9286
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 15200 9256 16000 9286
rect 12940 9215 13256 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 1485 8256 1551 8261
rect 1485 8200 1490 8256
rect 1546 8200 1551 8256
rect 1485 8195 1551 8200
rect 0 7986 800 8016
rect 1488 7986 1548 8195
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 0 7926 1548 7986
rect 14917 7986 14983 7989
rect 15200 7986 16000 8016
rect 14917 7984 16000 7986
rect 14917 7928 14922 7984
rect 14978 7928 16000 7984
rect 14917 7926 16000 7928
rect 0 7896 800 7926
rect 14917 7923 14983 7926
rect 15200 7896 16000 7926
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 12940 7039 13256 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 14917 6762 14983 6765
rect 14917 6760 15210 6762
rect 14917 6704 14922 6760
rect 14978 6704 15210 6760
rect 14917 6702 15210 6704
rect 14917 6699 14983 6702
rect 15150 6656 15210 6702
rect 15150 6566 16000 6656
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 15200 6536 16000 6566
rect 14653 6495 14969 6496
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 14549 5266 14615 5269
rect 15200 5266 16000 5296
rect 14549 5264 16000 5266
rect 14549 5208 14554 5264
rect 14610 5208 16000 5264
rect 14549 5206 16000 5208
rect 14549 5203 14615 5206
rect 15200 5176 16000 5206
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 14917 3906 14983 3909
rect 15200 3906 16000 3936
rect 14917 3904 16000 3906
rect 14917 3848 14922 3904
rect 14978 3848 16000 3904
rect 14917 3846 16000 3848
rect 14917 3843 14983 3846
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 15200 3816 16000 3846
rect 12940 3775 13256 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 1485 2682 1551 2685
rect 798 2680 1551 2682
rect 798 2624 1490 2680
rect 1546 2624 1551 2680
rect 798 2622 1551 2624
rect 798 2576 858 2622
rect 1485 2619 1551 2622
rect 0 2486 858 2576
rect 13721 2546 13787 2549
rect 15200 2546 16000 2576
rect 13721 2544 16000 2546
rect 13721 2488 13726 2544
rect 13782 2488 16000 2544
rect 13721 2486 16000 2488
rect 0 2456 800 2486
rect 13721 2483 13787 2486
rect 15200 2456 16000 2486
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 14549 1186 14615 1189
rect 15200 1186 16000 1216
rect 14549 1184 16000 1186
rect 14549 1128 14554 1184
rect 14610 1128 16000 1184
rect 14549 1126 16000 1128
rect 14549 1123 14615 1126
rect 15200 1096 16000 1126
<< via3 >>
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 13632 2977 13648
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 13088 4690 13648
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 13632 6404 13648
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 13088 8117 13648
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 13632 9831 13648
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 13088 11544 13648
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 13632 13258 13648
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 13088 14971 13648
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__inv_2  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform -1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform -1 0 4140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform -1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp 1688980957
transform -1 0 3772 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 1688980957
transform 1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform -1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform -1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _039_
timestamp 1688980957
transform 1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform -1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform -1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform -1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform -1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform -1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp 1688980957
transform 1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform -1 0 13984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform -1 0 13248 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp 1688980957
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 1688980957
transform -1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1688980957
transform 1 0 14168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform 1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1688980957
transform -1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1688980957
transform -1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1688980957
transform -1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform -1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _065_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _066_
timestamp 1688980957
transform -1 0 9844 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _067_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _068_
timestamp 1688980957
transform 1 0 1564 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _069_
timestamp 1688980957
transform -1 0 2852 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _070_
timestamp 1688980957
transform 1 0 4784 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _071_
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform -1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp 1688980957
transform -1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp 1688980957
transform -1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _084_
timestamp 1688980957
transform -1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _088_
timestamp 1688980957
transform -1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _090_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _091_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13708 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _092_
timestamp 1688980957
transform -1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _093_
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _093__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _094__44
timestamp 1688980957
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _094_
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _095_
timestamp 1688980957
transform -1 0 13432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _096_
timestamp 1688980957
transform -1 0 14168 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _097_
timestamp 1688980957
transform -1 0 10672 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _098__45
timestamp 1688980957
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _098_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _099_
timestamp 1688980957
transform 1 0 2024 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _100_
timestamp 1688980957
transform -1 0 3496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _101_
timestamp 1688980957
transform -1 0 3496 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _102_
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _103__46
timestamp 1688980957
transform 1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _103_
timestamp 1688980957
transform -1 0 7728 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _104_
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _105_
timestamp 1688980957
transform 1 0 5336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_42
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_66 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_73
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_80
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_94
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_107
timestamp 1688980957
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_124
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_132
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_33
timestamp 1688980957
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_45
timestamp 1688980957
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_66
timestamp 1688980957
transform 1 0 7176 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_78
timestamp 1688980957
transform 1 0 8280 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_145
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_12
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_24
timestamp 1688980957
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_36
timestamp 1688980957
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_145
timestamp 1688980957
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_21
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_45
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1688980957
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_143
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_16
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_28
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_40
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_145
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_36
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_48
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_144
timestamp 1688980957
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_130
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_8
timestamp 1688980957
transform 1 0 1840 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_16
timestamp 1688980957
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_22
timestamp 1688980957
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_132
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_143
timestamp 1688980957
transform 1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_38
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_62
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_68
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_106
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_110
timestamp 1688980957
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_37
timestamp 1688980957
transform 1 0 4508 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_73
timestamp 1688980957
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_77
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_104
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_145
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1688980957
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_59
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 1688980957
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_144
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_29
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_75
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_87
timestamp 1688980957
transform 1 0 9108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_129
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_139
timestamp 1688980957
transform 1 0 13892 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_10
timestamp 1688980957
transform 1 0 2024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_14
timestamp 1688980957
transform 1 0 2392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_38
timestamp 1688980957
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_54
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_63
timestamp 1688980957
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 1688980957
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_108
timestamp 1688980957
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_113
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_119
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_123
timestamp 1688980957
transform 1 0 12420 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_144
timestamp 1688980957
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 4784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 2392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 13524 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 6256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 14260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform -1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform -1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform -1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 13984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 12420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 4692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 11960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform -1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
<< labels >>
flabel metal3 s 15200 13336 16000 13456 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 15200 14696 16000 14816 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 15200 1096 16000 1216 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 15200 2456 16000 2576 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 3 nsew signal input
flabel metal3 s 15200 3816 16000 3936 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 4 nsew signal input
flabel metal3 s 15200 5176 16000 5296 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 5 nsew signal input
flabel metal3 s 15200 6536 16000 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 6 nsew signal input
flabel metal3 s 15200 7896 16000 8016 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 7 nsew signal input
flabel metal3 s 15200 9256 16000 9376 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 8 nsew signal input
flabel metal3 s 15200 10616 16000 10736 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 9 nsew signal input
flabel metal3 s 15200 11976 16000 12096 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 10 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 11 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 12 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 13 nsew signal tristate
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 14 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 15 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 16 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 17 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 18 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 19 nsew signal tristate
flabel metal2 s 1030 15200 1086 16000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 20 nsew signal input
flabel metal2 s 2410 15200 2466 16000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 21 nsew signal input
flabel metal2 s 3790 15200 3846 16000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 22 nsew signal input
flabel metal2 s 5170 15200 5226 16000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 23 nsew signal input
flabel metal2 s 6550 15200 6606 16000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 24 nsew signal input
flabel metal2 s 7930 15200 7986 16000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 25 nsew signal input
flabel metal2 s 9310 15200 9366 16000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 26 nsew signal input
flabel metal2 s 10690 15200 10746 16000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 27 nsew signal input
flabel metal2 s 12070 15200 12126 16000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 28 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chany_top_out[0]
port 29 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chany_top_out[1]
port 30 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chany_top_out[2]
port 31 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chany_top_out[3]
port 32 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_out[4]
port 33 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chany_top_out[5]
port 34 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chany_top_out[6]
port 35 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chany_top_out[7]
port 36 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chany_top_out[8]
port 37 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 38 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 39 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 prog_clk
port 40 nsew signal input
flabel metal2 s 13450 15200 13506 16000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 41 nsew signal input
flabel metal2 s 14830 15200 14886 16000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 42 nsew signal input
flabel metal4 s 2657 2128 2977 13648 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 6084 2128 6404 13648 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 9511 2128 9831 13648 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 12938 2128 13258 13648 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 4370 2128 4690 13648 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 13648 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 13648 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 13648 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 7958 13600 7958 13600 0 vdd
rlabel via1 8037 13056 8037 13056 0 vss
rlabel metal1 6624 12818 6624 12818 0 _000_
rlabel metal1 4140 12818 4140 12818 0 _001_
rlabel metal1 2622 12274 2622 12274 0 _002_
rlabel metal1 3174 11186 3174 11186 0 _003_
rlabel metal1 13754 11152 13754 11152 0 _004_
rlabel metal1 7452 11118 7452 11118 0 _005_
rlabel metal1 11776 10030 11776 10030 0 _006_
rlabel metal1 13754 10064 13754 10064 0 _007_
rlabel metal1 13248 12410 13248 12410 0 _008_
rlabel metal1 13202 9690 13202 9690 0 _009_
rlabel metal1 14076 9554 14076 9554 0 _010_
rlabel metal1 12282 9928 12282 9928 0 _011_
rlabel metal1 7912 11050 7912 11050 0 _012_
rlabel metal1 13432 11322 13432 11322 0 _013_
rlabel metal1 13800 11730 13800 11730 0 _014_
rlabel metal1 10028 11322 10028 11322 0 _015_
rlabel metal1 4002 11016 4002 11016 0 _016_
rlabel metal1 2346 12410 2346 12410 0 _017_
rlabel metal2 1886 13056 1886 13056 0 _018_
rlabel metal1 3450 12614 3450 12614 0 _019_
rlabel metal1 4922 12716 4922 12716 0 _020_
rlabel metal1 7176 12886 7176 12886 0 _021_
rlabel metal1 6210 12410 6210 12410 0 _022_
rlabel metal1 5060 12954 5060 12954 0 _023_
rlabel metal1 14536 12818 14536 12818 0 ccff_head
rlabel metal1 13800 13498 13800 13498 0 ccff_tail
rlabel metal1 14536 2414 14536 2414 0 chanx_left_in[0]
rlabel metal2 13754 2771 13754 2771 0 chanx_left_in[1]
rlabel metal1 14720 4114 14720 4114 0 chanx_left_in[2]
rlabel metal1 14536 5678 14536 5678 0 chanx_left_in[3]
rlabel metal1 14720 6766 14720 6766 0 chanx_left_in[4]
rlabel metal1 14720 8466 14720 8466 0 chanx_left_in[5]
rlabel metal1 14536 10030 14536 10030 0 chanx_left_in[6]
rlabel metal1 14536 11118 14536 11118 0 chanx_left_in[7]
rlabel metal1 13754 12240 13754 12240 0 chanx_left_in[8]
rlabel metal2 2530 1554 2530 1554 0 chanx_left_out[0]
rlabel metal2 4094 1554 4094 1554 0 chanx_left_out[1]
rlabel metal2 5658 1554 5658 1554 0 chanx_left_out[2]
rlabel metal2 7222 959 7222 959 0 chanx_left_out[3]
rlabel metal2 8786 823 8786 823 0 chanx_left_out[4]
rlabel metal2 10350 1520 10350 1520 0 chanx_left_out[5]
rlabel metal2 11914 1520 11914 1520 0 chanx_left_out[6]
rlabel metal2 13478 823 13478 823 0 chanx_left_out[7]
rlabel metal2 15042 1792 15042 1792 0 chanx_left_out[8]
rlabel metal1 2162 13260 2162 13260 0 chany_top_in[0]
rlabel metal1 2484 13294 2484 13294 0 chany_top_in[1]
rlabel metal1 4278 13294 4278 13294 0 chany_top_in[2]
rlabel metal1 5014 13294 5014 13294 0 chany_top_in[3]
rlabel metal1 6670 13328 6670 13328 0 chany_top_in[4]
rlabel metal1 8004 13294 8004 13294 0 chany_top_in[5]
rlabel metal1 9384 13294 9384 13294 0 chany_top_in[6]
rlabel metal1 10856 13294 10856 13294 0 chany_top_in[7]
rlabel metal1 12236 13294 12236 13294 0 chany_top_in[8]
rlabel metal3 751 2516 751 2516 0 chany_top_out[0]
rlabel metal3 820 3604 820 3604 0 chany_top_out[1]
rlabel metal3 820 4692 820 4692 0 chany_top_out[2]
rlabel metal3 820 5780 820 5780 0 chany_top_out[3]
rlabel metal3 1096 6868 1096 6868 0 chany_top_out[4]
rlabel metal3 1096 7956 1096 7956 0 chany_top_out[5]
rlabel metal3 820 9044 820 9044 0 chany_top_out[6]
rlabel metal3 820 10132 820 10132 0 chany_top_out[7]
rlabel metal3 1096 11220 1096 11220 0 chany_top_out[8]
rlabel metal1 6118 10710 6118 10710 0 clknet_0_prog_clk
rlabel metal1 1610 11764 1610 11764 0 clknet_1_0__leaf_prog_clk
rlabel metal2 11546 12585 11546 12585 0 clknet_1_1__leaf_prog_clk
rlabel metal3 1004 13396 1004 13396 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 843 14484 843 14484 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 7084 11118 7084 11118 0 mem_left_track_1.DFF_0_.D
rlabel metal1 1932 13294 1932 13294 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 3404 12750 3404 12750 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 4370 12818 4370 12818 0 mem_left_track_3.DFF_0_.Q
rlabel metal1 12834 12274 12834 12274 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 12742 11016 12742 11016 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 12788 11730 12788 11730 0 mem_top_track_2.DFF_0_.Q
rlabel metal1 3450 12886 3450 12886 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 2070 12852 2070 12852 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 2990 12614 2990 12614 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3956 11254 3956 11254 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5290 13362 5290 13362 0 mux_left_track_3.INVTX1_0_.out
rlabel metal1 4738 12852 4738 12852 0 mux_left_track_3.INVTX1_1_.out
rlabel metal1 5750 12750 5750 12750 0 mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 5612 12444 5612 12444 0 mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13156 12818 13156 12818 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 14536 9146 14536 9146 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 13708 9962 13708 9962 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 1794 2482 1794 2482 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 14122 11764 14122 11764 0 mux_top_track_2.INVTX1_0_.out
rlabel metal1 13386 11628 13386 11628 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 13110 11798 13110 11798 0 mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 8326 11220 8326 11220 0 mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13018 12750 13018 12750 0 net1
rlabel metal1 14214 11696 14214 11696 0 net10
rlabel metal1 3358 13362 3358 13362 0 net11
rlabel metal1 2714 13192 2714 13192 0 net12
rlabel metal1 4646 13158 4646 13158 0 net13
rlabel metal1 6164 2482 6164 2482 0 net14
rlabel metal1 6900 3026 6900 3026 0 net15
rlabel metal1 7958 13158 7958 13158 0 net16
rlabel metal2 9798 2516 9798 2516 0 net17
rlabel viali 6573 13294 6573 13294 0 net18
rlabel metal1 5382 13294 5382 13294 0 net19
rlabel metal1 14352 2618 14352 2618 0 net2
rlabel metal1 4094 13260 4094 13260 0 net20
rlabel metal1 1656 12410 1656 12410 0 net21
rlabel metal1 13202 13328 13202 13328 0 net22
rlabel metal1 14076 12206 14076 12206 0 net23
rlabel metal1 11086 13294 11086 13294 0 net24
rlabel metal1 3036 2414 3036 2414 0 net25
rlabel metal1 4784 2346 4784 2346 0 net26
rlabel metal2 6072 2516 6072 2516 0 net27
rlabel metal1 7682 2448 7682 2448 0 net28
rlabel metal1 9062 2312 9062 2312 0 net29
rlabel metal2 14076 9180 14076 9180 0 net3
rlabel metal1 9844 2346 9844 2346 0 net30
rlabel metal2 6578 2176 6578 2176 0 net31
rlabel metal1 4922 2006 4922 2006 0 net32
rlabel metal2 3496 12852 3496 12852 0 net33
rlabel metal1 1748 2618 1748 2618 0 net34
rlabel metal1 1932 4114 1932 4114 0 net35
rlabel metal2 1794 6085 1794 6085 0 net36
rlabel metal1 2277 6290 2277 6290 0 net37
rlabel metal1 2070 7446 2070 7446 0 net38
rlabel metal2 2070 7990 2070 7990 0 net39
rlabel metal1 14076 3910 14076 3910 0 net4
rlabel metal1 1886 8602 1886 8602 0 net40
rlabel metal2 1794 10438 1794 10438 0 net41
rlabel metal1 1794 10744 1794 10744 0 net42
rlabel metal1 12236 9690 12236 9690 0 net43
rlabel metal2 7958 11424 7958 11424 0 net44
rlabel metal1 3772 11050 3772 11050 0 net45
rlabel metal1 7682 12750 7682 12750 0 net46
rlabel metal1 3583 11798 3583 11798 0 net47
rlabel metal1 5290 11866 5290 11866 0 net48
rlabel metal1 1784 11730 1784 11730 0 net49
rlabel metal2 2162 7004 2162 7004 0 net5
rlabel metal2 12834 10846 12834 10846 0 net50
rlabel metal1 11771 11118 11771 11118 0 net51
rlabel metal1 3542 11118 3542 11118 0 net52
rlabel metal1 9951 11798 9951 11798 0 net53
rlabel metal1 2254 7310 2254 7310 0 net6
rlabel metal2 14306 7820 14306 7820 0 net7
rlabel metal2 14260 9044 14260 9044 0 net8
rlabel metal1 1794 10064 1794 10064 0 net9
rlabel via2 4094 12291 4094 12291 0 prog_clk
rlabel metal1 13892 13294 13892 13294 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 14214 12852 14214 12852 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
