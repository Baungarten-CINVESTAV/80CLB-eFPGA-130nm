VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_1__1_
  CLASS BLOCK ;
  FOREIGN cby_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 60.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 49.000 60.000 49.600 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 53.080 60.000 53.680 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.770 56.000 4.050 60.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 10.210 56.000 10.490 60.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.650 56.000 16.930 60.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 56.000 23.370 60.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.530 56.000 29.810 60.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 56.000 36.250 60.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 56.000 42.690 60.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 56.000 49.130 60.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 55.290 56.000 55.570 60.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 4.120 60.000 4.720 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 8.200 60.000 8.800 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 12.280 60.000 12.880 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 16.360 60.000 16.960 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 20.440 60.000 21.040 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 24.520 60.000 25.120 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 28.600 60.000 29.200 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 32.680 60.000 33.280 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 36.760 60.000 37.360 ;
    END
  END chany_top_out[8]
  PIN left_grid_right_width_0_height_0_subtile_0__pin_I_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END left_grid_right_width_0_height_0_subtile_0__pin_I_1_
  PIN left_grid_right_width_0_height_0_subtile_0__pin_I_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END left_grid_right_width_0_height_0_subtile_0__pin_I_5_
  PIN left_grid_right_width_0_height_0_subtile_0__pin_I_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END left_grid_right_width_0_height_0_subtile_0__pin_I_9_
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END prog_clk
  PIN right_grid_left_width_0_height_0_subtile_0__pin_I_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 56.000 40.840 60.000 41.440 ;
    END
  END right_grid_left_width_0_height_0_subtile_0__pin_I_3_
  PIN right_grid_left_width_0_height_0_subtile_0__pin_I_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 56.000 44.920 60.000 45.520 ;
    END
  END right_grid_left_width_0_height_0_subtile_0__pin_I_7_
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 49.200 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.910 10.640 18.510 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.100 10.640 30.700 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.290 10.640 42.890 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.480 10.640 55.080 49.200 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 49.045 ;
      LAYER met1 ;
        RECT 2.830 6.840 55.590 49.200 ;
      LAYER met2 ;
        RECT 2.860 55.720 3.490 56.285 ;
        RECT 4.330 55.720 9.930 56.285 ;
        RECT 10.770 55.720 16.370 56.285 ;
        RECT 17.210 55.720 22.810 56.285 ;
        RECT 23.650 55.720 29.250 56.285 ;
        RECT 30.090 55.720 35.690 56.285 ;
        RECT 36.530 55.720 42.130 56.285 ;
        RECT 42.970 55.720 48.570 56.285 ;
        RECT 49.410 55.720 55.010 56.285 ;
        RECT 2.860 4.280 55.560 55.720 ;
        RECT 3.410 4.000 8.550 4.280 ;
        RECT 9.390 4.000 14.530 4.280 ;
        RECT 15.370 4.000 20.510 4.280 ;
        RECT 21.350 4.000 26.490 4.280 ;
        RECT 27.330 4.000 32.470 4.280 ;
        RECT 33.310 4.000 38.450 4.280 ;
        RECT 39.290 4.000 44.430 4.280 ;
        RECT 45.270 4.000 50.410 4.280 ;
        RECT 51.250 4.000 55.560 4.280 ;
      LAYER met3 ;
        RECT 4.400 55.400 57.650 56.265 ;
        RECT 3.990 54.080 57.650 55.400 ;
        RECT 3.990 52.720 55.600 54.080 ;
        RECT 4.400 52.680 55.600 52.720 ;
        RECT 4.400 51.320 57.650 52.680 ;
        RECT 3.990 50.000 57.650 51.320 ;
        RECT 3.990 48.640 55.600 50.000 ;
        RECT 4.400 48.600 55.600 48.640 ;
        RECT 4.400 47.240 57.650 48.600 ;
        RECT 3.990 45.920 57.650 47.240 ;
        RECT 3.990 44.560 55.600 45.920 ;
        RECT 4.400 44.520 55.600 44.560 ;
        RECT 4.400 43.160 57.650 44.520 ;
        RECT 3.990 41.840 57.650 43.160 ;
        RECT 3.990 40.480 55.600 41.840 ;
        RECT 4.400 40.440 55.600 40.480 ;
        RECT 4.400 39.080 57.650 40.440 ;
        RECT 3.990 37.760 57.650 39.080 ;
        RECT 3.990 36.400 55.600 37.760 ;
        RECT 4.400 36.360 55.600 36.400 ;
        RECT 4.400 35.000 57.650 36.360 ;
        RECT 3.990 33.680 57.650 35.000 ;
        RECT 3.990 32.320 55.600 33.680 ;
        RECT 4.400 32.280 55.600 32.320 ;
        RECT 4.400 30.920 57.650 32.280 ;
        RECT 3.990 29.600 57.650 30.920 ;
        RECT 3.990 28.240 55.600 29.600 ;
        RECT 4.400 28.200 55.600 28.240 ;
        RECT 4.400 26.840 57.650 28.200 ;
        RECT 3.990 25.520 57.650 26.840 ;
        RECT 3.990 24.160 55.600 25.520 ;
        RECT 4.400 24.120 55.600 24.160 ;
        RECT 4.400 22.760 57.650 24.120 ;
        RECT 3.990 21.440 57.650 22.760 ;
        RECT 3.990 20.080 55.600 21.440 ;
        RECT 4.400 20.040 55.600 20.080 ;
        RECT 4.400 18.680 57.650 20.040 ;
        RECT 3.990 17.360 57.650 18.680 ;
        RECT 3.990 16.000 55.600 17.360 ;
        RECT 4.400 15.960 55.600 16.000 ;
        RECT 4.400 14.600 57.650 15.960 ;
        RECT 3.990 13.280 57.650 14.600 ;
        RECT 3.990 11.920 55.600 13.280 ;
        RECT 4.400 11.880 55.600 11.920 ;
        RECT 4.400 10.520 57.650 11.880 ;
        RECT 3.990 9.200 57.650 10.520 ;
        RECT 3.990 7.840 55.600 9.200 ;
        RECT 4.400 7.800 55.600 7.840 ;
        RECT 4.400 6.440 57.650 7.800 ;
        RECT 3.990 5.120 57.650 6.440 ;
        RECT 3.990 4.255 55.600 5.120 ;
  END
END cby_1__1_
END LIBRARY

