magic
tech sky130A
magscale 1 2
timestamp 1710357839
<< viali >>
rect 4537 13277 4571 13311
rect 1409 13209 1443 13243
rect 1777 13209 1811 13243
rect 4353 13141 4387 13175
rect 2881 12937 2915 12971
rect 3065 12801 3099 12835
rect 4537 10217 4571 10251
rect 3157 6273 3191 6307
rect 3424 6273 3458 6307
rect 4537 6069 4571 6103
rect 4353 5865 4387 5899
rect 4537 5661 4571 5695
rect 4353 2601 4387 2635
rect 4537 2397 4571 2431
<< metal1 >>
rect 1104 13626 4876 13648
rect 1104 13574 1421 13626
rect 1473 13574 1485 13626
rect 1537 13574 1549 13626
rect 1601 13574 1613 13626
rect 1665 13574 1677 13626
rect 1729 13574 2364 13626
rect 2416 13574 2428 13626
rect 2480 13574 2492 13626
rect 2544 13574 2556 13626
rect 2608 13574 2620 13626
rect 2672 13574 3307 13626
rect 3359 13574 3371 13626
rect 3423 13574 3435 13626
rect 3487 13574 3499 13626
rect 3551 13574 3563 13626
rect 3615 13574 4250 13626
rect 4302 13574 4314 13626
rect 4366 13574 4378 13626
rect 4430 13574 4442 13626
rect 4494 13574 4506 13626
rect 4558 13574 4876 13626
rect 1104 13552 4876 13574
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13308 4583 13311
rect 4890 13308 4896 13320
rect 4571 13280 4896 13308
rect 4571 13277 4583 13280
rect 4525 13271 4583 13277
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 1394 13200 1400 13252
rect 1452 13200 1458 13252
rect 1762 13200 1768 13252
rect 1820 13200 1826 13252
rect 4338 13132 4344 13184
rect 4396 13132 4402 13184
rect 1104 13082 5035 13104
rect 1104 13030 1892 13082
rect 1944 13030 1956 13082
rect 2008 13030 2020 13082
rect 2072 13030 2084 13082
rect 2136 13030 2148 13082
rect 2200 13030 2835 13082
rect 2887 13030 2899 13082
rect 2951 13030 2963 13082
rect 3015 13030 3027 13082
rect 3079 13030 3091 13082
rect 3143 13030 3778 13082
rect 3830 13030 3842 13082
rect 3894 13030 3906 13082
rect 3958 13030 3970 13082
rect 4022 13030 4034 13082
rect 4086 13030 4721 13082
rect 4773 13030 4785 13082
rect 4837 13030 4849 13082
rect 4901 13030 4913 13082
rect 4965 13030 4977 13082
rect 5029 13030 5035 13082
rect 1104 13008 5035 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 1820 12940 2881 12968
rect 1820 12928 1826 12940
rect 2869 12937 2881 12940
rect 2915 12937 2927 12971
rect 2869 12931 2927 12937
rect 4338 12928 4344 12980
rect 4396 12928 4402 12980
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 4356 12832 4384 12928
rect 3099 12804 4384 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 1104 12538 4876 12560
rect 1104 12486 1421 12538
rect 1473 12486 1485 12538
rect 1537 12486 1549 12538
rect 1601 12486 1613 12538
rect 1665 12486 1677 12538
rect 1729 12486 2364 12538
rect 2416 12486 2428 12538
rect 2480 12486 2492 12538
rect 2544 12486 2556 12538
rect 2608 12486 2620 12538
rect 2672 12486 3307 12538
rect 3359 12486 3371 12538
rect 3423 12486 3435 12538
rect 3487 12486 3499 12538
rect 3551 12486 3563 12538
rect 3615 12486 4250 12538
rect 4302 12486 4314 12538
rect 4366 12486 4378 12538
rect 4430 12486 4442 12538
rect 4494 12486 4506 12538
rect 4558 12486 4876 12538
rect 1104 12464 4876 12486
rect 1104 11994 5035 12016
rect 1104 11942 1892 11994
rect 1944 11942 1956 11994
rect 2008 11942 2020 11994
rect 2072 11942 2084 11994
rect 2136 11942 2148 11994
rect 2200 11942 2835 11994
rect 2887 11942 2899 11994
rect 2951 11942 2963 11994
rect 3015 11942 3027 11994
rect 3079 11942 3091 11994
rect 3143 11942 3778 11994
rect 3830 11942 3842 11994
rect 3894 11942 3906 11994
rect 3958 11942 3970 11994
rect 4022 11942 4034 11994
rect 4086 11942 4721 11994
rect 4773 11942 4785 11994
rect 4837 11942 4849 11994
rect 4901 11942 4913 11994
rect 4965 11942 4977 11994
rect 5029 11942 5035 11994
rect 1104 11920 5035 11942
rect 1104 11450 4876 11472
rect 1104 11398 1421 11450
rect 1473 11398 1485 11450
rect 1537 11398 1549 11450
rect 1601 11398 1613 11450
rect 1665 11398 1677 11450
rect 1729 11398 2364 11450
rect 2416 11398 2428 11450
rect 2480 11398 2492 11450
rect 2544 11398 2556 11450
rect 2608 11398 2620 11450
rect 2672 11398 3307 11450
rect 3359 11398 3371 11450
rect 3423 11398 3435 11450
rect 3487 11398 3499 11450
rect 3551 11398 3563 11450
rect 3615 11398 4250 11450
rect 4302 11398 4314 11450
rect 4366 11398 4378 11450
rect 4430 11398 4442 11450
rect 4494 11398 4506 11450
rect 4558 11398 4876 11450
rect 1104 11376 4876 11398
rect 1104 10906 5035 10928
rect 1104 10854 1892 10906
rect 1944 10854 1956 10906
rect 2008 10854 2020 10906
rect 2072 10854 2084 10906
rect 2136 10854 2148 10906
rect 2200 10854 2835 10906
rect 2887 10854 2899 10906
rect 2951 10854 2963 10906
rect 3015 10854 3027 10906
rect 3079 10854 3091 10906
rect 3143 10854 3778 10906
rect 3830 10854 3842 10906
rect 3894 10854 3906 10906
rect 3958 10854 3970 10906
rect 4022 10854 4034 10906
rect 4086 10854 4721 10906
rect 4773 10854 4785 10906
rect 4837 10854 4849 10906
rect 4901 10854 4913 10906
rect 4965 10854 4977 10906
rect 5029 10854 5035 10906
rect 1104 10832 5035 10854
rect 1104 10362 4876 10384
rect 1104 10310 1421 10362
rect 1473 10310 1485 10362
rect 1537 10310 1549 10362
rect 1601 10310 1613 10362
rect 1665 10310 1677 10362
rect 1729 10310 2364 10362
rect 2416 10310 2428 10362
rect 2480 10310 2492 10362
rect 2544 10310 2556 10362
rect 2608 10310 2620 10362
rect 2672 10310 3307 10362
rect 3359 10310 3371 10362
rect 3423 10310 3435 10362
rect 3487 10310 3499 10362
rect 3551 10310 3563 10362
rect 3615 10310 4250 10362
rect 4302 10310 4314 10362
rect 4366 10310 4378 10362
rect 4430 10310 4442 10362
rect 4494 10310 4506 10362
rect 4558 10310 4876 10362
rect 1104 10288 4876 10310
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 4540 10124 4568 10211
rect 4522 10072 4528 10124
rect 4580 10072 4586 10124
rect 1104 9818 5035 9840
rect 1104 9766 1892 9818
rect 1944 9766 1956 9818
rect 2008 9766 2020 9818
rect 2072 9766 2084 9818
rect 2136 9766 2148 9818
rect 2200 9766 2835 9818
rect 2887 9766 2899 9818
rect 2951 9766 2963 9818
rect 3015 9766 3027 9818
rect 3079 9766 3091 9818
rect 3143 9766 3778 9818
rect 3830 9766 3842 9818
rect 3894 9766 3906 9818
rect 3958 9766 3970 9818
rect 4022 9766 4034 9818
rect 4086 9766 4721 9818
rect 4773 9766 4785 9818
rect 4837 9766 4849 9818
rect 4901 9766 4913 9818
rect 4965 9766 4977 9818
rect 5029 9766 5035 9818
rect 1104 9744 5035 9766
rect 1104 9274 4876 9296
rect 1104 9222 1421 9274
rect 1473 9222 1485 9274
rect 1537 9222 1549 9274
rect 1601 9222 1613 9274
rect 1665 9222 1677 9274
rect 1729 9222 2364 9274
rect 2416 9222 2428 9274
rect 2480 9222 2492 9274
rect 2544 9222 2556 9274
rect 2608 9222 2620 9274
rect 2672 9222 3307 9274
rect 3359 9222 3371 9274
rect 3423 9222 3435 9274
rect 3487 9222 3499 9274
rect 3551 9222 3563 9274
rect 3615 9222 4250 9274
rect 4302 9222 4314 9274
rect 4366 9222 4378 9274
rect 4430 9222 4442 9274
rect 4494 9222 4506 9274
rect 4558 9222 4876 9274
rect 1104 9200 4876 9222
rect 1104 8730 5035 8752
rect 1104 8678 1892 8730
rect 1944 8678 1956 8730
rect 2008 8678 2020 8730
rect 2072 8678 2084 8730
rect 2136 8678 2148 8730
rect 2200 8678 2835 8730
rect 2887 8678 2899 8730
rect 2951 8678 2963 8730
rect 3015 8678 3027 8730
rect 3079 8678 3091 8730
rect 3143 8678 3778 8730
rect 3830 8678 3842 8730
rect 3894 8678 3906 8730
rect 3958 8678 3970 8730
rect 4022 8678 4034 8730
rect 4086 8678 4721 8730
rect 4773 8678 4785 8730
rect 4837 8678 4849 8730
rect 4901 8678 4913 8730
rect 4965 8678 4977 8730
rect 5029 8678 5035 8730
rect 1104 8656 5035 8678
rect 1104 8186 4876 8208
rect 1104 8134 1421 8186
rect 1473 8134 1485 8186
rect 1537 8134 1549 8186
rect 1601 8134 1613 8186
rect 1665 8134 1677 8186
rect 1729 8134 2364 8186
rect 2416 8134 2428 8186
rect 2480 8134 2492 8186
rect 2544 8134 2556 8186
rect 2608 8134 2620 8186
rect 2672 8134 3307 8186
rect 3359 8134 3371 8186
rect 3423 8134 3435 8186
rect 3487 8134 3499 8186
rect 3551 8134 3563 8186
rect 3615 8134 4250 8186
rect 4302 8134 4314 8186
rect 4366 8134 4378 8186
rect 4430 8134 4442 8186
rect 4494 8134 4506 8186
rect 4558 8134 4876 8186
rect 1104 8112 4876 8134
rect 1104 7642 5035 7664
rect 1104 7590 1892 7642
rect 1944 7590 1956 7642
rect 2008 7590 2020 7642
rect 2072 7590 2084 7642
rect 2136 7590 2148 7642
rect 2200 7590 2835 7642
rect 2887 7590 2899 7642
rect 2951 7590 2963 7642
rect 3015 7590 3027 7642
rect 3079 7590 3091 7642
rect 3143 7590 3778 7642
rect 3830 7590 3842 7642
rect 3894 7590 3906 7642
rect 3958 7590 3970 7642
rect 4022 7590 4034 7642
rect 4086 7590 4721 7642
rect 4773 7590 4785 7642
rect 4837 7590 4849 7642
rect 4901 7590 4913 7642
rect 4965 7590 4977 7642
rect 5029 7590 5035 7642
rect 1104 7568 5035 7590
rect 1104 7098 4876 7120
rect 1104 7046 1421 7098
rect 1473 7046 1485 7098
rect 1537 7046 1549 7098
rect 1601 7046 1613 7098
rect 1665 7046 1677 7098
rect 1729 7046 2364 7098
rect 2416 7046 2428 7098
rect 2480 7046 2492 7098
rect 2544 7046 2556 7098
rect 2608 7046 2620 7098
rect 2672 7046 3307 7098
rect 3359 7046 3371 7098
rect 3423 7046 3435 7098
rect 3487 7046 3499 7098
rect 3551 7046 3563 7098
rect 3615 7046 4250 7098
rect 4302 7046 4314 7098
rect 4366 7046 4378 7098
rect 4430 7046 4442 7098
rect 4494 7046 4506 7098
rect 4558 7046 4876 7098
rect 1104 7024 4876 7046
rect 1104 6554 5035 6576
rect 1104 6502 1892 6554
rect 1944 6502 1956 6554
rect 2008 6502 2020 6554
rect 2072 6502 2084 6554
rect 2136 6502 2148 6554
rect 2200 6502 2835 6554
rect 2887 6502 2899 6554
rect 2951 6502 2963 6554
rect 3015 6502 3027 6554
rect 3079 6502 3091 6554
rect 3143 6502 3778 6554
rect 3830 6502 3842 6554
rect 3894 6502 3906 6554
rect 3958 6502 3970 6554
rect 4022 6502 4034 6554
rect 4086 6502 4721 6554
rect 4773 6502 4785 6554
rect 4837 6502 4849 6554
rect 4901 6502 4913 6554
rect 4965 6502 4977 6554
rect 5029 6502 5035 6554
rect 1104 6480 5035 6502
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 1820 6276 3157 6304
rect 1820 6264 1826 6276
rect 3145 6273 3157 6276
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 3412 6307 3470 6313
rect 3412 6273 3424 6307
rect 3458 6304 3470 6307
rect 4154 6304 4160 6316
rect 3458 6276 4160 6304
rect 3458 6273 3470 6276
rect 3412 6267 3470 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 1104 6010 4876 6032
rect 1104 5958 1421 6010
rect 1473 5958 1485 6010
rect 1537 5958 1549 6010
rect 1601 5958 1613 6010
rect 1665 5958 1677 6010
rect 1729 5958 2364 6010
rect 2416 5958 2428 6010
rect 2480 5958 2492 6010
rect 2544 5958 2556 6010
rect 2608 5958 2620 6010
rect 2672 5958 3307 6010
rect 3359 5958 3371 6010
rect 3423 5958 3435 6010
rect 3487 5958 3499 6010
rect 3551 5958 3563 6010
rect 3615 5958 4250 6010
rect 4302 5958 4314 6010
rect 4366 5958 4378 6010
rect 4430 5958 4442 6010
rect 4494 5958 4506 6010
rect 4558 5958 4876 6010
rect 1104 5936 4876 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4798 5896 4804 5908
rect 4387 5868 4804 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4614 5692 4620 5704
rect 4571 5664 4620 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 1104 5466 5035 5488
rect 1104 5414 1892 5466
rect 1944 5414 1956 5466
rect 2008 5414 2020 5466
rect 2072 5414 2084 5466
rect 2136 5414 2148 5466
rect 2200 5414 2835 5466
rect 2887 5414 2899 5466
rect 2951 5414 2963 5466
rect 3015 5414 3027 5466
rect 3079 5414 3091 5466
rect 3143 5414 3778 5466
rect 3830 5414 3842 5466
rect 3894 5414 3906 5466
rect 3958 5414 3970 5466
rect 4022 5414 4034 5466
rect 4086 5414 4721 5466
rect 4773 5414 4785 5466
rect 4837 5414 4849 5466
rect 4901 5414 4913 5466
rect 4965 5414 4977 5466
rect 5029 5414 5035 5466
rect 1104 5392 5035 5414
rect 1104 4922 4876 4944
rect 1104 4870 1421 4922
rect 1473 4870 1485 4922
rect 1537 4870 1549 4922
rect 1601 4870 1613 4922
rect 1665 4870 1677 4922
rect 1729 4870 2364 4922
rect 2416 4870 2428 4922
rect 2480 4870 2492 4922
rect 2544 4870 2556 4922
rect 2608 4870 2620 4922
rect 2672 4870 3307 4922
rect 3359 4870 3371 4922
rect 3423 4870 3435 4922
rect 3487 4870 3499 4922
rect 3551 4870 3563 4922
rect 3615 4870 4250 4922
rect 4302 4870 4314 4922
rect 4366 4870 4378 4922
rect 4430 4870 4442 4922
rect 4494 4870 4506 4922
rect 4558 4870 4876 4922
rect 1104 4848 4876 4870
rect 1104 4378 5035 4400
rect 1104 4326 1892 4378
rect 1944 4326 1956 4378
rect 2008 4326 2020 4378
rect 2072 4326 2084 4378
rect 2136 4326 2148 4378
rect 2200 4326 2835 4378
rect 2887 4326 2899 4378
rect 2951 4326 2963 4378
rect 3015 4326 3027 4378
rect 3079 4326 3091 4378
rect 3143 4326 3778 4378
rect 3830 4326 3842 4378
rect 3894 4326 3906 4378
rect 3958 4326 3970 4378
rect 4022 4326 4034 4378
rect 4086 4326 4721 4378
rect 4773 4326 4785 4378
rect 4837 4326 4849 4378
rect 4901 4326 4913 4378
rect 4965 4326 4977 4378
rect 5029 4326 5035 4378
rect 1104 4304 5035 4326
rect 1104 3834 4876 3856
rect 1104 3782 1421 3834
rect 1473 3782 1485 3834
rect 1537 3782 1549 3834
rect 1601 3782 1613 3834
rect 1665 3782 1677 3834
rect 1729 3782 2364 3834
rect 2416 3782 2428 3834
rect 2480 3782 2492 3834
rect 2544 3782 2556 3834
rect 2608 3782 2620 3834
rect 2672 3782 3307 3834
rect 3359 3782 3371 3834
rect 3423 3782 3435 3834
rect 3487 3782 3499 3834
rect 3551 3782 3563 3834
rect 3615 3782 4250 3834
rect 4302 3782 4314 3834
rect 4366 3782 4378 3834
rect 4430 3782 4442 3834
rect 4494 3782 4506 3834
rect 4558 3782 4876 3834
rect 1104 3760 4876 3782
rect 1104 3290 5035 3312
rect 1104 3238 1892 3290
rect 1944 3238 1956 3290
rect 2008 3238 2020 3290
rect 2072 3238 2084 3290
rect 2136 3238 2148 3290
rect 2200 3238 2835 3290
rect 2887 3238 2899 3290
rect 2951 3238 2963 3290
rect 3015 3238 3027 3290
rect 3079 3238 3091 3290
rect 3143 3238 3778 3290
rect 3830 3238 3842 3290
rect 3894 3238 3906 3290
rect 3958 3238 3970 3290
rect 4022 3238 4034 3290
rect 4086 3238 4721 3290
rect 4773 3238 4785 3290
rect 4837 3238 4849 3290
rect 4901 3238 4913 3290
rect 4965 3238 4977 3290
rect 5029 3238 5035 3290
rect 1104 3216 5035 3238
rect 1104 2746 4876 2768
rect 1104 2694 1421 2746
rect 1473 2694 1485 2746
rect 1537 2694 1549 2746
rect 1601 2694 1613 2746
rect 1665 2694 1677 2746
rect 1729 2694 2364 2746
rect 2416 2694 2428 2746
rect 2480 2694 2492 2746
rect 2544 2694 2556 2746
rect 2608 2694 2620 2746
rect 2672 2694 3307 2746
rect 3359 2694 3371 2746
rect 3423 2694 3435 2746
rect 3487 2694 3499 2746
rect 3551 2694 3563 2746
rect 3615 2694 4250 2746
rect 4302 2694 4314 2746
rect 4366 2694 4378 2746
rect 4430 2694 4442 2746
rect 4494 2694 4506 2746
rect 4558 2694 4876 2746
rect 1104 2672 4876 2694
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4341 2635 4399 2641
rect 4341 2632 4353 2635
rect 4212 2604 4353 2632
rect 4212 2592 4218 2604
rect 4341 2601 4353 2604
rect 4387 2601 4399 2635
rect 4341 2595 4399 2601
rect 4890 2456 4896 2508
rect 4948 2456 4954 2508
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4908 2428 4936 2456
rect 4571 2400 4936 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 1104 2202 5035 2224
rect 1104 2150 1892 2202
rect 1944 2150 1956 2202
rect 2008 2150 2020 2202
rect 2072 2150 2084 2202
rect 2136 2150 2148 2202
rect 2200 2150 2835 2202
rect 2887 2150 2899 2202
rect 2951 2150 2963 2202
rect 3015 2150 3027 2202
rect 3079 2150 3091 2202
rect 3143 2150 3778 2202
rect 3830 2150 3842 2202
rect 3894 2150 3906 2202
rect 3958 2150 3970 2202
rect 4022 2150 4034 2202
rect 4086 2150 4721 2202
rect 4773 2150 4785 2202
rect 4837 2150 4849 2202
rect 4901 2150 4913 2202
rect 4965 2150 4977 2202
rect 5029 2150 5035 2202
rect 1104 2128 5035 2150
<< via1 >>
rect 1421 13574 1473 13626
rect 1485 13574 1537 13626
rect 1549 13574 1601 13626
rect 1613 13574 1665 13626
rect 1677 13574 1729 13626
rect 2364 13574 2416 13626
rect 2428 13574 2480 13626
rect 2492 13574 2544 13626
rect 2556 13574 2608 13626
rect 2620 13574 2672 13626
rect 3307 13574 3359 13626
rect 3371 13574 3423 13626
rect 3435 13574 3487 13626
rect 3499 13574 3551 13626
rect 3563 13574 3615 13626
rect 4250 13574 4302 13626
rect 4314 13574 4366 13626
rect 4378 13574 4430 13626
rect 4442 13574 4494 13626
rect 4506 13574 4558 13626
rect 4896 13268 4948 13320
rect 1400 13243 1452 13252
rect 1400 13209 1409 13243
rect 1409 13209 1443 13243
rect 1443 13209 1452 13243
rect 1400 13200 1452 13209
rect 1768 13243 1820 13252
rect 1768 13209 1777 13243
rect 1777 13209 1811 13243
rect 1811 13209 1820 13243
rect 1768 13200 1820 13209
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 1892 13030 1944 13082
rect 1956 13030 2008 13082
rect 2020 13030 2072 13082
rect 2084 13030 2136 13082
rect 2148 13030 2200 13082
rect 2835 13030 2887 13082
rect 2899 13030 2951 13082
rect 2963 13030 3015 13082
rect 3027 13030 3079 13082
rect 3091 13030 3143 13082
rect 3778 13030 3830 13082
rect 3842 13030 3894 13082
rect 3906 13030 3958 13082
rect 3970 13030 4022 13082
rect 4034 13030 4086 13082
rect 4721 13030 4773 13082
rect 4785 13030 4837 13082
rect 4849 13030 4901 13082
rect 4913 13030 4965 13082
rect 4977 13030 5029 13082
rect 1768 12928 1820 12980
rect 4344 12928 4396 12980
rect 1421 12486 1473 12538
rect 1485 12486 1537 12538
rect 1549 12486 1601 12538
rect 1613 12486 1665 12538
rect 1677 12486 1729 12538
rect 2364 12486 2416 12538
rect 2428 12486 2480 12538
rect 2492 12486 2544 12538
rect 2556 12486 2608 12538
rect 2620 12486 2672 12538
rect 3307 12486 3359 12538
rect 3371 12486 3423 12538
rect 3435 12486 3487 12538
rect 3499 12486 3551 12538
rect 3563 12486 3615 12538
rect 4250 12486 4302 12538
rect 4314 12486 4366 12538
rect 4378 12486 4430 12538
rect 4442 12486 4494 12538
rect 4506 12486 4558 12538
rect 1892 11942 1944 11994
rect 1956 11942 2008 11994
rect 2020 11942 2072 11994
rect 2084 11942 2136 11994
rect 2148 11942 2200 11994
rect 2835 11942 2887 11994
rect 2899 11942 2951 11994
rect 2963 11942 3015 11994
rect 3027 11942 3079 11994
rect 3091 11942 3143 11994
rect 3778 11942 3830 11994
rect 3842 11942 3894 11994
rect 3906 11942 3958 11994
rect 3970 11942 4022 11994
rect 4034 11942 4086 11994
rect 4721 11942 4773 11994
rect 4785 11942 4837 11994
rect 4849 11942 4901 11994
rect 4913 11942 4965 11994
rect 4977 11942 5029 11994
rect 1421 11398 1473 11450
rect 1485 11398 1537 11450
rect 1549 11398 1601 11450
rect 1613 11398 1665 11450
rect 1677 11398 1729 11450
rect 2364 11398 2416 11450
rect 2428 11398 2480 11450
rect 2492 11398 2544 11450
rect 2556 11398 2608 11450
rect 2620 11398 2672 11450
rect 3307 11398 3359 11450
rect 3371 11398 3423 11450
rect 3435 11398 3487 11450
rect 3499 11398 3551 11450
rect 3563 11398 3615 11450
rect 4250 11398 4302 11450
rect 4314 11398 4366 11450
rect 4378 11398 4430 11450
rect 4442 11398 4494 11450
rect 4506 11398 4558 11450
rect 1892 10854 1944 10906
rect 1956 10854 2008 10906
rect 2020 10854 2072 10906
rect 2084 10854 2136 10906
rect 2148 10854 2200 10906
rect 2835 10854 2887 10906
rect 2899 10854 2951 10906
rect 2963 10854 3015 10906
rect 3027 10854 3079 10906
rect 3091 10854 3143 10906
rect 3778 10854 3830 10906
rect 3842 10854 3894 10906
rect 3906 10854 3958 10906
rect 3970 10854 4022 10906
rect 4034 10854 4086 10906
rect 4721 10854 4773 10906
rect 4785 10854 4837 10906
rect 4849 10854 4901 10906
rect 4913 10854 4965 10906
rect 4977 10854 5029 10906
rect 1421 10310 1473 10362
rect 1485 10310 1537 10362
rect 1549 10310 1601 10362
rect 1613 10310 1665 10362
rect 1677 10310 1729 10362
rect 2364 10310 2416 10362
rect 2428 10310 2480 10362
rect 2492 10310 2544 10362
rect 2556 10310 2608 10362
rect 2620 10310 2672 10362
rect 3307 10310 3359 10362
rect 3371 10310 3423 10362
rect 3435 10310 3487 10362
rect 3499 10310 3551 10362
rect 3563 10310 3615 10362
rect 4250 10310 4302 10362
rect 4314 10310 4366 10362
rect 4378 10310 4430 10362
rect 4442 10310 4494 10362
rect 4506 10310 4558 10362
rect 4528 10072 4580 10124
rect 1892 9766 1944 9818
rect 1956 9766 2008 9818
rect 2020 9766 2072 9818
rect 2084 9766 2136 9818
rect 2148 9766 2200 9818
rect 2835 9766 2887 9818
rect 2899 9766 2951 9818
rect 2963 9766 3015 9818
rect 3027 9766 3079 9818
rect 3091 9766 3143 9818
rect 3778 9766 3830 9818
rect 3842 9766 3894 9818
rect 3906 9766 3958 9818
rect 3970 9766 4022 9818
rect 4034 9766 4086 9818
rect 4721 9766 4773 9818
rect 4785 9766 4837 9818
rect 4849 9766 4901 9818
rect 4913 9766 4965 9818
rect 4977 9766 5029 9818
rect 1421 9222 1473 9274
rect 1485 9222 1537 9274
rect 1549 9222 1601 9274
rect 1613 9222 1665 9274
rect 1677 9222 1729 9274
rect 2364 9222 2416 9274
rect 2428 9222 2480 9274
rect 2492 9222 2544 9274
rect 2556 9222 2608 9274
rect 2620 9222 2672 9274
rect 3307 9222 3359 9274
rect 3371 9222 3423 9274
rect 3435 9222 3487 9274
rect 3499 9222 3551 9274
rect 3563 9222 3615 9274
rect 4250 9222 4302 9274
rect 4314 9222 4366 9274
rect 4378 9222 4430 9274
rect 4442 9222 4494 9274
rect 4506 9222 4558 9274
rect 1892 8678 1944 8730
rect 1956 8678 2008 8730
rect 2020 8678 2072 8730
rect 2084 8678 2136 8730
rect 2148 8678 2200 8730
rect 2835 8678 2887 8730
rect 2899 8678 2951 8730
rect 2963 8678 3015 8730
rect 3027 8678 3079 8730
rect 3091 8678 3143 8730
rect 3778 8678 3830 8730
rect 3842 8678 3894 8730
rect 3906 8678 3958 8730
rect 3970 8678 4022 8730
rect 4034 8678 4086 8730
rect 4721 8678 4773 8730
rect 4785 8678 4837 8730
rect 4849 8678 4901 8730
rect 4913 8678 4965 8730
rect 4977 8678 5029 8730
rect 1421 8134 1473 8186
rect 1485 8134 1537 8186
rect 1549 8134 1601 8186
rect 1613 8134 1665 8186
rect 1677 8134 1729 8186
rect 2364 8134 2416 8186
rect 2428 8134 2480 8186
rect 2492 8134 2544 8186
rect 2556 8134 2608 8186
rect 2620 8134 2672 8186
rect 3307 8134 3359 8186
rect 3371 8134 3423 8186
rect 3435 8134 3487 8186
rect 3499 8134 3551 8186
rect 3563 8134 3615 8186
rect 4250 8134 4302 8186
rect 4314 8134 4366 8186
rect 4378 8134 4430 8186
rect 4442 8134 4494 8186
rect 4506 8134 4558 8186
rect 1892 7590 1944 7642
rect 1956 7590 2008 7642
rect 2020 7590 2072 7642
rect 2084 7590 2136 7642
rect 2148 7590 2200 7642
rect 2835 7590 2887 7642
rect 2899 7590 2951 7642
rect 2963 7590 3015 7642
rect 3027 7590 3079 7642
rect 3091 7590 3143 7642
rect 3778 7590 3830 7642
rect 3842 7590 3894 7642
rect 3906 7590 3958 7642
rect 3970 7590 4022 7642
rect 4034 7590 4086 7642
rect 4721 7590 4773 7642
rect 4785 7590 4837 7642
rect 4849 7590 4901 7642
rect 4913 7590 4965 7642
rect 4977 7590 5029 7642
rect 1421 7046 1473 7098
rect 1485 7046 1537 7098
rect 1549 7046 1601 7098
rect 1613 7046 1665 7098
rect 1677 7046 1729 7098
rect 2364 7046 2416 7098
rect 2428 7046 2480 7098
rect 2492 7046 2544 7098
rect 2556 7046 2608 7098
rect 2620 7046 2672 7098
rect 3307 7046 3359 7098
rect 3371 7046 3423 7098
rect 3435 7046 3487 7098
rect 3499 7046 3551 7098
rect 3563 7046 3615 7098
rect 4250 7046 4302 7098
rect 4314 7046 4366 7098
rect 4378 7046 4430 7098
rect 4442 7046 4494 7098
rect 4506 7046 4558 7098
rect 1892 6502 1944 6554
rect 1956 6502 2008 6554
rect 2020 6502 2072 6554
rect 2084 6502 2136 6554
rect 2148 6502 2200 6554
rect 2835 6502 2887 6554
rect 2899 6502 2951 6554
rect 2963 6502 3015 6554
rect 3027 6502 3079 6554
rect 3091 6502 3143 6554
rect 3778 6502 3830 6554
rect 3842 6502 3894 6554
rect 3906 6502 3958 6554
rect 3970 6502 4022 6554
rect 4034 6502 4086 6554
rect 4721 6502 4773 6554
rect 4785 6502 4837 6554
rect 4849 6502 4901 6554
rect 4913 6502 4965 6554
rect 4977 6502 5029 6554
rect 1768 6264 1820 6316
rect 4160 6264 4212 6316
rect 4620 6060 4672 6112
rect 1421 5958 1473 6010
rect 1485 5958 1537 6010
rect 1549 5958 1601 6010
rect 1613 5958 1665 6010
rect 1677 5958 1729 6010
rect 2364 5958 2416 6010
rect 2428 5958 2480 6010
rect 2492 5958 2544 6010
rect 2556 5958 2608 6010
rect 2620 5958 2672 6010
rect 3307 5958 3359 6010
rect 3371 5958 3423 6010
rect 3435 5958 3487 6010
rect 3499 5958 3551 6010
rect 3563 5958 3615 6010
rect 4250 5958 4302 6010
rect 4314 5958 4366 6010
rect 4378 5958 4430 6010
rect 4442 5958 4494 6010
rect 4506 5958 4558 6010
rect 4804 5856 4856 5908
rect 4620 5652 4672 5704
rect 1892 5414 1944 5466
rect 1956 5414 2008 5466
rect 2020 5414 2072 5466
rect 2084 5414 2136 5466
rect 2148 5414 2200 5466
rect 2835 5414 2887 5466
rect 2899 5414 2951 5466
rect 2963 5414 3015 5466
rect 3027 5414 3079 5466
rect 3091 5414 3143 5466
rect 3778 5414 3830 5466
rect 3842 5414 3894 5466
rect 3906 5414 3958 5466
rect 3970 5414 4022 5466
rect 4034 5414 4086 5466
rect 4721 5414 4773 5466
rect 4785 5414 4837 5466
rect 4849 5414 4901 5466
rect 4913 5414 4965 5466
rect 4977 5414 5029 5466
rect 1421 4870 1473 4922
rect 1485 4870 1537 4922
rect 1549 4870 1601 4922
rect 1613 4870 1665 4922
rect 1677 4870 1729 4922
rect 2364 4870 2416 4922
rect 2428 4870 2480 4922
rect 2492 4870 2544 4922
rect 2556 4870 2608 4922
rect 2620 4870 2672 4922
rect 3307 4870 3359 4922
rect 3371 4870 3423 4922
rect 3435 4870 3487 4922
rect 3499 4870 3551 4922
rect 3563 4870 3615 4922
rect 4250 4870 4302 4922
rect 4314 4870 4366 4922
rect 4378 4870 4430 4922
rect 4442 4870 4494 4922
rect 4506 4870 4558 4922
rect 1892 4326 1944 4378
rect 1956 4326 2008 4378
rect 2020 4326 2072 4378
rect 2084 4326 2136 4378
rect 2148 4326 2200 4378
rect 2835 4326 2887 4378
rect 2899 4326 2951 4378
rect 2963 4326 3015 4378
rect 3027 4326 3079 4378
rect 3091 4326 3143 4378
rect 3778 4326 3830 4378
rect 3842 4326 3894 4378
rect 3906 4326 3958 4378
rect 3970 4326 4022 4378
rect 4034 4326 4086 4378
rect 4721 4326 4773 4378
rect 4785 4326 4837 4378
rect 4849 4326 4901 4378
rect 4913 4326 4965 4378
rect 4977 4326 5029 4378
rect 1421 3782 1473 3834
rect 1485 3782 1537 3834
rect 1549 3782 1601 3834
rect 1613 3782 1665 3834
rect 1677 3782 1729 3834
rect 2364 3782 2416 3834
rect 2428 3782 2480 3834
rect 2492 3782 2544 3834
rect 2556 3782 2608 3834
rect 2620 3782 2672 3834
rect 3307 3782 3359 3834
rect 3371 3782 3423 3834
rect 3435 3782 3487 3834
rect 3499 3782 3551 3834
rect 3563 3782 3615 3834
rect 4250 3782 4302 3834
rect 4314 3782 4366 3834
rect 4378 3782 4430 3834
rect 4442 3782 4494 3834
rect 4506 3782 4558 3834
rect 1892 3238 1944 3290
rect 1956 3238 2008 3290
rect 2020 3238 2072 3290
rect 2084 3238 2136 3290
rect 2148 3238 2200 3290
rect 2835 3238 2887 3290
rect 2899 3238 2951 3290
rect 2963 3238 3015 3290
rect 3027 3238 3079 3290
rect 3091 3238 3143 3290
rect 3778 3238 3830 3290
rect 3842 3238 3894 3290
rect 3906 3238 3958 3290
rect 3970 3238 4022 3290
rect 4034 3238 4086 3290
rect 4721 3238 4773 3290
rect 4785 3238 4837 3290
rect 4849 3238 4901 3290
rect 4913 3238 4965 3290
rect 4977 3238 5029 3290
rect 1421 2694 1473 2746
rect 1485 2694 1537 2746
rect 1549 2694 1601 2746
rect 1613 2694 1665 2746
rect 1677 2694 1729 2746
rect 2364 2694 2416 2746
rect 2428 2694 2480 2746
rect 2492 2694 2544 2746
rect 2556 2694 2608 2746
rect 2620 2694 2672 2746
rect 3307 2694 3359 2746
rect 3371 2694 3423 2746
rect 3435 2694 3487 2746
rect 3499 2694 3551 2746
rect 3563 2694 3615 2746
rect 4250 2694 4302 2746
rect 4314 2694 4366 2746
rect 4378 2694 4430 2746
rect 4442 2694 4494 2746
rect 4506 2694 4558 2746
rect 4160 2592 4212 2644
rect 4896 2456 4948 2508
rect 1892 2150 1944 2202
rect 1956 2150 2008 2202
rect 2020 2150 2072 2202
rect 2084 2150 2136 2202
rect 2148 2150 2200 2202
rect 2835 2150 2887 2202
rect 2899 2150 2951 2202
rect 2963 2150 3015 2202
rect 3027 2150 3079 2202
rect 3091 2150 3143 2202
rect 3778 2150 3830 2202
rect 3842 2150 3894 2202
rect 3906 2150 3958 2202
rect 3970 2150 4022 2202
rect 4034 2150 4086 2202
rect 4721 2150 4773 2202
rect 4785 2150 4837 2202
rect 4849 2150 4901 2202
rect 4913 2150 4965 2202
rect 4977 2150 5029 2202
<< metal2 >>
rect 4894 13696 4950 13705
rect 1421 13628 1729 13637
rect 1421 13626 1427 13628
rect 1483 13626 1507 13628
rect 1563 13626 1587 13628
rect 1643 13626 1667 13628
rect 1723 13626 1729 13628
rect 1483 13574 1485 13626
rect 1665 13574 1667 13626
rect 1421 13572 1427 13574
rect 1483 13572 1507 13574
rect 1563 13572 1587 13574
rect 1643 13572 1667 13574
rect 1723 13572 1729 13574
rect 1421 13563 1729 13572
rect 2364 13628 2672 13637
rect 2364 13626 2370 13628
rect 2426 13626 2450 13628
rect 2506 13626 2530 13628
rect 2586 13626 2610 13628
rect 2666 13626 2672 13628
rect 2426 13574 2428 13626
rect 2608 13574 2610 13626
rect 2364 13572 2370 13574
rect 2426 13572 2450 13574
rect 2506 13572 2530 13574
rect 2586 13572 2610 13574
rect 2666 13572 2672 13574
rect 2364 13563 2672 13572
rect 3307 13628 3615 13637
rect 3307 13626 3313 13628
rect 3369 13626 3393 13628
rect 3449 13626 3473 13628
rect 3529 13626 3553 13628
rect 3609 13626 3615 13628
rect 3369 13574 3371 13626
rect 3551 13574 3553 13626
rect 3307 13572 3313 13574
rect 3369 13572 3393 13574
rect 3449 13572 3473 13574
rect 3529 13572 3553 13574
rect 3609 13572 3615 13574
rect 3307 13563 3615 13572
rect 4250 13628 4558 13637
rect 4894 13631 4950 13640
rect 4250 13626 4256 13628
rect 4312 13626 4336 13628
rect 4392 13626 4416 13628
rect 4472 13626 4496 13628
rect 4552 13626 4558 13628
rect 4312 13574 4314 13626
rect 4494 13574 4496 13626
rect 4250 13572 4256 13574
rect 4312 13572 4336 13574
rect 4392 13572 4416 13574
rect 4472 13572 4496 13574
rect 4552 13572 4558 13574
rect 4250 13563 4558 13572
rect 4908 13326 4936 13631
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1412 13161 1440 13194
rect 1398 13152 1454 13161
rect 1398 13087 1454 13096
rect 1780 12986 1808 13194
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 1892 13084 2200 13093
rect 1892 13082 1898 13084
rect 1954 13082 1978 13084
rect 2034 13082 2058 13084
rect 2114 13082 2138 13084
rect 2194 13082 2200 13084
rect 1954 13030 1956 13082
rect 2136 13030 2138 13082
rect 1892 13028 1898 13030
rect 1954 13028 1978 13030
rect 2034 13028 2058 13030
rect 2114 13028 2138 13030
rect 2194 13028 2200 13030
rect 1892 13019 2200 13028
rect 2835 13084 3143 13093
rect 2835 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3081 13084
rect 3137 13082 3143 13084
rect 2897 13030 2899 13082
rect 3079 13030 3081 13082
rect 2835 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3081 13030
rect 3137 13028 3143 13030
rect 2835 13019 3143 13028
rect 3778 13084 4086 13093
rect 3778 13082 3784 13084
rect 3840 13082 3864 13084
rect 3920 13082 3944 13084
rect 4000 13082 4024 13084
rect 4080 13082 4086 13084
rect 3840 13030 3842 13082
rect 4022 13030 4024 13082
rect 3778 13028 3784 13030
rect 3840 13028 3864 13030
rect 3920 13028 3944 13030
rect 4000 13028 4024 13030
rect 4080 13028 4086 13030
rect 3778 13019 4086 13028
rect 4356 12986 4384 13126
rect 4721 13084 5029 13093
rect 4721 13082 4727 13084
rect 4783 13082 4807 13084
rect 4863 13082 4887 13084
rect 4943 13082 4967 13084
rect 5023 13082 5029 13084
rect 4783 13030 4785 13082
rect 4965 13030 4967 13082
rect 4721 13028 4727 13030
rect 4783 13028 4807 13030
rect 4863 13028 4887 13030
rect 4943 13028 4967 13030
rect 5023 13028 5029 13030
rect 4721 13019 5029 13028
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 1421 12540 1729 12549
rect 1421 12538 1427 12540
rect 1483 12538 1507 12540
rect 1563 12538 1587 12540
rect 1643 12538 1667 12540
rect 1723 12538 1729 12540
rect 1483 12486 1485 12538
rect 1665 12486 1667 12538
rect 1421 12484 1427 12486
rect 1483 12484 1507 12486
rect 1563 12484 1587 12486
rect 1643 12484 1667 12486
rect 1723 12484 1729 12486
rect 1421 12475 1729 12484
rect 2364 12540 2672 12549
rect 2364 12538 2370 12540
rect 2426 12538 2450 12540
rect 2506 12538 2530 12540
rect 2586 12538 2610 12540
rect 2666 12538 2672 12540
rect 2426 12486 2428 12538
rect 2608 12486 2610 12538
rect 2364 12484 2370 12486
rect 2426 12484 2450 12486
rect 2506 12484 2530 12486
rect 2586 12484 2610 12486
rect 2666 12484 2672 12486
rect 2364 12475 2672 12484
rect 3307 12540 3615 12549
rect 3307 12538 3313 12540
rect 3369 12538 3393 12540
rect 3449 12538 3473 12540
rect 3529 12538 3553 12540
rect 3609 12538 3615 12540
rect 3369 12486 3371 12538
rect 3551 12486 3553 12538
rect 3307 12484 3313 12486
rect 3369 12484 3393 12486
rect 3449 12484 3473 12486
rect 3529 12484 3553 12486
rect 3609 12484 3615 12486
rect 3307 12475 3615 12484
rect 4250 12540 4558 12549
rect 4250 12538 4256 12540
rect 4312 12538 4336 12540
rect 4392 12538 4416 12540
rect 4472 12538 4496 12540
rect 4552 12538 4558 12540
rect 4312 12486 4314 12538
rect 4494 12486 4496 12538
rect 4250 12484 4256 12486
rect 4312 12484 4336 12486
rect 4392 12484 4416 12486
rect 4472 12484 4496 12486
rect 4552 12484 4558 12486
rect 4250 12475 4558 12484
rect 1892 11996 2200 12005
rect 1892 11994 1898 11996
rect 1954 11994 1978 11996
rect 2034 11994 2058 11996
rect 2114 11994 2138 11996
rect 2194 11994 2200 11996
rect 1954 11942 1956 11994
rect 2136 11942 2138 11994
rect 1892 11940 1898 11942
rect 1954 11940 1978 11942
rect 2034 11940 2058 11942
rect 2114 11940 2138 11942
rect 2194 11940 2200 11942
rect 1892 11931 2200 11940
rect 2835 11996 3143 12005
rect 2835 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3081 11996
rect 3137 11994 3143 11996
rect 2897 11942 2899 11994
rect 3079 11942 3081 11994
rect 2835 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3081 11942
rect 3137 11940 3143 11942
rect 2835 11931 3143 11940
rect 3778 11996 4086 12005
rect 3778 11994 3784 11996
rect 3840 11994 3864 11996
rect 3920 11994 3944 11996
rect 4000 11994 4024 11996
rect 4080 11994 4086 11996
rect 3840 11942 3842 11994
rect 4022 11942 4024 11994
rect 3778 11940 3784 11942
rect 3840 11940 3864 11942
rect 3920 11940 3944 11942
rect 4000 11940 4024 11942
rect 4080 11940 4086 11942
rect 3778 11931 4086 11940
rect 4721 11996 5029 12005
rect 4721 11994 4727 11996
rect 4783 11994 4807 11996
rect 4863 11994 4887 11996
rect 4943 11994 4967 11996
rect 5023 11994 5029 11996
rect 4783 11942 4785 11994
rect 4965 11942 4967 11994
rect 4721 11940 4727 11942
rect 4783 11940 4807 11942
rect 4863 11940 4887 11942
rect 4943 11940 4967 11942
rect 5023 11940 5029 11942
rect 4721 11931 5029 11940
rect 1421 11452 1729 11461
rect 1421 11450 1427 11452
rect 1483 11450 1507 11452
rect 1563 11450 1587 11452
rect 1643 11450 1667 11452
rect 1723 11450 1729 11452
rect 1483 11398 1485 11450
rect 1665 11398 1667 11450
rect 1421 11396 1427 11398
rect 1483 11396 1507 11398
rect 1563 11396 1587 11398
rect 1643 11396 1667 11398
rect 1723 11396 1729 11398
rect 1421 11387 1729 11396
rect 2364 11452 2672 11461
rect 2364 11450 2370 11452
rect 2426 11450 2450 11452
rect 2506 11450 2530 11452
rect 2586 11450 2610 11452
rect 2666 11450 2672 11452
rect 2426 11398 2428 11450
rect 2608 11398 2610 11450
rect 2364 11396 2370 11398
rect 2426 11396 2450 11398
rect 2506 11396 2530 11398
rect 2586 11396 2610 11398
rect 2666 11396 2672 11398
rect 2364 11387 2672 11396
rect 3307 11452 3615 11461
rect 3307 11450 3313 11452
rect 3369 11450 3393 11452
rect 3449 11450 3473 11452
rect 3529 11450 3553 11452
rect 3609 11450 3615 11452
rect 3369 11398 3371 11450
rect 3551 11398 3553 11450
rect 3307 11396 3313 11398
rect 3369 11396 3393 11398
rect 3449 11396 3473 11398
rect 3529 11396 3553 11398
rect 3609 11396 3615 11398
rect 3307 11387 3615 11396
rect 4250 11452 4558 11461
rect 4250 11450 4256 11452
rect 4312 11450 4336 11452
rect 4392 11450 4416 11452
rect 4472 11450 4496 11452
rect 4552 11450 4558 11452
rect 4312 11398 4314 11450
rect 4494 11398 4496 11450
rect 4250 11396 4256 11398
rect 4312 11396 4336 11398
rect 4392 11396 4416 11398
rect 4472 11396 4496 11398
rect 4552 11396 4558 11398
rect 4250 11387 4558 11396
rect 1892 10908 2200 10917
rect 1892 10906 1898 10908
rect 1954 10906 1978 10908
rect 2034 10906 2058 10908
rect 2114 10906 2138 10908
rect 2194 10906 2200 10908
rect 1954 10854 1956 10906
rect 2136 10854 2138 10906
rect 1892 10852 1898 10854
rect 1954 10852 1978 10854
rect 2034 10852 2058 10854
rect 2114 10852 2138 10854
rect 2194 10852 2200 10854
rect 1892 10843 2200 10852
rect 2835 10908 3143 10917
rect 2835 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3081 10908
rect 3137 10906 3143 10908
rect 2897 10854 2899 10906
rect 3079 10854 3081 10906
rect 2835 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3081 10854
rect 3137 10852 3143 10854
rect 2835 10843 3143 10852
rect 3778 10908 4086 10917
rect 3778 10906 3784 10908
rect 3840 10906 3864 10908
rect 3920 10906 3944 10908
rect 4000 10906 4024 10908
rect 4080 10906 4086 10908
rect 3840 10854 3842 10906
rect 4022 10854 4024 10906
rect 3778 10852 3784 10854
rect 3840 10852 3864 10854
rect 3920 10852 3944 10854
rect 4000 10852 4024 10854
rect 4080 10852 4086 10854
rect 3778 10843 4086 10852
rect 4721 10908 5029 10917
rect 4721 10906 4727 10908
rect 4783 10906 4807 10908
rect 4863 10906 4887 10908
rect 4943 10906 4967 10908
rect 5023 10906 5029 10908
rect 4783 10854 4785 10906
rect 4965 10854 4967 10906
rect 4721 10852 4727 10854
rect 4783 10852 4807 10854
rect 4863 10852 4887 10854
rect 4943 10852 4967 10854
rect 5023 10852 5029 10854
rect 4721 10843 5029 10852
rect 1421 10364 1729 10373
rect 1421 10362 1427 10364
rect 1483 10362 1507 10364
rect 1563 10362 1587 10364
rect 1643 10362 1667 10364
rect 1723 10362 1729 10364
rect 1483 10310 1485 10362
rect 1665 10310 1667 10362
rect 1421 10308 1427 10310
rect 1483 10308 1507 10310
rect 1563 10308 1587 10310
rect 1643 10308 1667 10310
rect 1723 10308 1729 10310
rect 1421 10299 1729 10308
rect 2364 10364 2672 10373
rect 2364 10362 2370 10364
rect 2426 10362 2450 10364
rect 2506 10362 2530 10364
rect 2586 10362 2610 10364
rect 2666 10362 2672 10364
rect 2426 10310 2428 10362
rect 2608 10310 2610 10362
rect 2364 10308 2370 10310
rect 2426 10308 2450 10310
rect 2506 10308 2530 10310
rect 2586 10308 2610 10310
rect 2666 10308 2672 10310
rect 2364 10299 2672 10308
rect 3307 10364 3615 10373
rect 3307 10362 3313 10364
rect 3369 10362 3393 10364
rect 3449 10362 3473 10364
rect 3529 10362 3553 10364
rect 3609 10362 3615 10364
rect 3369 10310 3371 10362
rect 3551 10310 3553 10362
rect 3307 10308 3313 10310
rect 3369 10308 3393 10310
rect 3449 10308 3473 10310
rect 3529 10308 3553 10310
rect 3609 10308 3615 10310
rect 3307 10299 3615 10308
rect 4250 10364 4558 10373
rect 4250 10362 4256 10364
rect 4312 10362 4336 10364
rect 4392 10362 4416 10364
rect 4472 10362 4496 10364
rect 4552 10362 4558 10364
rect 4312 10310 4314 10362
rect 4494 10310 4496 10362
rect 4250 10308 4256 10310
rect 4312 10308 4336 10310
rect 4392 10308 4416 10310
rect 4472 10308 4496 10310
rect 4552 10308 4558 10310
rect 4250 10299 4558 10308
rect 4526 10160 4582 10169
rect 4526 10095 4528 10104
rect 4580 10095 4582 10104
rect 4528 10066 4580 10072
rect 1892 9820 2200 9829
rect 1892 9818 1898 9820
rect 1954 9818 1978 9820
rect 2034 9818 2058 9820
rect 2114 9818 2138 9820
rect 2194 9818 2200 9820
rect 1954 9766 1956 9818
rect 2136 9766 2138 9818
rect 1892 9764 1898 9766
rect 1954 9764 1978 9766
rect 2034 9764 2058 9766
rect 2114 9764 2138 9766
rect 2194 9764 2200 9766
rect 1892 9755 2200 9764
rect 2835 9820 3143 9829
rect 2835 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3081 9820
rect 3137 9818 3143 9820
rect 2897 9766 2899 9818
rect 3079 9766 3081 9818
rect 2835 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3081 9766
rect 3137 9764 3143 9766
rect 2835 9755 3143 9764
rect 3778 9820 4086 9829
rect 3778 9818 3784 9820
rect 3840 9818 3864 9820
rect 3920 9818 3944 9820
rect 4000 9818 4024 9820
rect 4080 9818 4086 9820
rect 3840 9766 3842 9818
rect 4022 9766 4024 9818
rect 3778 9764 3784 9766
rect 3840 9764 3864 9766
rect 3920 9764 3944 9766
rect 4000 9764 4024 9766
rect 4080 9764 4086 9766
rect 3778 9755 4086 9764
rect 4721 9820 5029 9829
rect 4721 9818 4727 9820
rect 4783 9818 4807 9820
rect 4863 9818 4887 9820
rect 4943 9818 4967 9820
rect 5023 9818 5029 9820
rect 4783 9766 4785 9818
rect 4965 9766 4967 9818
rect 4721 9764 4727 9766
rect 4783 9764 4807 9766
rect 4863 9764 4887 9766
rect 4943 9764 4967 9766
rect 5023 9764 5029 9766
rect 4721 9755 5029 9764
rect 1421 9276 1729 9285
rect 1421 9274 1427 9276
rect 1483 9274 1507 9276
rect 1563 9274 1587 9276
rect 1643 9274 1667 9276
rect 1723 9274 1729 9276
rect 1483 9222 1485 9274
rect 1665 9222 1667 9274
rect 1421 9220 1427 9222
rect 1483 9220 1507 9222
rect 1563 9220 1587 9222
rect 1643 9220 1667 9222
rect 1723 9220 1729 9222
rect 1421 9211 1729 9220
rect 2364 9276 2672 9285
rect 2364 9274 2370 9276
rect 2426 9274 2450 9276
rect 2506 9274 2530 9276
rect 2586 9274 2610 9276
rect 2666 9274 2672 9276
rect 2426 9222 2428 9274
rect 2608 9222 2610 9274
rect 2364 9220 2370 9222
rect 2426 9220 2450 9222
rect 2506 9220 2530 9222
rect 2586 9220 2610 9222
rect 2666 9220 2672 9222
rect 2364 9211 2672 9220
rect 3307 9276 3615 9285
rect 3307 9274 3313 9276
rect 3369 9274 3393 9276
rect 3449 9274 3473 9276
rect 3529 9274 3553 9276
rect 3609 9274 3615 9276
rect 3369 9222 3371 9274
rect 3551 9222 3553 9274
rect 3307 9220 3313 9222
rect 3369 9220 3393 9222
rect 3449 9220 3473 9222
rect 3529 9220 3553 9222
rect 3609 9220 3615 9222
rect 3307 9211 3615 9220
rect 4250 9276 4558 9285
rect 4250 9274 4256 9276
rect 4312 9274 4336 9276
rect 4392 9274 4416 9276
rect 4472 9274 4496 9276
rect 4552 9274 4558 9276
rect 4312 9222 4314 9274
rect 4494 9222 4496 9274
rect 4250 9220 4256 9222
rect 4312 9220 4336 9222
rect 4392 9220 4416 9222
rect 4472 9220 4496 9222
rect 4552 9220 4558 9222
rect 4250 9211 4558 9220
rect 1892 8732 2200 8741
rect 1892 8730 1898 8732
rect 1954 8730 1978 8732
rect 2034 8730 2058 8732
rect 2114 8730 2138 8732
rect 2194 8730 2200 8732
rect 1954 8678 1956 8730
rect 2136 8678 2138 8730
rect 1892 8676 1898 8678
rect 1954 8676 1978 8678
rect 2034 8676 2058 8678
rect 2114 8676 2138 8678
rect 2194 8676 2200 8678
rect 1892 8667 2200 8676
rect 2835 8732 3143 8741
rect 2835 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3081 8732
rect 3137 8730 3143 8732
rect 2897 8678 2899 8730
rect 3079 8678 3081 8730
rect 2835 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3081 8678
rect 3137 8676 3143 8678
rect 2835 8667 3143 8676
rect 3778 8732 4086 8741
rect 3778 8730 3784 8732
rect 3840 8730 3864 8732
rect 3920 8730 3944 8732
rect 4000 8730 4024 8732
rect 4080 8730 4086 8732
rect 3840 8678 3842 8730
rect 4022 8678 4024 8730
rect 3778 8676 3784 8678
rect 3840 8676 3864 8678
rect 3920 8676 3944 8678
rect 4000 8676 4024 8678
rect 4080 8676 4086 8678
rect 3778 8667 4086 8676
rect 4721 8732 5029 8741
rect 4721 8730 4727 8732
rect 4783 8730 4807 8732
rect 4863 8730 4887 8732
rect 4943 8730 4967 8732
rect 5023 8730 5029 8732
rect 4783 8678 4785 8730
rect 4965 8678 4967 8730
rect 4721 8676 4727 8678
rect 4783 8676 4807 8678
rect 4863 8676 4887 8678
rect 4943 8676 4967 8678
rect 5023 8676 5029 8678
rect 4721 8667 5029 8676
rect 1421 8188 1729 8197
rect 1421 8186 1427 8188
rect 1483 8186 1507 8188
rect 1563 8186 1587 8188
rect 1643 8186 1667 8188
rect 1723 8186 1729 8188
rect 1483 8134 1485 8186
rect 1665 8134 1667 8186
rect 1421 8132 1427 8134
rect 1483 8132 1507 8134
rect 1563 8132 1587 8134
rect 1643 8132 1667 8134
rect 1723 8132 1729 8134
rect 1421 8123 1729 8132
rect 2364 8188 2672 8197
rect 2364 8186 2370 8188
rect 2426 8186 2450 8188
rect 2506 8186 2530 8188
rect 2586 8186 2610 8188
rect 2666 8186 2672 8188
rect 2426 8134 2428 8186
rect 2608 8134 2610 8186
rect 2364 8132 2370 8134
rect 2426 8132 2450 8134
rect 2506 8132 2530 8134
rect 2586 8132 2610 8134
rect 2666 8132 2672 8134
rect 2364 8123 2672 8132
rect 3307 8188 3615 8197
rect 3307 8186 3313 8188
rect 3369 8186 3393 8188
rect 3449 8186 3473 8188
rect 3529 8186 3553 8188
rect 3609 8186 3615 8188
rect 3369 8134 3371 8186
rect 3551 8134 3553 8186
rect 3307 8132 3313 8134
rect 3369 8132 3393 8134
rect 3449 8132 3473 8134
rect 3529 8132 3553 8134
rect 3609 8132 3615 8134
rect 3307 8123 3615 8132
rect 4250 8188 4558 8197
rect 4250 8186 4256 8188
rect 4312 8186 4336 8188
rect 4392 8186 4416 8188
rect 4472 8186 4496 8188
rect 4552 8186 4558 8188
rect 4312 8134 4314 8186
rect 4494 8134 4496 8186
rect 4250 8132 4256 8134
rect 4312 8132 4336 8134
rect 4392 8132 4416 8134
rect 4472 8132 4496 8134
rect 4552 8132 4558 8134
rect 4250 8123 4558 8132
rect 1766 7984 1822 7993
rect 1766 7919 1822 7928
rect 1421 7100 1729 7109
rect 1421 7098 1427 7100
rect 1483 7098 1507 7100
rect 1563 7098 1587 7100
rect 1643 7098 1667 7100
rect 1723 7098 1729 7100
rect 1483 7046 1485 7098
rect 1665 7046 1667 7098
rect 1421 7044 1427 7046
rect 1483 7044 1507 7046
rect 1563 7044 1587 7046
rect 1643 7044 1667 7046
rect 1723 7044 1729 7046
rect 1421 7035 1729 7044
rect 1780 6322 1808 7919
rect 1892 7644 2200 7653
rect 1892 7642 1898 7644
rect 1954 7642 1978 7644
rect 2034 7642 2058 7644
rect 2114 7642 2138 7644
rect 2194 7642 2200 7644
rect 1954 7590 1956 7642
rect 2136 7590 2138 7642
rect 1892 7588 1898 7590
rect 1954 7588 1978 7590
rect 2034 7588 2058 7590
rect 2114 7588 2138 7590
rect 2194 7588 2200 7590
rect 1892 7579 2200 7588
rect 2835 7644 3143 7653
rect 2835 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3081 7644
rect 3137 7642 3143 7644
rect 2897 7590 2899 7642
rect 3079 7590 3081 7642
rect 2835 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3081 7590
rect 3137 7588 3143 7590
rect 2835 7579 3143 7588
rect 3778 7644 4086 7653
rect 3778 7642 3784 7644
rect 3840 7642 3864 7644
rect 3920 7642 3944 7644
rect 4000 7642 4024 7644
rect 4080 7642 4086 7644
rect 3840 7590 3842 7642
rect 4022 7590 4024 7642
rect 3778 7588 3784 7590
rect 3840 7588 3864 7590
rect 3920 7588 3944 7590
rect 4000 7588 4024 7590
rect 4080 7588 4086 7590
rect 3778 7579 4086 7588
rect 4721 7644 5029 7653
rect 4721 7642 4727 7644
rect 4783 7642 4807 7644
rect 4863 7642 4887 7644
rect 4943 7642 4967 7644
rect 5023 7642 5029 7644
rect 4783 7590 4785 7642
rect 4965 7590 4967 7642
rect 4721 7588 4727 7590
rect 4783 7588 4807 7590
rect 4863 7588 4887 7590
rect 4943 7588 4967 7590
rect 5023 7588 5029 7590
rect 4721 7579 5029 7588
rect 2364 7100 2672 7109
rect 2364 7098 2370 7100
rect 2426 7098 2450 7100
rect 2506 7098 2530 7100
rect 2586 7098 2610 7100
rect 2666 7098 2672 7100
rect 2426 7046 2428 7098
rect 2608 7046 2610 7098
rect 2364 7044 2370 7046
rect 2426 7044 2450 7046
rect 2506 7044 2530 7046
rect 2586 7044 2610 7046
rect 2666 7044 2672 7046
rect 2364 7035 2672 7044
rect 3307 7100 3615 7109
rect 3307 7098 3313 7100
rect 3369 7098 3393 7100
rect 3449 7098 3473 7100
rect 3529 7098 3553 7100
rect 3609 7098 3615 7100
rect 3369 7046 3371 7098
rect 3551 7046 3553 7098
rect 3307 7044 3313 7046
rect 3369 7044 3393 7046
rect 3449 7044 3473 7046
rect 3529 7044 3553 7046
rect 3609 7044 3615 7046
rect 3307 7035 3615 7044
rect 4250 7100 4558 7109
rect 4250 7098 4256 7100
rect 4312 7098 4336 7100
rect 4392 7098 4416 7100
rect 4472 7098 4496 7100
rect 4552 7098 4558 7100
rect 4312 7046 4314 7098
rect 4494 7046 4496 7098
rect 4250 7044 4256 7046
rect 4312 7044 4336 7046
rect 4392 7044 4416 7046
rect 4472 7044 4496 7046
rect 4552 7044 4558 7046
rect 4250 7035 4558 7044
rect 1892 6556 2200 6565
rect 1892 6554 1898 6556
rect 1954 6554 1978 6556
rect 2034 6554 2058 6556
rect 2114 6554 2138 6556
rect 2194 6554 2200 6556
rect 1954 6502 1956 6554
rect 2136 6502 2138 6554
rect 1892 6500 1898 6502
rect 1954 6500 1978 6502
rect 2034 6500 2058 6502
rect 2114 6500 2138 6502
rect 2194 6500 2200 6502
rect 1892 6491 2200 6500
rect 2835 6556 3143 6565
rect 2835 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3081 6556
rect 3137 6554 3143 6556
rect 2897 6502 2899 6554
rect 3079 6502 3081 6554
rect 2835 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3081 6502
rect 3137 6500 3143 6502
rect 2835 6491 3143 6500
rect 3778 6556 4086 6565
rect 3778 6554 3784 6556
rect 3840 6554 3864 6556
rect 3920 6554 3944 6556
rect 4000 6554 4024 6556
rect 4080 6554 4086 6556
rect 3840 6502 3842 6554
rect 4022 6502 4024 6554
rect 3778 6500 3784 6502
rect 3840 6500 3864 6502
rect 3920 6500 3944 6502
rect 4000 6500 4024 6502
rect 4080 6500 4086 6502
rect 3778 6491 4086 6500
rect 4721 6556 5029 6565
rect 4721 6554 4727 6556
rect 4783 6554 4807 6556
rect 4863 6554 4887 6556
rect 4943 6554 4967 6556
rect 5023 6554 5029 6556
rect 4783 6502 4785 6554
rect 4965 6502 4967 6554
rect 4721 6500 4727 6502
rect 4783 6500 4807 6502
rect 4863 6500 4887 6502
rect 4943 6500 4967 6502
rect 5023 6500 5029 6502
rect 4721 6491 5029 6500
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 1421 6012 1729 6021
rect 1421 6010 1427 6012
rect 1483 6010 1507 6012
rect 1563 6010 1587 6012
rect 1643 6010 1667 6012
rect 1723 6010 1729 6012
rect 1483 5958 1485 6010
rect 1665 5958 1667 6010
rect 1421 5956 1427 5958
rect 1483 5956 1507 5958
rect 1563 5956 1587 5958
rect 1643 5956 1667 5958
rect 1723 5956 1729 5958
rect 1421 5947 1729 5956
rect 2364 6012 2672 6021
rect 2364 6010 2370 6012
rect 2426 6010 2450 6012
rect 2506 6010 2530 6012
rect 2586 6010 2610 6012
rect 2666 6010 2672 6012
rect 2426 5958 2428 6010
rect 2608 5958 2610 6010
rect 2364 5956 2370 5958
rect 2426 5956 2450 5958
rect 2506 5956 2530 5958
rect 2586 5956 2610 5958
rect 2666 5956 2672 5958
rect 2364 5947 2672 5956
rect 3307 6012 3615 6021
rect 3307 6010 3313 6012
rect 3369 6010 3393 6012
rect 3449 6010 3473 6012
rect 3529 6010 3553 6012
rect 3609 6010 3615 6012
rect 3369 5958 3371 6010
rect 3551 5958 3553 6010
rect 3307 5956 3313 5958
rect 3369 5956 3393 5958
rect 3449 5956 3473 5958
rect 3529 5956 3553 5958
rect 3609 5956 3615 5958
rect 3307 5947 3615 5956
rect 1892 5468 2200 5477
rect 1892 5466 1898 5468
rect 1954 5466 1978 5468
rect 2034 5466 2058 5468
rect 2114 5466 2138 5468
rect 2194 5466 2200 5468
rect 1954 5414 1956 5466
rect 2136 5414 2138 5466
rect 1892 5412 1898 5414
rect 1954 5412 1978 5414
rect 2034 5412 2058 5414
rect 2114 5412 2138 5414
rect 2194 5412 2200 5414
rect 1892 5403 2200 5412
rect 2835 5468 3143 5477
rect 2835 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3081 5468
rect 3137 5466 3143 5468
rect 2897 5414 2899 5466
rect 3079 5414 3081 5466
rect 2835 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3081 5414
rect 3137 5412 3143 5414
rect 2835 5403 3143 5412
rect 3778 5468 4086 5477
rect 3778 5466 3784 5468
rect 3840 5466 3864 5468
rect 3920 5466 3944 5468
rect 4000 5466 4024 5468
rect 4080 5466 4086 5468
rect 3840 5414 3842 5466
rect 4022 5414 4024 5466
rect 3778 5412 3784 5414
rect 3840 5412 3864 5414
rect 3920 5412 3944 5414
rect 4000 5412 4024 5414
rect 4080 5412 4086 5414
rect 3778 5403 4086 5412
rect 1421 4924 1729 4933
rect 1421 4922 1427 4924
rect 1483 4922 1507 4924
rect 1563 4922 1587 4924
rect 1643 4922 1667 4924
rect 1723 4922 1729 4924
rect 1483 4870 1485 4922
rect 1665 4870 1667 4922
rect 1421 4868 1427 4870
rect 1483 4868 1507 4870
rect 1563 4868 1587 4870
rect 1643 4868 1667 4870
rect 1723 4868 1729 4870
rect 1421 4859 1729 4868
rect 2364 4924 2672 4933
rect 2364 4922 2370 4924
rect 2426 4922 2450 4924
rect 2506 4922 2530 4924
rect 2586 4922 2610 4924
rect 2666 4922 2672 4924
rect 2426 4870 2428 4922
rect 2608 4870 2610 4922
rect 2364 4868 2370 4870
rect 2426 4868 2450 4870
rect 2506 4868 2530 4870
rect 2586 4868 2610 4870
rect 2666 4868 2672 4870
rect 2364 4859 2672 4868
rect 3307 4924 3615 4933
rect 3307 4922 3313 4924
rect 3369 4922 3393 4924
rect 3449 4922 3473 4924
rect 3529 4922 3553 4924
rect 3609 4922 3615 4924
rect 3369 4870 3371 4922
rect 3551 4870 3553 4922
rect 3307 4868 3313 4870
rect 3369 4868 3393 4870
rect 3449 4868 3473 4870
rect 3529 4868 3553 4870
rect 3609 4868 3615 4870
rect 3307 4859 3615 4868
rect 1892 4380 2200 4389
rect 1892 4378 1898 4380
rect 1954 4378 1978 4380
rect 2034 4378 2058 4380
rect 2114 4378 2138 4380
rect 2194 4378 2200 4380
rect 1954 4326 1956 4378
rect 2136 4326 2138 4378
rect 1892 4324 1898 4326
rect 1954 4324 1978 4326
rect 2034 4324 2058 4326
rect 2114 4324 2138 4326
rect 2194 4324 2200 4326
rect 1892 4315 2200 4324
rect 2835 4380 3143 4389
rect 2835 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3081 4380
rect 3137 4378 3143 4380
rect 2897 4326 2899 4378
rect 3079 4326 3081 4378
rect 2835 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3081 4326
rect 3137 4324 3143 4326
rect 2835 4315 3143 4324
rect 3778 4380 4086 4389
rect 3778 4378 3784 4380
rect 3840 4378 3864 4380
rect 3920 4378 3944 4380
rect 4000 4378 4024 4380
rect 4080 4378 4086 4380
rect 3840 4326 3842 4378
rect 4022 4326 4024 4378
rect 3778 4324 3784 4326
rect 3840 4324 3864 4326
rect 3920 4324 3944 4326
rect 4000 4324 4024 4326
rect 4080 4324 4086 4326
rect 3778 4315 4086 4324
rect 1421 3836 1729 3845
rect 1421 3834 1427 3836
rect 1483 3834 1507 3836
rect 1563 3834 1587 3836
rect 1643 3834 1667 3836
rect 1723 3834 1729 3836
rect 1483 3782 1485 3834
rect 1665 3782 1667 3834
rect 1421 3780 1427 3782
rect 1483 3780 1507 3782
rect 1563 3780 1587 3782
rect 1643 3780 1667 3782
rect 1723 3780 1729 3782
rect 1421 3771 1729 3780
rect 2364 3836 2672 3845
rect 2364 3834 2370 3836
rect 2426 3834 2450 3836
rect 2506 3834 2530 3836
rect 2586 3834 2610 3836
rect 2666 3834 2672 3836
rect 2426 3782 2428 3834
rect 2608 3782 2610 3834
rect 2364 3780 2370 3782
rect 2426 3780 2450 3782
rect 2506 3780 2530 3782
rect 2586 3780 2610 3782
rect 2666 3780 2672 3782
rect 2364 3771 2672 3780
rect 3307 3836 3615 3845
rect 3307 3834 3313 3836
rect 3369 3834 3393 3836
rect 3449 3834 3473 3836
rect 3529 3834 3553 3836
rect 3609 3834 3615 3836
rect 3369 3782 3371 3834
rect 3551 3782 3553 3834
rect 3307 3780 3313 3782
rect 3369 3780 3393 3782
rect 3449 3780 3473 3782
rect 3529 3780 3553 3782
rect 3609 3780 3615 3782
rect 3307 3771 3615 3780
rect 1892 3292 2200 3301
rect 1892 3290 1898 3292
rect 1954 3290 1978 3292
rect 2034 3290 2058 3292
rect 2114 3290 2138 3292
rect 2194 3290 2200 3292
rect 1954 3238 1956 3290
rect 2136 3238 2138 3290
rect 1892 3236 1898 3238
rect 1954 3236 1978 3238
rect 2034 3236 2058 3238
rect 2114 3236 2138 3238
rect 2194 3236 2200 3238
rect 1892 3227 2200 3236
rect 2835 3292 3143 3301
rect 2835 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3081 3292
rect 3137 3290 3143 3292
rect 2897 3238 2899 3290
rect 3079 3238 3081 3290
rect 2835 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3081 3238
rect 3137 3236 3143 3238
rect 2835 3227 3143 3236
rect 3778 3292 4086 3301
rect 3778 3290 3784 3292
rect 3840 3290 3864 3292
rect 3920 3290 3944 3292
rect 4000 3290 4024 3292
rect 4080 3290 4086 3292
rect 3840 3238 3842 3290
rect 4022 3238 4024 3290
rect 3778 3236 3784 3238
rect 3840 3236 3864 3238
rect 3920 3236 3944 3238
rect 4000 3236 4024 3238
rect 4080 3236 4086 3238
rect 3778 3227 4086 3236
rect 1421 2748 1729 2757
rect 1421 2746 1427 2748
rect 1483 2746 1507 2748
rect 1563 2746 1587 2748
rect 1643 2746 1667 2748
rect 1723 2746 1729 2748
rect 1483 2694 1485 2746
rect 1665 2694 1667 2746
rect 1421 2692 1427 2694
rect 1483 2692 1507 2694
rect 1563 2692 1587 2694
rect 1643 2692 1667 2694
rect 1723 2692 1729 2694
rect 1421 2683 1729 2692
rect 2364 2748 2672 2757
rect 2364 2746 2370 2748
rect 2426 2746 2450 2748
rect 2506 2746 2530 2748
rect 2586 2746 2610 2748
rect 2666 2746 2672 2748
rect 2426 2694 2428 2746
rect 2608 2694 2610 2746
rect 2364 2692 2370 2694
rect 2426 2692 2450 2694
rect 2506 2692 2530 2694
rect 2586 2692 2610 2694
rect 2666 2692 2672 2694
rect 2364 2683 2672 2692
rect 3307 2748 3615 2757
rect 3307 2746 3313 2748
rect 3369 2746 3393 2748
rect 3449 2746 3473 2748
rect 3529 2746 3553 2748
rect 3609 2746 3615 2748
rect 3369 2694 3371 2746
rect 3551 2694 3553 2746
rect 3307 2692 3313 2694
rect 3369 2692 3393 2694
rect 3449 2692 3473 2694
rect 3529 2692 3553 2694
rect 3609 2692 3615 2694
rect 3307 2683 3615 2692
rect 4172 2650 4200 6258
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4802 6080 4858 6089
rect 4250 6012 4558 6021
rect 4250 6010 4256 6012
rect 4312 6010 4336 6012
rect 4392 6010 4416 6012
rect 4472 6010 4496 6012
rect 4552 6010 4558 6012
rect 4312 5958 4314 6010
rect 4494 5958 4496 6010
rect 4250 5956 4256 5958
rect 4312 5956 4336 5958
rect 4392 5956 4416 5958
rect 4472 5956 4496 5958
rect 4552 5956 4558 5958
rect 4250 5947 4558 5956
rect 4632 5710 4660 6054
rect 4802 6015 4858 6024
rect 4816 5914 4844 6015
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4721 5468 5029 5477
rect 4721 5466 4727 5468
rect 4783 5466 4807 5468
rect 4863 5466 4887 5468
rect 4943 5466 4967 5468
rect 5023 5466 5029 5468
rect 4783 5414 4785 5466
rect 4965 5414 4967 5466
rect 4721 5412 4727 5414
rect 4783 5412 4807 5414
rect 4863 5412 4887 5414
rect 4943 5412 4967 5414
rect 5023 5412 5029 5414
rect 4721 5403 5029 5412
rect 4250 4924 4558 4933
rect 4250 4922 4256 4924
rect 4312 4922 4336 4924
rect 4392 4922 4416 4924
rect 4472 4922 4496 4924
rect 4552 4922 4558 4924
rect 4312 4870 4314 4922
rect 4494 4870 4496 4922
rect 4250 4868 4256 4870
rect 4312 4868 4336 4870
rect 4392 4868 4416 4870
rect 4472 4868 4496 4870
rect 4552 4868 4558 4870
rect 4250 4859 4558 4868
rect 4721 4380 5029 4389
rect 4721 4378 4727 4380
rect 4783 4378 4807 4380
rect 4863 4378 4887 4380
rect 4943 4378 4967 4380
rect 5023 4378 5029 4380
rect 4783 4326 4785 4378
rect 4965 4326 4967 4378
rect 4721 4324 4727 4326
rect 4783 4324 4807 4326
rect 4863 4324 4887 4326
rect 4943 4324 4967 4326
rect 5023 4324 5029 4326
rect 4721 4315 5029 4324
rect 4250 3836 4558 3845
rect 4250 3834 4256 3836
rect 4312 3834 4336 3836
rect 4392 3834 4416 3836
rect 4472 3834 4496 3836
rect 4552 3834 4558 3836
rect 4312 3782 4314 3834
rect 4494 3782 4496 3834
rect 4250 3780 4256 3782
rect 4312 3780 4336 3782
rect 4392 3780 4416 3782
rect 4472 3780 4496 3782
rect 4552 3780 4558 3782
rect 4250 3771 4558 3780
rect 4721 3292 5029 3301
rect 4721 3290 4727 3292
rect 4783 3290 4807 3292
rect 4863 3290 4887 3292
rect 4943 3290 4967 3292
rect 5023 3290 5029 3292
rect 4783 3238 4785 3290
rect 4965 3238 4967 3290
rect 4721 3236 4727 3238
rect 4783 3236 4807 3238
rect 4863 3236 4887 3238
rect 4943 3236 4967 3238
rect 5023 3236 5029 3238
rect 4721 3227 5029 3236
rect 4250 2748 4558 2757
rect 4250 2746 4256 2748
rect 4312 2746 4336 2748
rect 4392 2746 4416 2748
rect 4472 2746 4496 2748
rect 4552 2746 4558 2748
rect 4312 2694 4314 2746
rect 4494 2694 4496 2746
rect 4250 2692 4256 2694
rect 4312 2692 4336 2694
rect 4392 2692 4416 2694
rect 4472 2692 4496 2694
rect 4552 2692 4558 2694
rect 4250 2683 4558 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4894 2544 4950 2553
rect 4894 2479 4896 2488
rect 4948 2479 4950 2488
rect 4896 2450 4948 2456
rect 1892 2204 2200 2213
rect 1892 2202 1898 2204
rect 1954 2202 1978 2204
rect 2034 2202 2058 2204
rect 2114 2202 2138 2204
rect 2194 2202 2200 2204
rect 1954 2150 1956 2202
rect 2136 2150 2138 2202
rect 1892 2148 1898 2150
rect 1954 2148 1978 2150
rect 2034 2148 2058 2150
rect 2114 2148 2138 2150
rect 2194 2148 2200 2150
rect 1892 2139 2200 2148
rect 2835 2204 3143 2213
rect 2835 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3081 2204
rect 3137 2202 3143 2204
rect 2897 2150 2899 2202
rect 3079 2150 3081 2202
rect 2835 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3081 2150
rect 3137 2148 3143 2150
rect 2835 2139 3143 2148
rect 3778 2204 4086 2213
rect 3778 2202 3784 2204
rect 3840 2202 3864 2204
rect 3920 2202 3944 2204
rect 4000 2202 4024 2204
rect 4080 2202 4086 2204
rect 3840 2150 3842 2202
rect 4022 2150 4024 2202
rect 3778 2148 3784 2150
rect 3840 2148 3864 2150
rect 3920 2148 3944 2150
rect 4000 2148 4024 2150
rect 4080 2148 4086 2150
rect 3778 2139 4086 2148
rect 4721 2204 5029 2213
rect 4721 2202 4727 2204
rect 4783 2202 4807 2204
rect 4863 2202 4887 2204
rect 4943 2202 4967 2204
rect 5023 2202 5029 2204
rect 4783 2150 4785 2202
rect 4965 2150 4967 2202
rect 4721 2148 4727 2150
rect 4783 2148 4807 2150
rect 4863 2148 4887 2150
rect 4943 2148 4967 2150
rect 5023 2148 5029 2150
rect 4721 2139 5029 2148
<< via2 >>
rect 4894 13640 4950 13696
rect 1427 13626 1483 13628
rect 1507 13626 1563 13628
rect 1587 13626 1643 13628
rect 1667 13626 1723 13628
rect 1427 13574 1473 13626
rect 1473 13574 1483 13626
rect 1507 13574 1537 13626
rect 1537 13574 1549 13626
rect 1549 13574 1563 13626
rect 1587 13574 1601 13626
rect 1601 13574 1613 13626
rect 1613 13574 1643 13626
rect 1667 13574 1677 13626
rect 1677 13574 1723 13626
rect 1427 13572 1483 13574
rect 1507 13572 1563 13574
rect 1587 13572 1643 13574
rect 1667 13572 1723 13574
rect 2370 13626 2426 13628
rect 2450 13626 2506 13628
rect 2530 13626 2586 13628
rect 2610 13626 2666 13628
rect 2370 13574 2416 13626
rect 2416 13574 2426 13626
rect 2450 13574 2480 13626
rect 2480 13574 2492 13626
rect 2492 13574 2506 13626
rect 2530 13574 2544 13626
rect 2544 13574 2556 13626
rect 2556 13574 2586 13626
rect 2610 13574 2620 13626
rect 2620 13574 2666 13626
rect 2370 13572 2426 13574
rect 2450 13572 2506 13574
rect 2530 13572 2586 13574
rect 2610 13572 2666 13574
rect 3313 13626 3369 13628
rect 3393 13626 3449 13628
rect 3473 13626 3529 13628
rect 3553 13626 3609 13628
rect 3313 13574 3359 13626
rect 3359 13574 3369 13626
rect 3393 13574 3423 13626
rect 3423 13574 3435 13626
rect 3435 13574 3449 13626
rect 3473 13574 3487 13626
rect 3487 13574 3499 13626
rect 3499 13574 3529 13626
rect 3553 13574 3563 13626
rect 3563 13574 3609 13626
rect 3313 13572 3369 13574
rect 3393 13572 3449 13574
rect 3473 13572 3529 13574
rect 3553 13572 3609 13574
rect 4256 13626 4312 13628
rect 4336 13626 4392 13628
rect 4416 13626 4472 13628
rect 4496 13626 4552 13628
rect 4256 13574 4302 13626
rect 4302 13574 4312 13626
rect 4336 13574 4366 13626
rect 4366 13574 4378 13626
rect 4378 13574 4392 13626
rect 4416 13574 4430 13626
rect 4430 13574 4442 13626
rect 4442 13574 4472 13626
rect 4496 13574 4506 13626
rect 4506 13574 4552 13626
rect 4256 13572 4312 13574
rect 4336 13572 4392 13574
rect 4416 13572 4472 13574
rect 4496 13572 4552 13574
rect 1398 13096 1454 13152
rect 1898 13082 1954 13084
rect 1978 13082 2034 13084
rect 2058 13082 2114 13084
rect 2138 13082 2194 13084
rect 1898 13030 1944 13082
rect 1944 13030 1954 13082
rect 1978 13030 2008 13082
rect 2008 13030 2020 13082
rect 2020 13030 2034 13082
rect 2058 13030 2072 13082
rect 2072 13030 2084 13082
rect 2084 13030 2114 13082
rect 2138 13030 2148 13082
rect 2148 13030 2194 13082
rect 1898 13028 1954 13030
rect 1978 13028 2034 13030
rect 2058 13028 2114 13030
rect 2138 13028 2194 13030
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 3081 13082 3137 13084
rect 2841 13030 2887 13082
rect 2887 13030 2897 13082
rect 2921 13030 2951 13082
rect 2951 13030 2963 13082
rect 2963 13030 2977 13082
rect 3001 13030 3015 13082
rect 3015 13030 3027 13082
rect 3027 13030 3057 13082
rect 3081 13030 3091 13082
rect 3091 13030 3137 13082
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 3081 13028 3137 13030
rect 3784 13082 3840 13084
rect 3864 13082 3920 13084
rect 3944 13082 4000 13084
rect 4024 13082 4080 13084
rect 3784 13030 3830 13082
rect 3830 13030 3840 13082
rect 3864 13030 3894 13082
rect 3894 13030 3906 13082
rect 3906 13030 3920 13082
rect 3944 13030 3958 13082
rect 3958 13030 3970 13082
rect 3970 13030 4000 13082
rect 4024 13030 4034 13082
rect 4034 13030 4080 13082
rect 3784 13028 3840 13030
rect 3864 13028 3920 13030
rect 3944 13028 4000 13030
rect 4024 13028 4080 13030
rect 4727 13082 4783 13084
rect 4807 13082 4863 13084
rect 4887 13082 4943 13084
rect 4967 13082 5023 13084
rect 4727 13030 4773 13082
rect 4773 13030 4783 13082
rect 4807 13030 4837 13082
rect 4837 13030 4849 13082
rect 4849 13030 4863 13082
rect 4887 13030 4901 13082
rect 4901 13030 4913 13082
rect 4913 13030 4943 13082
rect 4967 13030 4977 13082
rect 4977 13030 5023 13082
rect 4727 13028 4783 13030
rect 4807 13028 4863 13030
rect 4887 13028 4943 13030
rect 4967 13028 5023 13030
rect 1427 12538 1483 12540
rect 1507 12538 1563 12540
rect 1587 12538 1643 12540
rect 1667 12538 1723 12540
rect 1427 12486 1473 12538
rect 1473 12486 1483 12538
rect 1507 12486 1537 12538
rect 1537 12486 1549 12538
rect 1549 12486 1563 12538
rect 1587 12486 1601 12538
rect 1601 12486 1613 12538
rect 1613 12486 1643 12538
rect 1667 12486 1677 12538
rect 1677 12486 1723 12538
rect 1427 12484 1483 12486
rect 1507 12484 1563 12486
rect 1587 12484 1643 12486
rect 1667 12484 1723 12486
rect 2370 12538 2426 12540
rect 2450 12538 2506 12540
rect 2530 12538 2586 12540
rect 2610 12538 2666 12540
rect 2370 12486 2416 12538
rect 2416 12486 2426 12538
rect 2450 12486 2480 12538
rect 2480 12486 2492 12538
rect 2492 12486 2506 12538
rect 2530 12486 2544 12538
rect 2544 12486 2556 12538
rect 2556 12486 2586 12538
rect 2610 12486 2620 12538
rect 2620 12486 2666 12538
rect 2370 12484 2426 12486
rect 2450 12484 2506 12486
rect 2530 12484 2586 12486
rect 2610 12484 2666 12486
rect 3313 12538 3369 12540
rect 3393 12538 3449 12540
rect 3473 12538 3529 12540
rect 3553 12538 3609 12540
rect 3313 12486 3359 12538
rect 3359 12486 3369 12538
rect 3393 12486 3423 12538
rect 3423 12486 3435 12538
rect 3435 12486 3449 12538
rect 3473 12486 3487 12538
rect 3487 12486 3499 12538
rect 3499 12486 3529 12538
rect 3553 12486 3563 12538
rect 3563 12486 3609 12538
rect 3313 12484 3369 12486
rect 3393 12484 3449 12486
rect 3473 12484 3529 12486
rect 3553 12484 3609 12486
rect 4256 12538 4312 12540
rect 4336 12538 4392 12540
rect 4416 12538 4472 12540
rect 4496 12538 4552 12540
rect 4256 12486 4302 12538
rect 4302 12486 4312 12538
rect 4336 12486 4366 12538
rect 4366 12486 4378 12538
rect 4378 12486 4392 12538
rect 4416 12486 4430 12538
rect 4430 12486 4442 12538
rect 4442 12486 4472 12538
rect 4496 12486 4506 12538
rect 4506 12486 4552 12538
rect 4256 12484 4312 12486
rect 4336 12484 4392 12486
rect 4416 12484 4472 12486
rect 4496 12484 4552 12486
rect 1898 11994 1954 11996
rect 1978 11994 2034 11996
rect 2058 11994 2114 11996
rect 2138 11994 2194 11996
rect 1898 11942 1944 11994
rect 1944 11942 1954 11994
rect 1978 11942 2008 11994
rect 2008 11942 2020 11994
rect 2020 11942 2034 11994
rect 2058 11942 2072 11994
rect 2072 11942 2084 11994
rect 2084 11942 2114 11994
rect 2138 11942 2148 11994
rect 2148 11942 2194 11994
rect 1898 11940 1954 11942
rect 1978 11940 2034 11942
rect 2058 11940 2114 11942
rect 2138 11940 2194 11942
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 3081 11994 3137 11996
rect 2841 11942 2887 11994
rect 2887 11942 2897 11994
rect 2921 11942 2951 11994
rect 2951 11942 2963 11994
rect 2963 11942 2977 11994
rect 3001 11942 3015 11994
rect 3015 11942 3027 11994
rect 3027 11942 3057 11994
rect 3081 11942 3091 11994
rect 3091 11942 3137 11994
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 3081 11940 3137 11942
rect 3784 11994 3840 11996
rect 3864 11994 3920 11996
rect 3944 11994 4000 11996
rect 4024 11994 4080 11996
rect 3784 11942 3830 11994
rect 3830 11942 3840 11994
rect 3864 11942 3894 11994
rect 3894 11942 3906 11994
rect 3906 11942 3920 11994
rect 3944 11942 3958 11994
rect 3958 11942 3970 11994
rect 3970 11942 4000 11994
rect 4024 11942 4034 11994
rect 4034 11942 4080 11994
rect 3784 11940 3840 11942
rect 3864 11940 3920 11942
rect 3944 11940 4000 11942
rect 4024 11940 4080 11942
rect 4727 11994 4783 11996
rect 4807 11994 4863 11996
rect 4887 11994 4943 11996
rect 4967 11994 5023 11996
rect 4727 11942 4773 11994
rect 4773 11942 4783 11994
rect 4807 11942 4837 11994
rect 4837 11942 4849 11994
rect 4849 11942 4863 11994
rect 4887 11942 4901 11994
rect 4901 11942 4913 11994
rect 4913 11942 4943 11994
rect 4967 11942 4977 11994
rect 4977 11942 5023 11994
rect 4727 11940 4783 11942
rect 4807 11940 4863 11942
rect 4887 11940 4943 11942
rect 4967 11940 5023 11942
rect 1427 11450 1483 11452
rect 1507 11450 1563 11452
rect 1587 11450 1643 11452
rect 1667 11450 1723 11452
rect 1427 11398 1473 11450
rect 1473 11398 1483 11450
rect 1507 11398 1537 11450
rect 1537 11398 1549 11450
rect 1549 11398 1563 11450
rect 1587 11398 1601 11450
rect 1601 11398 1613 11450
rect 1613 11398 1643 11450
rect 1667 11398 1677 11450
rect 1677 11398 1723 11450
rect 1427 11396 1483 11398
rect 1507 11396 1563 11398
rect 1587 11396 1643 11398
rect 1667 11396 1723 11398
rect 2370 11450 2426 11452
rect 2450 11450 2506 11452
rect 2530 11450 2586 11452
rect 2610 11450 2666 11452
rect 2370 11398 2416 11450
rect 2416 11398 2426 11450
rect 2450 11398 2480 11450
rect 2480 11398 2492 11450
rect 2492 11398 2506 11450
rect 2530 11398 2544 11450
rect 2544 11398 2556 11450
rect 2556 11398 2586 11450
rect 2610 11398 2620 11450
rect 2620 11398 2666 11450
rect 2370 11396 2426 11398
rect 2450 11396 2506 11398
rect 2530 11396 2586 11398
rect 2610 11396 2666 11398
rect 3313 11450 3369 11452
rect 3393 11450 3449 11452
rect 3473 11450 3529 11452
rect 3553 11450 3609 11452
rect 3313 11398 3359 11450
rect 3359 11398 3369 11450
rect 3393 11398 3423 11450
rect 3423 11398 3435 11450
rect 3435 11398 3449 11450
rect 3473 11398 3487 11450
rect 3487 11398 3499 11450
rect 3499 11398 3529 11450
rect 3553 11398 3563 11450
rect 3563 11398 3609 11450
rect 3313 11396 3369 11398
rect 3393 11396 3449 11398
rect 3473 11396 3529 11398
rect 3553 11396 3609 11398
rect 4256 11450 4312 11452
rect 4336 11450 4392 11452
rect 4416 11450 4472 11452
rect 4496 11450 4552 11452
rect 4256 11398 4302 11450
rect 4302 11398 4312 11450
rect 4336 11398 4366 11450
rect 4366 11398 4378 11450
rect 4378 11398 4392 11450
rect 4416 11398 4430 11450
rect 4430 11398 4442 11450
rect 4442 11398 4472 11450
rect 4496 11398 4506 11450
rect 4506 11398 4552 11450
rect 4256 11396 4312 11398
rect 4336 11396 4392 11398
rect 4416 11396 4472 11398
rect 4496 11396 4552 11398
rect 1898 10906 1954 10908
rect 1978 10906 2034 10908
rect 2058 10906 2114 10908
rect 2138 10906 2194 10908
rect 1898 10854 1944 10906
rect 1944 10854 1954 10906
rect 1978 10854 2008 10906
rect 2008 10854 2020 10906
rect 2020 10854 2034 10906
rect 2058 10854 2072 10906
rect 2072 10854 2084 10906
rect 2084 10854 2114 10906
rect 2138 10854 2148 10906
rect 2148 10854 2194 10906
rect 1898 10852 1954 10854
rect 1978 10852 2034 10854
rect 2058 10852 2114 10854
rect 2138 10852 2194 10854
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 3081 10906 3137 10908
rect 2841 10854 2887 10906
rect 2887 10854 2897 10906
rect 2921 10854 2951 10906
rect 2951 10854 2963 10906
rect 2963 10854 2977 10906
rect 3001 10854 3015 10906
rect 3015 10854 3027 10906
rect 3027 10854 3057 10906
rect 3081 10854 3091 10906
rect 3091 10854 3137 10906
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 3081 10852 3137 10854
rect 3784 10906 3840 10908
rect 3864 10906 3920 10908
rect 3944 10906 4000 10908
rect 4024 10906 4080 10908
rect 3784 10854 3830 10906
rect 3830 10854 3840 10906
rect 3864 10854 3894 10906
rect 3894 10854 3906 10906
rect 3906 10854 3920 10906
rect 3944 10854 3958 10906
rect 3958 10854 3970 10906
rect 3970 10854 4000 10906
rect 4024 10854 4034 10906
rect 4034 10854 4080 10906
rect 3784 10852 3840 10854
rect 3864 10852 3920 10854
rect 3944 10852 4000 10854
rect 4024 10852 4080 10854
rect 4727 10906 4783 10908
rect 4807 10906 4863 10908
rect 4887 10906 4943 10908
rect 4967 10906 5023 10908
rect 4727 10854 4773 10906
rect 4773 10854 4783 10906
rect 4807 10854 4837 10906
rect 4837 10854 4849 10906
rect 4849 10854 4863 10906
rect 4887 10854 4901 10906
rect 4901 10854 4913 10906
rect 4913 10854 4943 10906
rect 4967 10854 4977 10906
rect 4977 10854 5023 10906
rect 4727 10852 4783 10854
rect 4807 10852 4863 10854
rect 4887 10852 4943 10854
rect 4967 10852 5023 10854
rect 1427 10362 1483 10364
rect 1507 10362 1563 10364
rect 1587 10362 1643 10364
rect 1667 10362 1723 10364
rect 1427 10310 1473 10362
rect 1473 10310 1483 10362
rect 1507 10310 1537 10362
rect 1537 10310 1549 10362
rect 1549 10310 1563 10362
rect 1587 10310 1601 10362
rect 1601 10310 1613 10362
rect 1613 10310 1643 10362
rect 1667 10310 1677 10362
rect 1677 10310 1723 10362
rect 1427 10308 1483 10310
rect 1507 10308 1563 10310
rect 1587 10308 1643 10310
rect 1667 10308 1723 10310
rect 2370 10362 2426 10364
rect 2450 10362 2506 10364
rect 2530 10362 2586 10364
rect 2610 10362 2666 10364
rect 2370 10310 2416 10362
rect 2416 10310 2426 10362
rect 2450 10310 2480 10362
rect 2480 10310 2492 10362
rect 2492 10310 2506 10362
rect 2530 10310 2544 10362
rect 2544 10310 2556 10362
rect 2556 10310 2586 10362
rect 2610 10310 2620 10362
rect 2620 10310 2666 10362
rect 2370 10308 2426 10310
rect 2450 10308 2506 10310
rect 2530 10308 2586 10310
rect 2610 10308 2666 10310
rect 3313 10362 3369 10364
rect 3393 10362 3449 10364
rect 3473 10362 3529 10364
rect 3553 10362 3609 10364
rect 3313 10310 3359 10362
rect 3359 10310 3369 10362
rect 3393 10310 3423 10362
rect 3423 10310 3435 10362
rect 3435 10310 3449 10362
rect 3473 10310 3487 10362
rect 3487 10310 3499 10362
rect 3499 10310 3529 10362
rect 3553 10310 3563 10362
rect 3563 10310 3609 10362
rect 3313 10308 3369 10310
rect 3393 10308 3449 10310
rect 3473 10308 3529 10310
rect 3553 10308 3609 10310
rect 4256 10362 4312 10364
rect 4336 10362 4392 10364
rect 4416 10362 4472 10364
rect 4496 10362 4552 10364
rect 4256 10310 4302 10362
rect 4302 10310 4312 10362
rect 4336 10310 4366 10362
rect 4366 10310 4378 10362
rect 4378 10310 4392 10362
rect 4416 10310 4430 10362
rect 4430 10310 4442 10362
rect 4442 10310 4472 10362
rect 4496 10310 4506 10362
rect 4506 10310 4552 10362
rect 4256 10308 4312 10310
rect 4336 10308 4392 10310
rect 4416 10308 4472 10310
rect 4496 10308 4552 10310
rect 4526 10124 4582 10160
rect 4526 10104 4528 10124
rect 4528 10104 4580 10124
rect 4580 10104 4582 10124
rect 1898 9818 1954 9820
rect 1978 9818 2034 9820
rect 2058 9818 2114 9820
rect 2138 9818 2194 9820
rect 1898 9766 1944 9818
rect 1944 9766 1954 9818
rect 1978 9766 2008 9818
rect 2008 9766 2020 9818
rect 2020 9766 2034 9818
rect 2058 9766 2072 9818
rect 2072 9766 2084 9818
rect 2084 9766 2114 9818
rect 2138 9766 2148 9818
rect 2148 9766 2194 9818
rect 1898 9764 1954 9766
rect 1978 9764 2034 9766
rect 2058 9764 2114 9766
rect 2138 9764 2194 9766
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 3081 9818 3137 9820
rect 2841 9766 2887 9818
rect 2887 9766 2897 9818
rect 2921 9766 2951 9818
rect 2951 9766 2963 9818
rect 2963 9766 2977 9818
rect 3001 9766 3015 9818
rect 3015 9766 3027 9818
rect 3027 9766 3057 9818
rect 3081 9766 3091 9818
rect 3091 9766 3137 9818
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 3081 9764 3137 9766
rect 3784 9818 3840 9820
rect 3864 9818 3920 9820
rect 3944 9818 4000 9820
rect 4024 9818 4080 9820
rect 3784 9766 3830 9818
rect 3830 9766 3840 9818
rect 3864 9766 3894 9818
rect 3894 9766 3906 9818
rect 3906 9766 3920 9818
rect 3944 9766 3958 9818
rect 3958 9766 3970 9818
rect 3970 9766 4000 9818
rect 4024 9766 4034 9818
rect 4034 9766 4080 9818
rect 3784 9764 3840 9766
rect 3864 9764 3920 9766
rect 3944 9764 4000 9766
rect 4024 9764 4080 9766
rect 4727 9818 4783 9820
rect 4807 9818 4863 9820
rect 4887 9818 4943 9820
rect 4967 9818 5023 9820
rect 4727 9766 4773 9818
rect 4773 9766 4783 9818
rect 4807 9766 4837 9818
rect 4837 9766 4849 9818
rect 4849 9766 4863 9818
rect 4887 9766 4901 9818
rect 4901 9766 4913 9818
rect 4913 9766 4943 9818
rect 4967 9766 4977 9818
rect 4977 9766 5023 9818
rect 4727 9764 4783 9766
rect 4807 9764 4863 9766
rect 4887 9764 4943 9766
rect 4967 9764 5023 9766
rect 1427 9274 1483 9276
rect 1507 9274 1563 9276
rect 1587 9274 1643 9276
rect 1667 9274 1723 9276
rect 1427 9222 1473 9274
rect 1473 9222 1483 9274
rect 1507 9222 1537 9274
rect 1537 9222 1549 9274
rect 1549 9222 1563 9274
rect 1587 9222 1601 9274
rect 1601 9222 1613 9274
rect 1613 9222 1643 9274
rect 1667 9222 1677 9274
rect 1677 9222 1723 9274
rect 1427 9220 1483 9222
rect 1507 9220 1563 9222
rect 1587 9220 1643 9222
rect 1667 9220 1723 9222
rect 2370 9274 2426 9276
rect 2450 9274 2506 9276
rect 2530 9274 2586 9276
rect 2610 9274 2666 9276
rect 2370 9222 2416 9274
rect 2416 9222 2426 9274
rect 2450 9222 2480 9274
rect 2480 9222 2492 9274
rect 2492 9222 2506 9274
rect 2530 9222 2544 9274
rect 2544 9222 2556 9274
rect 2556 9222 2586 9274
rect 2610 9222 2620 9274
rect 2620 9222 2666 9274
rect 2370 9220 2426 9222
rect 2450 9220 2506 9222
rect 2530 9220 2586 9222
rect 2610 9220 2666 9222
rect 3313 9274 3369 9276
rect 3393 9274 3449 9276
rect 3473 9274 3529 9276
rect 3553 9274 3609 9276
rect 3313 9222 3359 9274
rect 3359 9222 3369 9274
rect 3393 9222 3423 9274
rect 3423 9222 3435 9274
rect 3435 9222 3449 9274
rect 3473 9222 3487 9274
rect 3487 9222 3499 9274
rect 3499 9222 3529 9274
rect 3553 9222 3563 9274
rect 3563 9222 3609 9274
rect 3313 9220 3369 9222
rect 3393 9220 3449 9222
rect 3473 9220 3529 9222
rect 3553 9220 3609 9222
rect 4256 9274 4312 9276
rect 4336 9274 4392 9276
rect 4416 9274 4472 9276
rect 4496 9274 4552 9276
rect 4256 9222 4302 9274
rect 4302 9222 4312 9274
rect 4336 9222 4366 9274
rect 4366 9222 4378 9274
rect 4378 9222 4392 9274
rect 4416 9222 4430 9274
rect 4430 9222 4442 9274
rect 4442 9222 4472 9274
rect 4496 9222 4506 9274
rect 4506 9222 4552 9274
rect 4256 9220 4312 9222
rect 4336 9220 4392 9222
rect 4416 9220 4472 9222
rect 4496 9220 4552 9222
rect 1898 8730 1954 8732
rect 1978 8730 2034 8732
rect 2058 8730 2114 8732
rect 2138 8730 2194 8732
rect 1898 8678 1944 8730
rect 1944 8678 1954 8730
rect 1978 8678 2008 8730
rect 2008 8678 2020 8730
rect 2020 8678 2034 8730
rect 2058 8678 2072 8730
rect 2072 8678 2084 8730
rect 2084 8678 2114 8730
rect 2138 8678 2148 8730
rect 2148 8678 2194 8730
rect 1898 8676 1954 8678
rect 1978 8676 2034 8678
rect 2058 8676 2114 8678
rect 2138 8676 2194 8678
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 3081 8730 3137 8732
rect 2841 8678 2887 8730
rect 2887 8678 2897 8730
rect 2921 8678 2951 8730
rect 2951 8678 2963 8730
rect 2963 8678 2977 8730
rect 3001 8678 3015 8730
rect 3015 8678 3027 8730
rect 3027 8678 3057 8730
rect 3081 8678 3091 8730
rect 3091 8678 3137 8730
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 3081 8676 3137 8678
rect 3784 8730 3840 8732
rect 3864 8730 3920 8732
rect 3944 8730 4000 8732
rect 4024 8730 4080 8732
rect 3784 8678 3830 8730
rect 3830 8678 3840 8730
rect 3864 8678 3894 8730
rect 3894 8678 3906 8730
rect 3906 8678 3920 8730
rect 3944 8678 3958 8730
rect 3958 8678 3970 8730
rect 3970 8678 4000 8730
rect 4024 8678 4034 8730
rect 4034 8678 4080 8730
rect 3784 8676 3840 8678
rect 3864 8676 3920 8678
rect 3944 8676 4000 8678
rect 4024 8676 4080 8678
rect 4727 8730 4783 8732
rect 4807 8730 4863 8732
rect 4887 8730 4943 8732
rect 4967 8730 5023 8732
rect 4727 8678 4773 8730
rect 4773 8678 4783 8730
rect 4807 8678 4837 8730
rect 4837 8678 4849 8730
rect 4849 8678 4863 8730
rect 4887 8678 4901 8730
rect 4901 8678 4913 8730
rect 4913 8678 4943 8730
rect 4967 8678 4977 8730
rect 4977 8678 5023 8730
rect 4727 8676 4783 8678
rect 4807 8676 4863 8678
rect 4887 8676 4943 8678
rect 4967 8676 5023 8678
rect 1427 8186 1483 8188
rect 1507 8186 1563 8188
rect 1587 8186 1643 8188
rect 1667 8186 1723 8188
rect 1427 8134 1473 8186
rect 1473 8134 1483 8186
rect 1507 8134 1537 8186
rect 1537 8134 1549 8186
rect 1549 8134 1563 8186
rect 1587 8134 1601 8186
rect 1601 8134 1613 8186
rect 1613 8134 1643 8186
rect 1667 8134 1677 8186
rect 1677 8134 1723 8186
rect 1427 8132 1483 8134
rect 1507 8132 1563 8134
rect 1587 8132 1643 8134
rect 1667 8132 1723 8134
rect 2370 8186 2426 8188
rect 2450 8186 2506 8188
rect 2530 8186 2586 8188
rect 2610 8186 2666 8188
rect 2370 8134 2416 8186
rect 2416 8134 2426 8186
rect 2450 8134 2480 8186
rect 2480 8134 2492 8186
rect 2492 8134 2506 8186
rect 2530 8134 2544 8186
rect 2544 8134 2556 8186
rect 2556 8134 2586 8186
rect 2610 8134 2620 8186
rect 2620 8134 2666 8186
rect 2370 8132 2426 8134
rect 2450 8132 2506 8134
rect 2530 8132 2586 8134
rect 2610 8132 2666 8134
rect 3313 8186 3369 8188
rect 3393 8186 3449 8188
rect 3473 8186 3529 8188
rect 3553 8186 3609 8188
rect 3313 8134 3359 8186
rect 3359 8134 3369 8186
rect 3393 8134 3423 8186
rect 3423 8134 3435 8186
rect 3435 8134 3449 8186
rect 3473 8134 3487 8186
rect 3487 8134 3499 8186
rect 3499 8134 3529 8186
rect 3553 8134 3563 8186
rect 3563 8134 3609 8186
rect 3313 8132 3369 8134
rect 3393 8132 3449 8134
rect 3473 8132 3529 8134
rect 3553 8132 3609 8134
rect 4256 8186 4312 8188
rect 4336 8186 4392 8188
rect 4416 8186 4472 8188
rect 4496 8186 4552 8188
rect 4256 8134 4302 8186
rect 4302 8134 4312 8186
rect 4336 8134 4366 8186
rect 4366 8134 4378 8186
rect 4378 8134 4392 8186
rect 4416 8134 4430 8186
rect 4430 8134 4442 8186
rect 4442 8134 4472 8186
rect 4496 8134 4506 8186
rect 4506 8134 4552 8186
rect 4256 8132 4312 8134
rect 4336 8132 4392 8134
rect 4416 8132 4472 8134
rect 4496 8132 4552 8134
rect 1766 7928 1822 7984
rect 1427 7098 1483 7100
rect 1507 7098 1563 7100
rect 1587 7098 1643 7100
rect 1667 7098 1723 7100
rect 1427 7046 1473 7098
rect 1473 7046 1483 7098
rect 1507 7046 1537 7098
rect 1537 7046 1549 7098
rect 1549 7046 1563 7098
rect 1587 7046 1601 7098
rect 1601 7046 1613 7098
rect 1613 7046 1643 7098
rect 1667 7046 1677 7098
rect 1677 7046 1723 7098
rect 1427 7044 1483 7046
rect 1507 7044 1563 7046
rect 1587 7044 1643 7046
rect 1667 7044 1723 7046
rect 1898 7642 1954 7644
rect 1978 7642 2034 7644
rect 2058 7642 2114 7644
rect 2138 7642 2194 7644
rect 1898 7590 1944 7642
rect 1944 7590 1954 7642
rect 1978 7590 2008 7642
rect 2008 7590 2020 7642
rect 2020 7590 2034 7642
rect 2058 7590 2072 7642
rect 2072 7590 2084 7642
rect 2084 7590 2114 7642
rect 2138 7590 2148 7642
rect 2148 7590 2194 7642
rect 1898 7588 1954 7590
rect 1978 7588 2034 7590
rect 2058 7588 2114 7590
rect 2138 7588 2194 7590
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 3081 7642 3137 7644
rect 2841 7590 2887 7642
rect 2887 7590 2897 7642
rect 2921 7590 2951 7642
rect 2951 7590 2963 7642
rect 2963 7590 2977 7642
rect 3001 7590 3015 7642
rect 3015 7590 3027 7642
rect 3027 7590 3057 7642
rect 3081 7590 3091 7642
rect 3091 7590 3137 7642
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 3081 7588 3137 7590
rect 3784 7642 3840 7644
rect 3864 7642 3920 7644
rect 3944 7642 4000 7644
rect 4024 7642 4080 7644
rect 3784 7590 3830 7642
rect 3830 7590 3840 7642
rect 3864 7590 3894 7642
rect 3894 7590 3906 7642
rect 3906 7590 3920 7642
rect 3944 7590 3958 7642
rect 3958 7590 3970 7642
rect 3970 7590 4000 7642
rect 4024 7590 4034 7642
rect 4034 7590 4080 7642
rect 3784 7588 3840 7590
rect 3864 7588 3920 7590
rect 3944 7588 4000 7590
rect 4024 7588 4080 7590
rect 4727 7642 4783 7644
rect 4807 7642 4863 7644
rect 4887 7642 4943 7644
rect 4967 7642 5023 7644
rect 4727 7590 4773 7642
rect 4773 7590 4783 7642
rect 4807 7590 4837 7642
rect 4837 7590 4849 7642
rect 4849 7590 4863 7642
rect 4887 7590 4901 7642
rect 4901 7590 4913 7642
rect 4913 7590 4943 7642
rect 4967 7590 4977 7642
rect 4977 7590 5023 7642
rect 4727 7588 4783 7590
rect 4807 7588 4863 7590
rect 4887 7588 4943 7590
rect 4967 7588 5023 7590
rect 2370 7098 2426 7100
rect 2450 7098 2506 7100
rect 2530 7098 2586 7100
rect 2610 7098 2666 7100
rect 2370 7046 2416 7098
rect 2416 7046 2426 7098
rect 2450 7046 2480 7098
rect 2480 7046 2492 7098
rect 2492 7046 2506 7098
rect 2530 7046 2544 7098
rect 2544 7046 2556 7098
rect 2556 7046 2586 7098
rect 2610 7046 2620 7098
rect 2620 7046 2666 7098
rect 2370 7044 2426 7046
rect 2450 7044 2506 7046
rect 2530 7044 2586 7046
rect 2610 7044 2666 7046
rect 3313 7098 3369 7100
rect 3393 7098 3449 7100
rect 3473 7098 3529 7100
rect 3553 7098 3609 7100
rect 3313 7046 3359 7098
rect 3359 7046 3369 7098
rect 3393 7046 3423 7098
rect 3423 7046 3435 7098
rect 3435 7046 3449 7098
rect 3473 7046 3487 7098
rect 3487 7046 3499 7098
rect 3499 7046 3529 7098
rect 3553 7046 3563 7098
rect 3563 7046 3609 7098
rect 3313 7044 3369 7046
rect 3393 7044 3449 7046
rect 3473 7044 3529 7046
rect 3553 7044 3609 7046
rect 4256 7098 4312 7100
rect 4336 7098 4392 7100
rect 4416 7098 4472 7100
rect 4496 7098 4552 7100
rect 4256 7046 4302 7098
rect 4302 7046 4312 7098
rect 4336 7046 4366 7098
rect 4366 7046 4378 7098
rect 4378 7046 4392 7098
rect 4416 7046 4430 7098
rect 4430 7046 4442 7098
rect 4442 7046 4472 7098
rect 4496 7046 4506 7098
rect 4506 7046 4552 7098
rect 4256 7044 4312 7046
rect 4336 7044 4392 7046
rect 4416 7044 4472 7046
rect 4496 7044 4552 7046
rect 1898 6554 1954 6556
rect 1978 6554 2034 6556
rect 2058 6554 2114 6556
rect 2138 6554 2194 6556
rect 1898 6502 1944 6554
rect 1944 6502 1954 6554
rect 1978 6502 2008 6554
rect 2008 6502 2020 6554
rect 2020 6502 2034 6554
rect 2058 6502 2072 6554
rect 2072 6502 2084 6554
rect 2084 6502 2114 6554
rect 2138 6502 2148 6554
rect 2148 6502 2194 6554
rect 1898 6500 1954 6502
rect 1978 6500 2034 6502
rect 2058 6500 2114 6502
rect 2138 6500 2194 6502
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 3081 6554 3137 6556
rect 2841 6502 2887 6554
rect 2887 6502 2897 6554
rect 2921 6502 2951 6554
rect 2951 6502 2963 6554
rect 2963 6502 2977 6554
rect 3001 6502 3015 6554
rect 3015 6502 3027 6554
rect 3027 6502 3057 6554
rect 3081 6502 3091 6554
rect 3091 6502 3137 6554
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 3081 6500 3137 6502
rect 3784 6554 3840 6556
rect 3864 6554 3920 6556
rect 3944 6554 4000 6556
rect 4024 6554 4080 6556
rect 3784 6502 3830 6554
rect 3830 6502 3840 6554
rect 3864 6502 3894 6554
rect 3894 6502 3906 6554
rect 3906 6502 3920 6554
rect 3944 6502 3958 6554
rect 3958 6502 3970 6554
rect 3970 6502 4000 6554
rect 4024 6502 4034 6554
rect 4034 6502 4080 6554
rect 3784 6500 3840 6502
rect 3864 6500 3920 6502
rect 3944 6500 4000 6502
rect 4024 6500 4080 6502
rect 4727 6554 4783 6556
rect 4807 6554 4863 6556
rect 4887 6554 4943 6556
rect 4967 6554 5023 6556
rect 4727 6502 4773 6554
rect 4773 6502 4783 6554
rect 4807 6502 4837 6554
rect 4837 6502 4849 6554
rect 4849 6502 4863 6554
rect 4887 6502 4901 6554
rect 4901 6502 4913 6554
rect 4913 6502 4943 6554
rect 4967 6502 4977 6554
rect 4977 6502 5023 6554
rect 4727 6500 4783 6502
rect 4807 6500 4863 6502
rect 4887 6500 4943 6502
rect 4967 6500 5023 6502
rect 1427 6010 1483 6012
rect 1507 6010 1563 6012
rect 1587 6010 1643 6012
rect 1667 6010 1723 6012
rect 1427 5958 1473 6010
rect 1473 5958 1483 6010
rect 1507 5958 1537 6010
rect 1537 5958 1549 6010
rect 1549 5958 1563 6010
rect 1587 5958 1601 6010
rect 1601 5958 1613 6010
rect 1613 5958 1643 6010
rect 1667 5958 1677 6010
rect 1677 5958 1723 6010
rect 1427 5956 1483 5958
rect 1507 5956 1563 5958
rect 1587 5956 1643 5958
rect 1667 5956 1723 5958
rect 2370 6010 2426 6012
rect 2450 6010 2506 6012
rect 2530 6010 2586 6012
rect 2610 6010 2666 6012
rect 2370 5958 2416 6010
rect 2416 5958 2426 6010
rect 2450 5958 2480 6010
rect 2480 5958 2492 6010
rect 2492 5958 2506 6010
rect 2530 5958 2544 6010
rect 2544 5958 2556 6010
rect 2556 5958 2586 6010
rect 2610 5958 2620 6010
rect 2620 5958 2666 6010
rect 2370 5956 2426 5958
rect 2450 5956 2506 5958
rect 2530 5956 2586 5958
rect 2610 5956 2666 5958
rect 3313 6010 3369 6012
rect 3393 6010 3449 6012
rect 3473 6010 3529 6012
rect 3553 6010 3609 6012
rect 3313 5958 3359 6010
rect 3359 5958 3369 6010
rect 3393 5958 3423 6010
rect 3423 5958 3435 6010
rect 3435 5958 3449 6010
rect 3473 5958 3487 6010
rect 3487 5958 3499 6010
rect 3499 5958 3529 6010
rect 3553 5958 3563 6010
rect 3563 5958 3609 6010
rect 3313 5956 3369 5958
rect 3393 5956 3449 5958
rect 3473 5956 3529 5958
rect 3553 5956 3609 5958
rect 1898 5466 1954 5468
rect 1978 5466 2034 5468
rect 2058 5466 2114 5468
rect 2138 5466 2194 5468
rect 1898 5414 1944 5466
rect 1944 5414 1954 5466
rect 1978 5414 2008 5466
rect 2008 5414 2020 5466
rect 2020 5414 2034 5466
rect 2058 5414 2072 5466
rect 2072 5414 2084 5466
rect 2084 5414 2114 5466
rect 2138 5414 2148 5466
rect 2148 5414 2194 5466
rect 1898 5412 1954 5414
rect 1978 5412 2034 5414
rect 2058 5412 2114 5414
rect 2138 5412 2194 5414
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 3081 5466 3137 5468
rect 2841 5414 2887 5466
rect 2887 5414 2897 5466
rect 2921 5414 2951 5466
rect 2951 5414 2963 5466
rect 2963 5414 2977 5466
rect 3001 5414 3015 5466
rect 3015 5414 3027 5466
rect 3027 5414 3057 5466
rect 3081 5414 3091 5466
rect 3091 5414 3137 5466
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 3081 5412 3137 5414
rect 3784 5466 3840 5468
rect 3864 5466 3920 5468
rect 3944 5466 4000 5468
rect 4024 5466 4080 5468
rect 3784 5414 3830 5466
rect 3830 5414 3840 5466
rect 3864 5414 3894 5466
rect 3894 5414 3906 5466
rect 3906 5414 3920 5466
rect 3944 5414 3958 5466
rect 3958 5414 3970 5466
rect 3970 5414 4000 5466
rect 4024 5414 4034 5466
rect 4034 5414 4080 5466
rect 3784 5412 3840 5414
rect 3864 5412 3920 5414
rect 3944 5412 4000 5414
rect 4024 5412 4080 5414
rect 1427 4922 1483 4924
rect 1507 4922 1563 4924
rect 1587 4922 1643 4924
rect 1667 4922 1723 4924
rect 1427 4870 1473 4922
rect 1473 4870 1483 4922
rect 1507 4870 1537 4922
rect 1537 4870 1549 4922
rect 1549 4870 1563 4922
rect 1587 4870 1601 4922
rect 1601 4870 1613 4922
rect 1613 4870 1643 4922
rect 1667 4870 1677 4922
rect 1677 4870 1723 4922
rect 1427 4868 1483 4870
rect 1507 4868 1563 4870
rect 1587 4868 1643 4870
rect 1667 4868 1723 4870
rect 2370 4922 2426 4924
rect 2450 4922 2506 4924
rect 2530 4922 2586 4924
rect 2610 4922 2666 4924
rect 2370 4870 2416 4922
rect 2416 4870 2426 4922
rect 2450 4870 2480 4922
rect 2480 4870 2492 4922
rect 2492 4870 2506 4922
rect 2530 4870 2544 4922
rect 2544 4870 2556 4922
rect 2556 4870 2586 4922
rect 2610 4870 2620 4922
rect 2620 4870 2666 4922
rect 2370 4868 2426 4870
rect 2450 4868 2506 4870
rect 2530 4868 2586 4870
rect 2610 4868 2666 4870
rect 3313 4922 3369 4924
rect 3393 4922 3449 4924
rect 3473 4922 3529 4924
rect 3553 4922 3609 4924
rect 3313 4870 3359 4922
rect 3359 4870 3369 4922
rect 3393 4870 3423 4922
rect 3423 4870 3435 4922
rect 3435 4870 3449 4922
rect 3473 4870 3487 4922
rect 3487 4870 3499 4922
rect 3499 4870 3529 4922
rect 3553 4870 3563 4922
rect 3563 4870 3609 4922
rect 3313 4868 3369 4870
rect 3393 4868 3449 4870
rect 3473 4868 3529 4870
rect 3553 4868 3609 4870
rect 1898 4378 1954 4380
rect 1978 4378 2034 4380
rect 2058 4378 2114 4380
rect 2138 4378 2194 4380
rect 1898 4326 1944 4378
rect 1944 4326 1954 4378
rect 1978 4326 2008 4378
rect 2008 4326 2020 4378
rect 2020 4326 2034 4378
rect 2058 4326 2072 4378
rect 2072 4326 2084 4378
rect 2084 4326 2114 4378
rect 2138 4326 2148 4378
rect 2148 4326 2194 4378
rect 1898 4324 1954 4326
rect 1978 4324 2034 4326
rect 2058 4324 2114 4326
rect 2138 4324 2194 4326
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 3081 4378 3137 4380
rect 2841 4326 2887 4378
rect 2887 4326 2897 4378
rect 2921 4326 2951 4378
rect 2951 4326 2963 4378
rect 2963 4326 2977 4378
rect 3001 4326 3015 4378
rect 3015 4326 3027 4378
rect 3027 4326 3057 4378
rect 3081 4326 3091 4378
rect 3091 4326 3137 4378
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 3081 4324 3137 4326
rect 3784 4378 3840 4380
rect 3864 4378 3920 4380
rect 3944 4378 4000 4380
rect 4024 4378 4080 4380
rect 3784 4326 3830 4378
rect 3830 4326 3840 4378
rect 3864 4326 3894 4378
rect 3894 4326 3906 4378
rect 3906 4326 3920 4378
rect 3944 4326 3958 4378
rect 3958 4326 3970 4378
rect 3970 4326 4000 4378
rect 4024 4326 4034 4378
rect 4034 4326 4080 4378
rect 3784 4324 3840 4326
rect 3864 4324 3920 4326
rect 3944 4324 4000 4326
rect 4024 4324 4080 4326
rect 1427 3834 1483 3836
rect 1507 3834 1563 3836
rect 1587 3834 1643 3836
rect 1667 3834 1723 3836
rect 1427 3782 1473 3834
rect 1473 3782 1483 3834
rect 1507 3782 1537 3834
rect 1537 3782 1549 3834
rect 1549 3782 1563 3834
rect 1587 3782 1601 3834
rect 1601 3782 1613 3834
rect 1613 3782 1643 3834
rect 1667 3782 1677 3834
rect 1677 3782 1723 3834
rect 1427 3780 1483 3782
rect 1507 3780 1563 3782
rect 1587 3780 1643 3782
rect 1667 3780 1723 3782
rect 2370 3834 2426 3836
rect 2450 3834 2506 3836
rect 2530 3834 2586 3836
rect 2610 3834 2666 3836
rect 2370 3782 2416 3834
rect 2416 3782 2426 3834
rect 2450 3782 2480 3834
rect 2480 3782 2492 3834
rect 2492 3782 2506 3834
rect 2530 3782 2544 3834
rect 2544 3782 2556 3834
rect 2556 3782 2586 3834
rect 2610 3782 2620 3834
rect 2620 3782 2666 3834
rect 2370 3780 2426 3782
rect 2450 3780 2506 3782
rect 2530 3780 2586 3782
rect 2610 3780 2666 3782
rect 3313 3834 3369 3836
rect 3393 3834 3449 3836
rect 3473 3834 3529 3836
rect 3553 3834 3609 3836
rect 3313 3782 3359 3834
rect 3359 3782 3369 3834
rect 3393 3782 3423 3834
rect 3423 3782 3435 3834
rect 3435 3782 3449 3834
rect 3473 3782 3487 3834
rect 3487 3782 3499 3834
rect 3499 3782 3529 3834
rect 3553 3782 3563 3834
rect 3563 3782 3609 3834
rect 3313 3780 3369 3782
rect 3393 3780 3449 3782
rect 3473 3780 3529 3782
rect 3553 3780 3609 3782
rect 1898 3290 1954 3292
rect 1978 3290 2034 3292
rect 2058 3290 2114 3292
rect 2138 3290 2194 3292
rect 1898 3238 1944 3290
rect 1944 3238 1954 3290
rect 1978 3238 2008 3290
rect 2008 3238 2020 3290
rect 2020 3238 2034 3290
rect 2058 3238 2072 3290
rect 2072 3238 2084 3290
rect 2084 3238 2114 3290
rect 2138 3238 2148 3290
rect 2148 3238 2194 3290
rect 1898 3236 1954 3238
rect 1978 3236 2034 3238
rect 2058 3236 2114 3238
rect 2138 3236 2194 3238
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 3081 3290 3137 3292
rect 2841 3238 2887 3290
rect 2887 3238 2897 3290
rect 2921 3238 2951 3290
rect 2951 3238 2963 3290
rect 2963 3238 2977 3290
rect 3001 3238 3015 3290
rect 3015 3238 3027 3290
rect 3027 3238 3057 3290
rect 3081 3238 3091 3290
rect 3091 3238 3137 3290
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 3081 3236 3137 3238
rect 3784 3290 3840 3292
rect 3864 3290 3920 3292
rect 3944 3290 4000 3292
rect 4024 3290 4080 3292
rect 3784 3238 3830 3290
rect 3830 3238 3840 3290
rect 3864 3238 3894 3290
rect 3894 3238 3906 3290
rect 3906 3238 3920 3290
rect 3944 3238 3958 3290
rect 3958 3238 3970 3290
rect 3970 3238 4000 3290
rect 4024 3238 4034 3290
rect 4034 3238 4080 3290
rect 3784 3236 3840 3238
rect 3864 3236 3920 3238
rect 3944 3236 4000 3238
rect 4024 3236 4080 3238
rect 1427 2746 1483 2748
rect 1507 2746 1563 2748
rect 1587 2746 1643 2748
rect 1667 2746 1723 2748
rect 1427 2694 1473 2746
rect 1473 2694 1483 2746
rect 1507 2694 1537 2746
rect 1537 2694 1549 2746
rect 1549 2694 1563 2746
rect 1587 2694 1601 2746
rect 1601 2694 1613 2746
rect 1613 2694 1643 2746
rect 1667 2694 1677 2746
rect 1677 2694 1723 2746
rect 1427 2692 1483 2694
rect 1507 2692 1563 2694
rect 1587 2692 1643 2694
rect 1667 2692 1723 2694
rect 2370 2746 2426 2748
rect 2450 2746 2506 2748
rect 2530 2746 2586 2748
rect 2610 2746 2666 2748
rect 2370 2694 2416 2746
rect 2416 2694 2426 2746
rect 2450 2694 2480 2746
rect 2480 2694 2492 2746
rect 2492 2694 2506 2746
rect 2530 2694 2544 2746
rect 2544 2694 2556 2746
rect 2556 2694 2586 2746
rect 2610 2694 2620 2746
rect 2620 2694 2666 2746
rect 2370 2692 2426 2694
rect 2450 2692 2506 2694
rect 2530 2692 2586 2694
rect 2610 2692 2666 2694
rect 3313 2746 3369 2748
rect 3393 2746 3449 2748
rect 3473 2746 3529 2748
rect 3553 2746 3609 2748
rect 3313 2694 3359 2746
rect 3359 2694 3369 2746
rect 3393 2694 3423 2746
rect 3423 2694 3435 2746
rect 3435 2694 3449 2746
rect 3473 2694 3487 2746
rect 3487 2694 3499 2746
rect 3499 2694 3529 2746
rect 3553 2694 3563 2746
rect 3563 2694 3609 2746
rect 3313 2692 3369 2694
rect 3393 2692 3449 2694
rect 3473 2692 3529 2694
rect 3553 2692 3609 2694
rect 4256 6010 4312 6012
rect 4336 6010 4392 6012
rect 4416 6010 4472 6012
rect 4496 6010 4552 6012
rect 4256 5958 4302 6010
rect 4302 5958 4312 6010
rect 4336 5958 4366 6010
rect 4366 5958 4378 6010
rect 4378 5958 4392 6010
rect 4416 5958 4430 6010
rect 4430 5958 4442 6010
rect 4442 5958 4472 6010
rect 4496 5958 4506 6010
rect 4506 5958 4552 6010
rect 4256 5956 4312 5958
rect 4336 5956 4392 5958
rect 4416 5956 4472 5958
rect 4496 5956 4552 5958
rect 4802 6024 4858 6080
rect 4727 5466 4783 5468
rect 4807 5466 4863 5468
rect 4887 5466 4943 5468
rect 4967 5466 5023 5468
rect 4727 5414 4773 5466
rect 4773 5414 4783 5466
rect 4807 5414 4837 5466
rect 4837 5414 4849 5466
rect 4849 5414 4863 5466
rect 4887 5414 4901 5466
rect 4901 5414 4913 5466
rect 4913 5414 4943 5466
rect 4967 5414 4977 5466
rect 4977 5414 5023 5466
rect 4727 5412 4783 5414
rect 4807 5412 4863 5414
rect 4887 5412 4943 5414
rect 4967 5412 5023 5414
rect 4256 4922 4312 4924
rect 4336 4922 4392 4924
rect 4416 4922 4472 4924
rect 4496 4922 4552 4924
rect 4256 4870 4302 4922
rect 4302 4870 4312 4922
rect 4336 4870 4366 4922
rect 4366 4870 4378 4922
rect 4378 4870 4392 4922
rect 4416 4870 4430 4922
rect 4430 4870 4442 4922
rect 4442 4870 4472 4922
rect 4496 4870 4506 4922
rect 4506 4870 4552 4922
rect 4256 4868 4312 4870
rect 4336 4868 4392 4870
rect 4416 4868 4472 4870
rect 4496 4868 4552 4870
rect 4727 4378 4783 4380
rect 4807 4378 4863 4380
rect 4887 4378 4943 4380
rect 4967 4378 5023 4380
rect 4727 4326 4773 4378
rect 4773 4326 4783 4378
rect 4807 4326 4837 4378
rect 4837 4326 4849 4378
rect 4849 4326 4863 4378
rect 4887 4326 4901 4378
rect 4901 4326 4913 4378
rect 4913 4326 4943 4378
rect 4967 4326 4977 4378
rect 4977 4326 5023 4378
rect 4727 4324 4783 4326
rect 4807 4324 4863 4326
rect 4887 4324 4943 4326
rect 4967 4324 5023 4326
rect 4256 3834 4312 3836
rect 4336 3834 4392 3836
rect 4416 3834 4472 3836
rect 4496 3834 4552 3836
rect 4256 3782 4302 3834
rect 4302 3782 4312 3834
rect 4336 3782 4366 3834
rect 4366 3782 4378 3834
rect 4378 3782 4392 3834
rect 4416 3782 4430 3834
rect 4430 3782 4442 3834
rect 4442 3782 4472 3834
rect 4496 3782 4506 3834
rect 4506 3782 4552 3834
rect 4256 3780 4312 3782
rect 4336 3780 4392 3782
rect 4416 3780 4472 3782
rect 4496 3780 4552 3782
rect 4727 3290 4783 3292
rect 4807 3290 4863 3292
rect 4887 3290 4943 3292
rect 4967 3290 5023 3292
rect 4727 3238 4773 3290
rect 4773 3238 4783 3290
rect 4807 3238 4837 3290
rect 4837 3238 4849 3290
rect 4849 3238 4863 3290
rect 4887 3238 4901 3290
rect 4901 3238 4913 3290
rect 4913 3238 4943 3290
rect 4967 3238 4977 3290
rect 4977 3238 5023 3290
rect 4727 3236 4783 3238
rect 4807 3236 4863 3238
rect 4887 3236 4943 3238
rect 4967 3236 5023 3238
rect 4256 2746 4312 2748
rect 4336 2746 4392 2748
rect 4416 2746 4472 2748
rect 4496 2746 4552 2748
rect 4256 2694 4302 2746
rect 4302 2694 4312 2746
rect 4336 2694 4366 2746
rect 4366 2694 4378 2746
rect 4378 2694 4392 2746
rect 4416 2694 4430 2746
rect 4430 2694 4442 2746
rect 4442 2694 4472 2746
rect 4496 2694 4506 2746
rect 4506 2694 4552 2746
rect 4256 2692 4312 2694
rect 4336 2692 4392 2694
rect 4416 2692 4472 2694
rect 4496 2692 4552 2694
rect 4894 2508 4950 2544
rect 4894 2488 4896 2508
rect 4896 2488 4948 2508
rect 4948 2488 4950 2508
rect 1898 2202 1954 2204
rect 1978 2202 2034 2204
rect 2058 2202 2114 2204
rect 2138 2202 2194 2204
rect 1898 2150 1944 2202
rect 1944 2150 1954 2202
rect 1978 2150 2008 2202
rect 2008 2150 2020 2202
rect 2020 2150 2034 2202
rect 2058 2150 2072 2202
rect 2072 2150 2084 2202
rect 2084 2150 2114 2202
rect 2138 2150 2148 2202
rect 2148 2150 2194 2202
rect 1898 2148 1954 2150
rect 1978 2148 2034 2150
rect 2058 2148 2114 2150
rect 2138 2148 2194 2150
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 3081 2202 3137 2204
rect 2841 2150 2887 2202
rect 2887 2150 2897 2202
rect 2921 2150 2951 2202
rect 2951 2150 2963 2202
rect 2963 2150 2977 2202
rect 3001 2150 3015 2202
rect 3015 2150 3027 2202
rect 3027 2150 3057 2202
rect 3081 2150 3091 2202
rect 3091 2150 3137 2202
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 3081 2148 3137 2150
rect 3784 2202 3840 2204
rect 3864 2202 3920 2204
rect 3944 2202 4000 2204
rect 4024 2202 4080 2204
rect 3784 2150 3830 2202
rect 3830 2150 3840 2202
rect 3864 2150 3894 2202
rect 3894 2150 3906 2202
rect 3906 2150 3920 2202
rect 3944 2150 3958 2202
rect 3958 2150 3970 2202
rect 3970 2150 4000 2202
rect 4024 2150 4034 2202
rect 4034 2150 4080 2202
rect 3784 2148 3840 2150
rect 3864 2148 3920 2150
rect 3944 2148 4000 2150
rect 4024 2148 4080 2150
rect 4727 2202 4783 2204
rect 4807 2202 4863 2204
rect 4887 2202 4943 2204
rect 4967 2202 5023 2204
rect 4727 2150 4773 2202
rect 4773 2150 4783 2202
rect 4807 2150 4837 2202
rect 4837 2150 4849 2202
rect 4849 2150 4863 2202
rect 4887 2150 4901 2202
rect 4901 2150 4913 2202
rect 4913 2150 4943 2202
rect 4967 2150 4977 2202
rect 4977 2150 5023 2202
rect 4727 2148 4783 2150
rect 4807 2148 4863 2150
rect 4887 2148 4943 2150
rect 4967 2148 5023 2150
<< metal3 >>
rect 4889 13698 4955 13701
rect 5200 13698 6000 13728
rect 4889 13696 6000 13698
rect 4889 13640 4894 13696
rect 4950 13640 6000 13696
rect 4889 13638 6000 13640
rect 4889 13635 4955 13638
rect 1417 13632 1733 13633
rect 1417 13568 1423 13632
rect 1487 13568 1503 13632
rect 1567 13568 1583 13632
rect 1647 13568 1663 13632
rect 1727 13568 1733 13632
rect 1417 13567 1733 13568
rect 2360 13632 2676 13633
rect 2360 13568 2366 13632
rect 2430 13568 2446 13632
rect 2510 13568 2526 13632
rect 2590 13568 2606 13632
rect 2670 13568 2676 13632
rect 2360 13567 2676 13568
rect 3303 13632 3619 13633
rect 3303 13568 3309 13632
rect 3373 13568 3389 13632
rect 3453 13568 3469 13632
rect 3533 13568 3549 13632
rect 3613 13568 3619 13632
rect 3303 13567 3619 13568
rect 4246 13632 4562 13633
rect 4246 13568 4252 13632
rect 4316 13568 4332 13632
rect 4396 13568 4412 13632
rect 4476 13568 4492 13632
rect 4556 13568 4562 13632
rect 5200 13608 6000 13638
rect 4246 13567 4562 13568
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 1888 13088 2204 13089
rect 1888 13024 1894 13088
rect 1958 13024 1974 13088
rect 2038 13024 2054 13088
rect 2118 13024 2134 13088
rect 2198 13024 2204 13088
rect 1888 13023 2204 13024
rect 2831 13088 3147 13089
rect 2831 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3077 13088
rect 3141 13024 3147 13088
rect 2831 13023 3147 13024
rect 3774 13088 4090 13089
rect 3774 13024 3780 13088
rect 3844 13024 3860 13088
rect 3924 13024 3940 13088
rect 4004 13024 4020 13088
rect 4084 13024 4090 13088
rect 3774 13023 4090 13024
rect 4717 13088 5033 13089
rect 4717 13024 4723 13088
rect 4787 13024 4803 13088
rect 4867 13024 4883 13088
rect 4947 13024 4963 13088
rect 5027 13024 5033 13088
rect 4717 13023 5033 13024
rect 1417 12544 1733 12545
rect 1417 12480 1423 12544
rect 1487 12480 1503 12544
rect 1567 12480 1583 12544
rect 1647 12480 1663 12544
rect 1727 12480 1733 12544
rect 1417 12479 1733 12480
rect 2360 12544 2676 12545
rect 2360 12480 2366 12544
rect 2430 12480 2446 12544
rect 2510 12480 2526 12544
rect 2590 12480 2606 12544
rect 2670 12480 2676 12544
rect 2360 12479 2676 12480
rect 3303 12544 3619 12545
rect 3303 12480 3309 12544
rect 3373 12480 3389 12544
rect 3453 12480 3469 12544
rect 3533 12480 3549 12544
rect 3613 12480 3619 12544
rect 3303 12479 3619 12480
rect 4246 12544 4562 12545
rect 4246 12480 4252 12544
rect 4316 12480 4332 12544
rect 4396 12480 4412 12544
rect 4476 12480 4492 12544
rect 4556 12480 4562 12544
rect 4246 12479 4562 12480
rect 1888 12000 2204 12001
rect 1888 11936 1894 12000
rect 1958 11936 1974 12000
rect 2038 11936 2054 12000
rect 2118 11936 2134 12000
rect 2198 11936 2204 12000
rect 1888 11935 2204 11936
rect 2831 12000 3147 12001
rect 2831 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3077 12000
rect 3141 11936 3147 12000
rect 2831 11935 3147 11936
rect 3774 12000 4090 12001
rect 3774 11936 3780 12000
rect 3844 11936 3860 12000
rect 3924 11936 3940 12000
rect 4004 11936 4020 12000
rect 4084 11936 4090 12000
rect 3774 11935 4090 11936
rect 4717 12000 5033 12001
rect 4717 11936 4723 12000
rect 4787 11936 4803 12000
rect 4867 11936 4883 12000
rect 4947 11936 4963 12000
rect 5027 11936 5033 12000
rect 4717 11935 5033 11936
rect 1417 11456 1733 11457
rect 1417 11392 1423 11456
rect 1487 11392 1503 11456
rect 1567 11392 1583 11456
rect 1647 11392 1663 11456
rect 1727 11392 1733 11456
rect 1417 11391 1733 11392
rect 2360 11456 2676 11457
rect 2360 11392 2366 11456
rect 2430 11392 2446 11456
rect 2510 11392 2526 11456
rect 2590 11392 2606 11456
rect 2670 11392 2676 11456
rect 2360 11391 2676 11392
rect 3303 11456 3619 11457
rect 3303 11392 3309 11456
rect 3373 11392 3389 11456
rect 3453 11392 3469 11456
rect 3533 11392 3549 11456
rect 3613 11392 3619 11456
rect 3303 11391 3619 11392
rect 4246 11456 4562 11457
rect 4246 11392 4252 11456
rect 4316 11392 4332 11456
rect 4396 11392 4412 11456
rect 4476 11392 4492 11456
rect 4556 11392 4562 11456
rect 4246 11391 4562 11392
rect 1888 10912 2204 10913
rect 1888 10848 1894 10912
rect 1958 10848 1974 10912
rect 2038 10848 2054 10912
rect 2118 10848 2134 10912
rect 2198 10848 2204 10912
rect 1888 10847 2204 10848
rect 2831 10912 3147 10913
rect 2831 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3077 10912
rect 3141 10848 3147 10912
rect 2831 10847 3147 10848
rect 3774 10912 4090 10913
rect 3774 10848 3780 10912
rect 3844 10848 3860 10912
rect 3924 10848 3940 10912
rect 4004 10848 4020 10912
rect 4084 10848 4090 10912
rect 3774 10847 4090 10848
rect 4717 10912 5033 10913
rect 4717 10848 4723 10912
rect 4787 10848 4803 10912
rect 4867 10848 4883 10912
rect 4947 10848 4963 10912
rect 5027 10848 5033 10912
rect 4717 10847 5033 10848
rect 1417 10368 1733 10369
rect 1417 10304 1423 10368
rect 1487 10304 1503 10368
rect 1567 10304 1583 10368
rect 1647 10304 1663 10368
rect 1727 10304 1733 10368
rect 1417 10303 1733 10304
rect 2360 10368 2676 10369
rect 2360 10304 2366 10368
rect 2430 10304 2446 10368
rect 2510 10304 2526 10368
rect 2590 10304 2606 10368
rect 2670 10304 2676 10368
rect 2360 10303 2676 10304
rect 3303 10368 3619 10369
rect 3303 10304 3309 10368
rect 3373 10304 3389 10368
rect 3453 10304 3469 10368
rect 3533 10304 3549 10368
rect 3613 10304 3619 10368
rect 3303 10303 3619 10304
rect 4246 10368 4562 10369
rect 4246 10304 4252 10368
rect 4316 10304 4332 10368
rect 4396 10304 4412 10368
rect 4476 10304 4492 10368
rect 4556 10304 4562 10368
rect 4246 10303 4562 10304
rect 4521 10162 4587 10165
rect 4521 10160 5458 10162
rect 4521 10104 4526 10160
rect 4582 10104 5458 10160
rect 4521 10102 5458 10104
rect 4521 10099 4587 10102
rect 5398 9920 5458 10102
rect 1888 9824 2204 9825
rect 1888 9760 1894 9824
rect 1958 9760 1974 9824
rect 2038 9760 2054 9824
rect 2118 9760 2134 9824
rect 2198 9760 2204 9824
rect 1888 9759 2204 9760
rect 2831 9824 3147 9825
rect 2831 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3077 9824
rect 3141 9760 3147 9824
rect 2831 9759 3147 9760
rect 3774 9824 4090 9825
rect 3774 9760 3780 9824
rect 3844 9760 3860 9824
rect 3924 9760 3940 9824
rect 4004 9760 4020 9824
rect 4084 9760 4090 9824
rect 3774 9759 4090 9760
rect 4717 9824 5033 9825
rect 4717 9760 4723 9824
rect 4787 9760 4803 9824
rect 4867 9760 4883 9824
rect 4947 9760 4963 9824
rect 5027 9760 5033 9824
rect 5200 9800 6000 9920
rect 4717 9759 5033 9760
rect 1417 9280 1733 9281
rect 1417 9216 1423 9280
rect 1487 9216 1503 9280
rect 1567 9216 1583 9280
rect 1647 9216 1663 9280
rect 1727 9216 1733 9280
rect 1417 9215 1733 9216
rect 2360 9280 2676 9281
rect 2360 9216 2366 9280
rect 2430 9216 2446 9280
rect 2510 9216 2526 9280
rect 2590 9216 2606 9280
rect 2670 9216 2676 9280
rect 2360 9215 2676 9216
rect 3303 9280 3619 9281
rect 3303 9216 3309 9280
rect 3373 9216 3389 9280
rect 3453 9216 3469 9280
rect 3533 9216 3549 9280
rect 3613 9216 3619 9280
rect 3303 9215 3619 9216
rect 4246 9280 4562 9281
rect 4246 9216 4252 9280
rect 4316 9216 4332 9280
rect 4396 9216 4412 9280
rect 4476 9216 4492 9280
rect 4556 9216 4562 9280
rect 4246 9215 4562 9216
rect 1888 8736 2204 8737
rect 1888 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2204 8736
rect 1888 8671 2204 8672
rect 2831 8736 3147 8737
rect 2831 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3147 8736
rect 2831 8671 3147 8672
rect 3774 8736 4090 8737
rect 3774 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4090 8736
rect 3774 8671 4090 8672
rect 4717 8736 5033 8737
rect 4717 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5033 8736
rect 4717 8671 5033 8672
rect 1417 8192 1733 8193
rect 1417 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1733 8192
rect 1417 8127 1733 8128
rect 2360 8192 2676 8193
rect 2360 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2676 8192
rect 2360 8127 2676 8128
rect 3303 8192 3619 8193
rect 3303 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3619 8192
rect 3303 8127 3619 8128
rect 4246 8192 4562 8193
rect 4246 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4562 8192
rect 4246 8127 4562 8128
rect 0 7986 800 8016
rect 1761 7986 1827 7989
rect 0 7984 1827 7986
rect 0 7928 1766 7984
rect 1822 7928 1827 7984
rect 0 7926 1827 7928
rect 0 7896 800 7926
rect 1761 7923 1827 7926
rect 1888 7648 2204 7649
rect 1888 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2204 7648
rect 1888 7583 2204 7584
rect 2831 7648 3147 7649
rect 2831 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3147 7648
rect 2831 7583 3147 7584
rect 3774 7648 4090 7649
rect 3774 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4090 7648
rect 3774 7583 4090 7584
rect 4717 7648 5033 7649
rect 4717 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5033 7648
rect 4717 7583 5033 7584
rect 1417 7104 1733 7105
rect 1417 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1733 7104
rect 1417 7039 1733 7040
rect 2360 7104 2676 7105
rect 2360 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2676 7104
rect 2360 7039 2676 7040
rect 3303 7104 3619 7105
rect 3303 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3619 7104
rect 3303 7039 3619 7040
rect 4246 7104 4562 7105
rect 4246 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4562 7104
rect 4246 7039 4562 7040
rect 1888 6560 2204 6561
rect 1888 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2204 6560
rect 1888 6495 2204 6496
rect 2831 6560 3147 6561
rect 2831 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3147 6560
rect 2831 6495 3147 6496
rect 3774 6560 4090 6561
rect 3774 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4090 6560
rect 3774 6495 4090 6496
rect 4717 6560 5033 6561
rect 4717 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5033 6560
rect 4717 6495 5033 6496
rect 4797 6082 4863 6085
rect 5200 6082 6000 6112
rect 4797 6080 6000 6082
rect 4797 6024 4802 6080
rect 4858 6024 6000 6080
rect 4797 6022 6000 6024
rect 4797 6019 4863 6022
rect 1417 6016 1733 6017
rect 1417 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1733 6016
rect 1417 5951 1733 5952
rect 2360 6016 2676 6017
rect 2360 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2676 6016
rect 2360 5951 2676 5952
rect 3303 6016 3619 6017
rect 3303 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3619 6016
rect 3303 5951 3619 5952
rect 4246 6016 4562 6017
rect 4246 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4562 6016
rect 5200 5992 6000 6022
rect 4246 5951 4562 5952
rect 1888 5472 2204 5473
rect 1888 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2204 5472
rect 1888 5407 2204 5408
rect 2831 5472 3147 5473
rect 2831 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3147 5472
rect 2831 5407 3147 5408
rect 3774 5472 4090 5473
rect 3774 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4090 5472
rect 3774 5407 4090 5408
rect 4717 5472 5033 5473
rect 4717 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5033 5472
rect 4717 5407 5033 5408
rect 1417 4928 1733 4929
rect 1417 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1733 4928
rect 1417 4863 1733 4864
rect 2360 4928 2676 4929
rect 2360 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2676 4928
rect 2360 4863 2676 4864
rect 3303 4928 3619 4929
rect 3303 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3619 4928
rect 3303 4863 3619 4864
rect 4246 4928 4562 4929
rect 4246 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4562 4928
rect 4246 4863 4562 4864
rect 1888 4384 2204 4385
rect 1888 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2204 4384
rect 1888 4319 2204 4320
rect 2831 4384 3147 4385
rect 2831 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3147 4384
rect 2831 4319 3147 4320
rect 3774 4384 4090 4385
rect 3774 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4090 4384
rect 3774 4319 4090 4320
rect 4717 4384 5033 4385
rect 4717 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5033 4384
rect 4717 4319 5033 4320
rect 1417 3840 1733 3841
rect 1417 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1733 3840
rect 1417 3775 1733 3776
rect 2360 3840 2676 3841
rect 2360 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2676 3840
rect 2360 3775 2676 3776
rect 3303 3840 3619 3841
rect 3303 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3619 3840
rect 3303 3775 3619 3776
rect 4246 3840 4562 3841
rect 4246 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4562 3840
rect 4246 3775 4562 3776
rect 1888 3296 2204 3297
rect 1888 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2204 3296
rect 1888 3231 2204 3232
rect 2831 3296 3147 3297
rect 2831 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3147 3296
rect 2831 3231 3147 3232
rect 3774 3296 4090 3297
rect 3774 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4090 3296
rect 3774 3231 4090 3232
rect 4717 3296 5033 3297
rect 4717 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5033 3296
rect 4717 3231 5033 3232
rect 1417 2752 1733 2753
rect 1417 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1733 2752
rect 1417 2687 1733 2688
rect 2360 2752 2676 2753
rect 2360 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2676 2752
rect 2360 2687 2676 2688
rect 3303 2752 3619 2753
rect 3303 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3619 2752
rect 3303 2687 3619 2688
rect 4246 2752 4562 2753
rect 4246 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4562 2752
rect 4246 2687 4562 2688
rect 4889 2546 4955 2549
rect 4889 2544 5458 2546
rect 4889 2488 4894 2544
rect 4950 2488 5458 2544
rect 4889 2486 5458 2488
rect 4889 2483 4955 2486
rect 5398 2304 5458 2486
rect 1888 2208 2204 2209
rect 1888 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2204 2208
rect 1888 2143 2204 2144
rect 2831 2208 3147 2209
rect 2831 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3147 2208
rect 2831 2143 3147 2144
rect 3774 2208 4090 2209
rect 3774 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4090 2208
rect 3774 2143 4090 2144
rect 4717 2208 5033 2209
rect 4717 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5033 2208
rect 5200 2184 6000 2304
rect 4717 2143 5033 2144
<< via3 >>
rect 1423 13628 1487 13632
rect 1423 13572 1427 13628
rect 1427 13572 1483 13628
rect 1483 13572 1487 13628
rect 1423 13568 1487 13572
rect 1503 13628 1567 13632
rect 1503 13572 1507 13628
rect 1507 13572 1563 13628
rect 1563 13572 1567 13628
rect 1503 13568 1567 13572
rect 1583 13628 1647 13632
rect 1583 13572 1587 13628
rect 1587 13572 1643 13628
rect 1643 13572 1647 13628
rect 1583 13568 1647 13572
rect 1663 13628 1727 13632
rect 1663 13572 1667 13628
rect 1667 13572 1723 13628
rect 1723 13572 1727 13628
rect 1663 13568 1727 13572
rect 2366 13628 2430 13632
rect 2366 13572 2370 13628
rect 2370 13572 2426 13628
rect 2426 13572 2430 13628
rect 2366 13568 2430 13572
rect 2446 13628 2510 13632
rect 2446 13572 2450 13628
rect 2450 13572 2506 13628
rect 2506 13572 2510 13628
rect 2446 13568 2510 13572
rect 2526 13628 2590 13632
rect 2526 13572 2530 13628
rect 2530 13572 2586 13628
rect 2586 13572 2590 13628
rect 2526 13568 2590 13572
rect 2606 13628 2670 13632
rect 2606 13572 2610 13628
rect 2610 13572 2666 13628
rect 2666 13572 2670 13628
rect 2606 13568 2670 13572
rect 3309 13628 3373 13632
rect 3309 13572 3313 13628
rect 3313 13572 3369 13628
rect 3369 13572 3373 13628
rect 3309 13568 3373 13572
rect 3389 13628 3453 13632
rect 3389 13572 3393 13628
rect 3393 13572 3449 13628
rect 3449 13572 3453 13628
rect 3389 13568 3453 13572
rect 3469 13628 3533 13632
rect 3469 13572 3473 13628
rect 3473 13572 3529 13628
rect 3529 13572 3533 13628
rect 3469 13568 3533 13572
rect 3549 13628 3613 13632
rect 3549 13572 3553 13628
rect 3553 13572 3609 13628
rect 3609 13572 3613 13628
rect 3549 13568 3613 13572
rect 4252 13628 4316 13632
rect 4252 13572 4256 13628
rect 4256 13572 4312 13628
rect 4312 13572 4316 13628
rect 4252 13568 4316 13572
rect 4332 13628 4396 13632
rect 4332 13572 4336 13628
rect 4336 13572 4392 13628
rect 4392 13572 4396 13628
rect 4332 13568 4396 13572
rect 4412 13628 4476 13632
rect 4412 13572 4416 13628
rect 4416 13572 4472 13628
rect 4472 13572 4476 13628
rect 4412 13568 4476 13572
rect 4492 13628 4556 13632
rect 4492 13572 4496 13628
rect 4496 13572 4552 13628
rect 4552 13572 4556 13628
rect 4492 13568 4556 13572
rect 1894 13084 1958 13088
rect 1894 13028 1898 13084
rect 1898 13028 1954 13084
rect 1954 13028 1958 13084
rect 1894 13024 1958 13028
rect 1974 13084 2038 13088
rect 1974 13028 1978 13084
rect 1978 13028 2034 13084
rect 2034 13028 2038 13084
rect 1974 13024 2038 13028
rect 2054 13084 2118 13088
rect 2054 13028 2058 13084
rect 2058 13028 2114 13084
rect 2114 13028 2118 13084
rect 2054 13024 2118 13028
rect 2134 13084 2198 13088
rect 2134 13028 2138 13084
rect 2138 13028 2194 13084
rect 2194 13028 2198 13084
rect 2134 13024 2198 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 3077 13084 3141 13088
rect 3077 13028 3081 13084
rect 3081 13028 3137 13084
rect 3137 13028 3141 13084
rect 3077 13024 3141 13028
rect 3780 13084 3844 13088
rect 3780 13028 3784 13084
rect 3784 13028 3840 13084
rect 3840 13028 3844 13084
rect 3780 13024 3844 13028
rect 3860 13084 3924 13088
rect 3860 13028 3864 13084
rect 3864 13028 3920 13084
rect 3920 13028 3924 13084
rect 3860 13024 3924 13028
rect 3940 13084 4004 13088
rect 3940 13028 3944 13084
rect 3944 13028 4000 13084
rect 4000 13028 4004 13084
rect 3940 13024 4004 13028
rect 4020 13084 4084 13088
rect 4020 13028 4024 13084
rect 4024 13028 4080 13084
rect 4080 13028 4084 13084
rect 4020 13024 4084 13028
rect 4723 13084 4787 13088
rect 4723 13028 4727 13084
rect 4727 13028 4783 13084
rect 4783 13028 4787 13084
rect 4723 13024 4787 13028
rect 4803 13084 4867 13088
rect 4803 13028 4807 13084
rect 4807 13028 4863 13084
rect 4863 13028 4867 13084
rect 4803 13024 4867 13028
rect 4883 13084 4947 13088
rect 4883 13028 4887 13084
rect 4887 13028 4943 13084
rect 4943 13028 4947 13084
rect 4883 13024 4947 13028
rect 4963 13084 5027 13088
rect 4963 13028 4967 13084
rect 4967 13028 5023 13084
rect 5023 13028 5027 13084
rect 4963 13024 5027 13028
rect 1423 12540 1487 12544
rect 1423 12484 1427 12540
rect 1427 12484 1483 12540
rect 1483 12484 1487 12540
rect 1423 12480 1487 12484
rect 1503 12540 1567 12544
rect 1503 12484 1507 12540
rect 1507 12484 1563 12540
rect 1563 12484 1567 12540
rect 1503 12480 1567 12484
rect 1583 12540 1647 12544
rect 1583 12484 1587 12540
rect 1587 12484 1643 12540
rect 1643 12484 1647 12540
rect 1583 12480 1647 12484
rect 1663 12540 1727 12544
rect 1663 12484 1667 12540
rect 1667 12484 1723 12540
rect 1723 12484 1727 12540
rect 1663 12480 1727 12484
rect 2366 12540 2430 12544
rect 2366 12484 2370 12540
rect 2370 12484 2426 12540
rect 2426 12484 2430 12540
rect 2366 12480 2430 12484
rect 2446 12540 2510 12544
rect 2446 12484 2450 12540
rect 2450 12484 2506 12540
rect 2506 12484 2510 12540
rect 2446 12480 2510 12484
rect 2526 12540 2590 12544
rect 2526 12484 2530 12540
rect 2530 12484 2586 12540
rect 2586 12484 2590 12540
rect 2526 12480 2590 12484
rect 2606 12540 2670 12544
rect 2606 12484 2610 12540
rect 2610 12484 2666 12540
rect 2666 12484 2670 12540
rect 2606 12480 2670 12484
rect 3309 12540 3373 12544
rect 3309 12484 3313 12540
rect 3313 12484 3369 12540
rect 3369 12484 3373 12540
rect 3309 12480 3373 12484
rect 3389 12540 3453 12544
rect 3389 12484 3393 12540
rect 3393 12484 3449 12540
rect 3449 12484 3453 12540
rect 3389 12480 3453 12484
rect 3469 12540 3533 12544
rect 3469 12484 3473 12540
rect 3473 12484 3529 12540
rect 3529 12484 3533 12540
rect 3469 12480 3533 12484
rect 3549 12540 3613 12544
rect 3549 12484 3553 12540
rect 3553 12484 3609 12540
rect 3609 12484 3613 12540
rect 3549 12480 3613 12484
rect 4252 12540 4316 12544
rect 4252 12484 4256 12540
rect 4256 12484 4312 12540
rect 4312 12484 4316 12540
rect 4252 12480 4316 12484
rect 4332 12540 4396 12544
rect 4332 12484 4336 12540
rect 4336 12484 4392 12540
rect 4392 12484 4396 12540
rect 4332 12480 4396 12484
rect 4412 12540 4476 12544
rect 4412 12484 4416 12540
rect 4416 12484 4472 12540
rect 4472 12484 4476 12540
rect 4412 12480 4476 12484
rect 4492 12540 4556 12544
rect 4492 12484 4496 12540
rect 4496 12484 4552 12540
rect 4552 12484 4556 12540
rect 4492 12480 4556 12484
rect 1894 11996 1958 12000
rect 1894 11940 1898 11996
rect 1898 11940 1954 11996
rect 1954 11940 1958 11996
rect 1894 11936 1958 11940
rect 1974 11996 2038 12000
rect 1974 11940 1978 11996
rect 1978 11940 2034 11996
rect 2034 11940 2038 11996
rect 1974 11936 2038 11940
rect 2054 11996 2118 12000
rect 2054 11940 2058 11996
rect 2058 11940 2114 11996
rect 2114 11940 2118 11996
rect 2054 11936 2118 11940
rect 2134 11996 2198 12000
rect 2134 11940 2138 11996
rect 2138 11940 2194 11996
rect 2194 11940 2198 11996
rect 2134 11936 2198 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 3077 11996 3141 12000
rect 3077 11940 3081 11996
rect 3081 11940 3137 11996
rect 3137 11940 3141 11996
rect 3077 11936 3141 11940
rect 3780 11996 3844 12000
rect 3780 11940 3784 11996
rect 3784 11940 3840 11996
rect 3840 11940 3844 11996
rect 3780 11936 3844 11940
rect 3860 11996 3924 12000
rect 3860 11940 3864 11996
rect 3864 11940 3920 11996
rect 3920 11940 3924 11996
rect 3860 11936 3924 11940
rect 3940 11996 4004 12000
rect 3940 11940 3944 11996
rect 3944 11940 4000 11996
rect 4000 11940 4004 11996
rect 3940 11936 4004 11940
rect 4020 11996 4084 12000
rect 4020 11940 4024 11996
rect 4024 11940 4080 11996
rect 4080 11940 4084 11996
rect 4020 11936 4084 11940
rect 4723 11996 4787 12000
rect 4723 11940 4727 11996
rect 4727 11940 4783 11996
rect 4783 11940 4787 11996
rect 4723 11936 4787 11940
rect 4803 11996 4867 12000
rect 4803 11940 4807 11996
rect 4807 11940 4863 11996
rect 4863 11940 4867 11996
rect 4803 11936 4867 11940
rect 4883 11996 4947 12000
rect 4883 11940 4887 11996
rect 4887 11940 4943 11996
rect 4943 11940 4947 11996
rect 4883 11936 4947 11940
rect 4963 11996 5027 12000
rect 4963 11940 4967 11996
rect 4967 11940 5023 11996
rect 5023 11940 5027 11996
rect 4963 11936 5027 11940
rect 1423 11452 1487 11456
rect 1423 11396 1427 11452
rect 1427 11396 1483 11452
rect 1483 11396 1487 11452
rect 1423 11392 1487 11396
rect 1503 11452 1567 11456
rect 1503 11396 1507 11452
rect 1507 11396 1563 11452
rect 1563 11396 1567 11452
rect 1503 11392 1567 11396
rect 1583 11452 1647 11456
rect 1583 11396 1587 11452
rect 1587 11396 1643 11452
rect 1643 11396 1647 11452
rect 1583 11392 1647 11396
rect 1663 11452 1727 11456
rect 1663 11396 1667 11452
rect 1667 11396 1723 11452
rect 1723 11396 1727 11452
rect 1663 11392 1727 11396
rect 2366 11452 2430 11456
rect 2366 11396 2370 11452
rect 2370 11396 2426 11452
rect 2426 11396 2430 11452
rect 2366 11392 2430 11396
rect 2446 11452 2510 11456
rect 2446 11396 2450 11452
rect 2450 11396 2506 11452
rect 2506 11396 2510 11452
rect 2446 11392 2510 11396
rect 2526 11452 2590 11456
rect 2526 11396 2530 11452
rect 2530 11396 2586 11452
rect 2586 11396 2590 11452
rect 2526 11392 2590 11396
rect 2606 11452 2670 11456
rect 2606 11396 2610 11452
rect 2610 11396 2666 11452
rect 2666 11396 2670 11452
rect 2606 11392 2670 11396
rect 3309 11452 3373 11456
rect 3309 11396 3313 11452
rect 3313 11396 3369 11452
rect 3369 11396 3373 11452
rect 3309 11392 3373 11396
rect 3389 11452 3453 11456
rect 3389 11396 3393 11452
rect 3393 11396 3449 11452
rect 3449 11396 3453 11452
rect 3389 11392 3453 11396
rect 3469 11452 3533 11456
rect 3469 11396 3473 11452
rect 3473 11396 3529 11452
rect 3529 11396 3533 11452
rect 3469 11392 3533 11396
rect 3549 11452 3613 11456
rect 3549 11396 3553 11452
rect 3553 11396 3609 11452
rect 3609 11396 3613 11452
rect 3549 11392 3613 11396
rect 4252 11452 4316 11456
rect 4252 11396 4256 11452
rect 4256 11396 4312 11452
rect 4312 11396 4316 11452
rect 4252 11392 4316 11396
rect 4332 11452 4396 11456
rect 4332 11396 4336 11452
rect 4336 11396 4392 11452
rect 4392 11396 4396 11452
rect 4332 11392 4396 11396
rect 4412 11452 4476 11456
rect 4412 11396 4416 11452
rect 4416 11396 4472 11452
rect 4472 11396 4476 11452
rect 4412 11392 4476 11396
rect 4492 11452 4556 11456
rect 4492 11396 4496 11452
rect 4496 11396 4552 11452
rect 4552 11396 4556 11452
rect 4492 11392 4556 11396
rect 1894 10908 1958 10912
rect 1894 10852 1898 10908
rect 1898 10852 1954 10908
rect 1954 10852 1958 10908
rect 1894 10848 1958 10852
rect 1974 10908 2038 10912
rect 1974 10852 1978 10908
rect 1978 10852 2034 10908
rect 2034 10852 2038 10908
rect 1974 10848 2038 10852
rect 2054 10908 2118 10912
rect 2054 10852 2058 10908
rect 2058 10852 2114 10908
rect 2114 10852 2118 10908
rect 2054 10848 2118 10852
rect 2134 10908 2198 10912
rect 2134 10852 2138 10908
rect 2138 10852 2194 10908
rect 2194 10852 2198 10908
rect 2134 10848 2198 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 3077 10908 3141 10912
rect 3077 10852 3081 10908
rect 3081 10852 3137 10908
rect 3137 10852 3141 10908
rect 3077 10848 3141 10852
rect 3780 10908 3844 10912
rect 3780 10852 3784 10908
rect 3784 10852 3840 10908
rect 3840 10852 3844 10908
rect 3780 10848 3844 10852
rect 3860 10908 3924 10912
rect 3860 10852 3864 10908
rect 3864 10852 3920 10908
rect 3920 10852 3924 10908
rect 3860 10848 3924 10852
rect 3940 10908 4004 10912
rect 3940 10852 3944 10908
rect 3944 10852 4000 10908
rect 4000 10852 4004 10908
rect 3940 10848 4004 10852
rect 4020 10908 4084 10912
rect 4020 10852 4024 10908
rect 4024 10852 4080 10908
rect 4080 10852 4084 10908
rect 4020 10848 4084 10852
rect 4723 10908 4787 10912
rect 4723 10852 4727 10908
rect 4727 10852 4783 10908
rect 4783 10852 4787 10908
rect 4723 10848 4787 10852
rect 4803 10908 4867 10912
rect 4803 10852 4807 10908
rect 4807 10852 4863 10908
rect 4863 10852 4867 10908
rect 4803 10848 4867 10852
rect 4883 10908 4947 10912
rect 4883 10852 4887 10908
rect 4887 10852 4943 10908
rect 4943 10852 4947 10908
rect 4883 10848 4947 10852
rect 4963 10908 5027 10912
rect 4963 10852 4967 10908
rect 4967 10852 5023 10908
rect 5023 10852 5027 10908
rect 4963 10848 5027 10852
rect 1423 10364 1487 10368
rect 1423 10308 1427 10364
rect 1427 10308 1483 10364
rect 1483 10308 1487 10364
rect 1423 10304 1487 10308
rect 1503 10364 1567 10368
rect 1503 10308 1507 10364
rect 1507 10308 1563 10364
rect 1563 10308 1567 10364
rect 1503 10304 1567 10308
rect 1583 10364 1647 10368
rect 1583 10308 1587 10364
rect 1587 10308 1643 10364
rect 1643 10308 1647 10364
rect 1583 10304 1647 10308
rect 1663 10364 1727 10368
rect 1663 10308 1667 10364
rect 1667 10308 1723 10364
rect 1723 10308 1727 10364
rect 1663 10304 1727 10308
rect 2366 10364 2430 10368
rect 2366 10308 2370 10364
rect 2370 10308 2426 10364
rect 2426 10308 2430 10364
rect 2366 10304 2430 10308
rect 2446 10364 2510 10368
rect 2446 10308 2450 10364
rect 2450 10308 2506 10364
rect 2506 10308 2510 10364
rect 2446 10304 2510 10308
rect 2526 10364 2590 10368
rect 2526 10308 2530 10364
rect 2530 10308 2586 10364
rect 2586 10308 2590 10364
rect 2526 10304 2590 10308
rect 2606 10364 2670 10368
rect 2606 10308 2610 10364
rect 2610 10308 2666 10364
rect 2666 10308 2670 10364
rect 2606 10304 2670 10308
rect 3309 10364 3373 10368
rect 3309 10308 3313 10364
rect 3313 10308 3369 10364
rect 3369 10308 3373 10364
rect 3309 10304 3373 10308
rect 3389 10364 3453 10368
rect 3389 10308 3393 10364
rect 3393 10308 3449 10364
rect 3449 10308 3453 10364
rect 3389 10304 3453 10308
rect 3469 10364 3533 10368
rect 3469 10308 3473 10364
rect 3473 10308 3529 10364
rect 3529 10308 3533 10364
rect 3469 10304 3533 10308
rect 3549 10364 3613 10368
rect 3549 10308 3553 10364
rect 3553 10308 3609 10364
rect 3609 10308 3613 10364
rect 3549 10304 3613 10308
rect 4252 10364 4316 10368
rect 4252 10308 4256 10364
rect 4256 10308 4312 10364
rect 4312 10308 4316 10364
rect 4252 10304 4316 10308
rect 4332 10364 4396 10368
rect 4332 10308 4336 10364
rect 4336 10308 4392 10364
rect 4392 10308 4396 10364
rect 4332 10304 4396 10308
rect 4412 10364 4476 10368
rect 4412 10308 4416 10364
rect 4416 10308 4472 10364
rect 4472 10308 4476 10364
rect 4412 10304 4476 10308
rect 4492 10364 4556 10368
rect 4492 10308 4496 10364
rect 4496 10308 4552 10364
rect 4552 10308 4556 10364
rect 4492 10304 4556 10308
rect 1894 9820 1958 9824
rect 1894 9764 1898 9820
rect 1898 9764 1954 9820
rect 1954 9764 1958 9820
rect 1894 9760 1958 9764
rect 1974 9820 2038 9824
rect 1974 9764 1978 9820
rect 1978 9764 2034 9820
rect 2034 9764 2038 9820
rect 1974 9760 2038 9764
rect 2054 9820 2118 9824
rect 2054 9764 2058 9820
rect 2058 9764 2114 9820
rect 2114 9764 2118 9820
rect 2054 9760 2118 9764
rect 2134 9820 2198 9824
rect 2134 9764 2138 9820
rect 2138 9764 2194 9820
rect 2194 9764 2198 9820
rect 2134 9760 2198 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 3077 9820 3141 9824
rect 3077 9764 3081 9820
rect 3081 9764 3137 9820
rect 3137 9764 3141 9820
rect 3077 9760 3141 9764
rect 3780 9820 3844 9824
rect 3780 9764 3784 9820
rect 3784 9764 3840 9820
rect 3840 9764 3844 9820
rect 3780 9760 3844 9764
rect 3860 9820 3924 9824
rect 3860 9764 3864 9820
rect 3864 9764 3920 9820
rect 3920 9764 3924 9820
rect 3860 9760 3924 9764
rect 3940 9820 4004 9824
rect 3940 9764 3944 9820
rect 3944 9764 4000 9820
rect 4000 9764 4004 9820
rect 3940 9760 4004 9764
rect 4020 9820 4084 9824
rect 4020 9764 4024 9820
rect 4024 9764 4080 9820
rect 4080 9764 4084 9820
rect 4020 9760 4084 9764
rect 4723 9820 4787 9824
rect 4723 9764 4727 9820
rect 4727 9764 4783 9820
rect 4783 9764 4787 9820
rect 4723 9760 4787 9764
rect 4803 9820 4867 9824
rect 4803 9764 4807 9820
rect 4807 9764 4863 9820
rect 4863 9764 4867 9820
rect 4803 9760 4867 9764
rect 4883 9820 4947 9824
rect 4883 9764 4887 9820
rect 4887 9764 4943 9820
rect 4943 9764 4947 9820
rect 4883 9760 4947 9764
rect 4963 9820 5027 9824
rect 4963 9764 4967 9820
rect 4967 9764 5023 9820
rect 5023 9764 5027 9820
rect 4963 9760 5027 9764
rect 1423 9276 1487 9280
rect 1423 9220 1427 9276
rect 1427 9220 1483 9276
rect 1483 9220 1487 9276
rect 1423 9216 1487 9220
rect 1503 9276 1567 9280
rect 1503 9220 1507 9276
rect 1507 9220 1563 9276
rect 1563 9220 1567 9276
rect 1503 9216 1567 9220
rect 1583 9276 1647 9280
rect 1583 9220 1587 9276
rect 1587 9220 1643 9276
rect 1643 9220 1647 9276
rect 1583 9216 1647 9220
rect 1663 9276 1727 9280
rect 1663 9220 1667 9276
rect 1667 9220 1723 9276
rect 1723 9220 1727 9276
rect 1663 9216 1727 9220
rect 2366 9276 2430 9280
rect 2366 9220 2370 9276
rect 2370 9220 2426 9276
rect 2426 9220 2430 9276
rect 2366 9216 2430 9220
rect 2446 9276 2510 9280
rect 2446 9220 2450 9276
rect 2450 9220 2506 9276
rect 2506 9220 2510 9276
rect 2446 9216 2510 9220
rect 2526 9276 2590 9280
rect 2526 9220 2530 9276
rect 2530 9220 2586 9276
rect 2586 9220 2590 9276
rect 2526 9216 2590 9220
rect 2606 9276 2670 9280
rect 2606 9220 2610 9276
rect 2610 9220 2666 9276
rect 2666 9220 2670 9276
rect 2606 9216 2670 9220
rect 3309 9276 3373 9280
rect 3309 9220 3313 9276
rect 3313 9220 3369 9276
rect 3369 9220 3373 9276
rect 3309 9216 3373 9220
rect 3389 9276 3453 9280
rect 3389 9220 3393 9276
rect 3393 9220 3449 9276
rect 3449 9220 3453 9276
rect 3389 9216 3453 9220
rect 3469 9276 3533 9280
rect 3469 9220 3473 9276
rect 3473 9220 3529 9276
rect 3529 9220 3533 9276
rect 3469 9216 3533 9220
rect 3549 9276 3613 9280
rect 3549 9220 3553 9276
rect 3553 9220 3609 9276
rect 3609 9220 3613 9276
rect 3549 9216 3613 9220
rect 4252 9276 4316 9280
rect 4252 9220 4256 9276
rect 4256 9220 4312 9276
rect 4312 9220 4316 9276
rect 4252 9216 4316 9220
rect 4332 9276 4396 9280
rect 4332 9220 4336 9276
rect 4336 9220 4392 9276
rect 4392 9220 4396 9276
rect 4332 9216 4396 9220
rect 4412 9276 4476 9280
rect 4412 9220 4416 9276
rect 4416 9220 4472 9276
rect 4472 9220 4476 9276
rect 4412 9216 4476 9220
rect 4492 9276 4556 9280
rect 4492 9220 4496 9276
rect 4496 9220 4552 9276
rect 4552 9220 4556 9276
rect 4492 9216 4556 9220
rect 1894 8732 1958 8736
rect 1894 8676 1898 8732
rect 1898 8676 1954 8732
rect 1954 8676 1958 8732
rect 1894 8672 1958 8676
rect 1974 8732 2038 8736
rect 1974 8676 1978 8732
rect 1978 8676 2034 8732
rect 2034 8676 2038 8732
rect 1974 8672 2038 8676
rect 2054 8732 2118 8736
rect 2054 8676 2058 8732
rect 2058 8676 2114 8732
rect 2114 8676 2118 8732
rect 2054 8672 2118 8676
rect 2134 8732 2198 8736
rect 2134 8676 2138 8732
rect 2138 8676 2194 8732
rect 2194 8676 2198 8732
rect 2134 8672 2198 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 3077 8732 3141 8736
rect 3077 8676 3081 8732
rect 3081 8676 3137 8732
rect 3137 8676 3141 8732
rect 3077 8672 3141 8676
rect 3780 8732 3844 8736
rect 3780 8676 3784 8732
rect 3784 8676 3840 8732
rect 3840 8676 3844 8732
rect 3780 8672 3844 8676
rect 3860 8732 3924 8736
rect 3860 8676 3864 8732
rect 3864 8676 3920 8732
rect 3920 8676 3924 8732
rect 3860 8672 3924 8676
rect 3940 8732 4004 8736
rect 3940 8676 3944 8732
rect 3944 8676 4000 8732
rect 4000 8676 4004 8732
rect 3940 8672 4004 8676
rect 4020 8732 4084 8736
rect 4020 8676 4024 8732
rect 4024 8676 4080 8732
rect 4080 8676 4084 8732
rect 4020 8672 4084 8676
rect 4723 8732 4787 8736
rect 4723 8676 4727 8732
rect 4727 8676 4783 8732
rect 4783 8676 4787 8732
rect 4723 8672 4787 8676
rect 4803 8732 4867 8736
rect 4803 8676 4807 8732
rect 4807 8676 4863 8732
rect 4863 8676 4867 8732
rect 4803 8672 4867 8676
rect 4883 8732 4947 8736
rect 4883 8676 4887 8732
rect 4887 8676 4943 8732
rect 4943 8676 4947 8732
rect 4883 8672 4947 8676
rect 4963 8732 5027 8736
rect 4963 8676 4967 8732
rect 4967 8676 5023 8732
rect 5023 8676 5027 8732
rect 4963 8672 5027 8676
rect 1423 8188 1487 8192
rect 1423 8132 1427 8188
rect 1427 8132 1483 8188
rect 1483 8132 1487 8188
rect 1423 8128 1487 8132
rect 1503 8188 1567 8192
rect 1503 8132 1507 8188
rect 1507 8132 1563 8188
rect 1563 8132 1567 8188
rect 1503 8128 1567 8132
rect 1583 8188 1647 8192
rect 1583 8132 1587 8188
rect 1587 8132 1643 8188
rect 1643 8132 1647 8188
rect 1583 8128 1647 8132
rect 1663 8188 1727 8192
rect 1663 8132 1667 8188
rect 1667 8132 1723 8188
rect 1723 8132 1727 8188
rect 1663 8128 1727 8132
rect 2366 8188 2430 8192
rect 2366 8132 2370 8188
rect 2370 8132 2426 8188
rect 2426 8132 2430 8188
rect 2366 8128 2430 8132
rect 2446 8188 2510 8192
rect 2446 8132 2450 8188
rect 2450 8132 2506 8188
rect 2506 8132 2510 8188
rect 2446 8128 2510 8132
rect 2526 8188 2590 8192
rect 2526 8132 2530 8188
rect 2530 8132 2586 8188
rect 2586 8132 2590 8188
rect 2526 8128 2590 8132
rect 2606 8188 2670 8192
rect 2606 8132 2610 8188
rect 2610 8132 2666 8188
rect 2666 8132 2670 8188
rect 2606 8128 2670 8132
rect 3309 8188 3373 8192
rect 3309 8132 3313 8188
rect 3313 8132 3369 8188
rect 3369 8132 3373 8188
rect 3309 8128 3373 8132
rect 3389 8188 3453 8192
rect 3389 8132 3393 8188
rect 3393 8132 3449 8188
rect 3449 8132 3453 8188
rect 3389 8128 3453 8132
rect 3469 8188 3533 8192
rect 3469 8132 3473 8188
rect 3473 8132 3529 8188
rect 3529 8132 3533 8188
rect 3469 8128 3533 8132
rect 3549 8188 3613 8192
rect 3549 8132 3553 8188
rect 3553 8132 3609 8188
rect 3609 8132 3613 8188
rect 3549 8128 3613 8132
rect 4252 8188 4316 8192
rect 4252 8132 4256 8188
rect 4256 8132 4312 8188
rect 4312 8132 4316 8188
rect 4252 8128 4316 8132
rect 4332 8188 4396 8192
rect 4332 8132 4336 8188
rect 4336 8132 4392 8188
rect 4392 8132 4396 8188
rect 4332 8128 4396 8132
rect 4412 8188 4476 8192
rect 4412 8132 4416 8188
rect 4416 8132 4472 8188
rect 4472 8132 4476 8188
rect 4412 8128 4476 8132
rect 4492 8188 4556 8192
rect 4492 8132 4496 8188
rect 4496 8132 4552 8188
rect 4552 8132 4556 8188
rect 4492 8128 4556 8132
rect 1894 7644 1958 7648
rect 1894 7588 1898 7644
rect 1898 7588 1954 7644
rect 1954 7588 1958 7644
rect 1894 7584 1958 7588
rect 1974 7644 2038 7648
rect 1974 7588 1978 7644
rect 1978 7588 2034 7644
rect 2034 7588 2038 7644
rect 1974 7584 2038 7588
rect 2054 7644 2118 7648
rect 2054 7588 2058 7644
rect 2058 7588 2114 7644
rect 2114 7588 2118 7644
rect 2054 7584 2118 7588
rect 2134 7644 2198 7648
rect 2134 7588 2138 7644
rect 2138 7588 2194 7644
rect 2194 7588 2198 7644
rect 2134 7584 2198 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 3077 7644 3141 7648
rect 3077 7588 3081 7644
rect 3081 7588 3137 7644
rect 3137 7588 3141 7644
rect 3077 7584 3141 7588
rect 3780 7644 3844 7648
rect 3780 7588 3784 7644
rect 3784 7588 3840 7644
rect 3840 7588 3844 7644
rect 3780 7584 3844 7588
rect 3860 7644 3924 7648
rect 3860 7588 3864 7644
rect 3864 7588 3920 7644
rect 3920 7588 3924 7644
rect 3860 7584 3924 7588
rect 3940 7644 4004 7648
rect 3940 7588 3944 7644
rect 3944 7588 4000 7644
rect 4000 7588 4004 7644
rect 3940 7584 4004 7588
rect 4020 7644 4084 7648
rect 4020 7588 4024 7644
rect 4024 7588 4080 7644
rect 4080 7588 4084 7644
rect 4020 7584 4084 7588
rect 4723 7644 4787 7648
rect 4723 7588 4727 7644
rect 4727 7588 4783 7644
rect 4783 7588 4787 7644
rect 4723 7584 4787 7588
rect 4803 7644 4867 7648
rect 4803 7588 4807 7644
rect 4807 7588 4863 7644
rect 4863 7588 4867 7644
rect 4803 7584 4867 7588
rect 4883 7644 4947 7648
rect 4883 7588 4887 7644
rect 4887 7588 4943 7644
rect 4943 7588 4947 7644
rect 4883 7584 4947 7588
rect 4963 7644 5027 7648
rect 4963 7588 4967 7644
rect 4967 7588 5023 7644
rect 5023 7588 5027 7644
rect 4963 7584 5027 7588
rect 1423 7100 1487 7104
rect 1423 7044 1427 7100
rect 1427 7044 1483 7100
rect 1483 7044 1487 7100
rect 1423 7040 1487 7044
rect 1503 7100 1567 7104
rect 1503 7044 1507 7100
rect 1507 7044 1563 7100
rect 1563 7044 1567 7100
rect 1503 7040 1567 7044
rect 1583 7100 1647 7104
rect 1583 7044 1587 7100
rect 1587 7044 1643 7100
rect 1643 7044 1647 7100
rect 1583 7040 1647 7044
rect 1663 7100 1727 7104
rect 1663 7044 1667 7100
rect 1667 7044 1723 7100
rect 1723 7044 1727 7100
rect 1663 7040 1727 7044
rect 2366 7100 2430 7104
rect 2366 7044 2370 7100
rect 2370 7044 2426 7100
rect 2426 7044 2430 7100
rect 2366 7040 2430 7044
rect 2446 7100 2510 7104
rect 2446 7044 2450 7100
rect 2450 7044 2506 7100
rect 2506 7044 2510 7100
rect 2446 7040 2510 7044
rect 2526 7100 2590 7104
rect 2526 7044 2530 7100
rect 2530 7044 2586 7100
rect 2586 7044 2590 7100
rect 2526 7040 2590 7044
rect 2606 7100 2670 7104
rect 2606 7044 2610 7100
rect 2610 7044 2666 7100
rect 2666 7044 2670 7100
rect 2606 7040 2670 7044
rect 3309 7100 3373 7104
rect 3309 7044 3313 7100
rect 3313 7044 3369 7100
rect 3369 7044 3373 7100
rect 3309 7040 3373 7044
rect 3389 7100 3453 7104
rect 3389 7044 3393 7100
rect 3393 7044 3449 7100
rect 3449 7044 3453 7100
rect 3389 7040 3453 7044
rect 3469 7100 3533 7104
rect 3469 7044 3473 7100
rect 3473 7044 3529 7100
rect 3529 7044 3533 7100
rect 3469 7040 3533 7044
rect 3549 7100 3613 7104
rect 3549 7044 3553 7100
rect 3553 7044 3609 7100
rect 3609 7044 3613 7100
rect 3549 7040 3613 7044
rect 4252 7100 4316 7104
rect 4252 7044 4256 7100
rect 4256 7044 4312 7100
rect 4312 7044 4316 7100
rect 4252 7040 4316 7044
rect 4332 7100 4396 7104
rect 4332 7044 4336 7100
rect 4336 7044 4392 7100
rect 4392 7044 4396 7100
rect 4332 7040 4396 7044
rect 4412 7100 4476 7104
rect 4412 7044 4416 7100
rect 4416 7044 4472 7100
rect 4472 7044 4476 7100
rect 4412 7040 4476 7044
rect 4492 7100 4556 7104
rect 4492 7044 4496 7100
rect 4496 7044 4552 7100
rect 4552 7044 4556 7100
rect 4492 7040 4556 7044
rect 1894 6556 1958 6560
rect 1894 6500 1898 6556
rect 1898 6500 1954 6556
rect 1954 6500 1958 6556
rect 1894 6496 1958 6500
rect 1974 6556 2038 6560
rect 1974 6500 1978 6556
rect 1978 6500 2034 6556
rect 2034 6500 2038 6556
rect 1974 6496 2038 6500
rect 2054 6556 2118 6560
rect 2054 6500 2058 6556
rect 2058 6500 2114 6556
rect 2114 6500 2118 6556
rect 2054 6496 2118 6500
rect 2134 6556 2198 6560
rect 2134 6500 2138 6556
rect 2138 6500 2194 6556
rect 2194 6500 2198 6556
rect 2134 6496 2198 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 3077 6556 3141 6560
rect 3077 6500 3081 6556
rect 3081 6500 3137 6556
rect 3137 6500 3141 6556
rect 3077 6496 3141 6500
rect 3780 6556 3844 6560
rect 3780 6500 3784 6556
rect 3784 6500 3840 6556
rect 3840 6500 3844 6556
rect 3780 6496 3844 6500
rect 3860 6556 3924 6560
rect 3860 6500 3864 6556
rect 3864 6500 3920 6556
rect 3920 6500 3924 6556
rect 3860 6496 3924 6500
rect 3940 6556 4004 6560
rect 3940 6500 3944 6556
rect 3944 6500 4000 6556
rect 4000 6500 4004 6556
rect 3940 6496 4004 6500
rect 4020 6556 4084 6560
rect 4020 6500 4024 6556
rect 4024 6500 4080 6556
rect 4080 6500 4084 6556
rect 4020 6496 4084 6500
rect 4723 6556 4787 6560
rect 4723 6500 4727 6556
rect 4727 6500 4783 6556
rect 4783 6500 4787 6556
rect 4723 6496 4787 6500
rect 4803 6556 4867 6560
rect 4803 6500 4807 6556
rect 4807 6500 4863 6556
rect 4863 6500 4867 6556
rect 4803 6496 4867 6500
rect 4883 6556 4947 6560
rect 4883 6500 4887 6556
rect 4887 6500 4943 6556
rect 4943 6500 4947 6556
rect 4883 6496 4947 6500
rect 4963 6556 5027 6560
rect 4963 6500 4967 6556
rect 4967 6500 5023 6556
rect 5023 6500 5027 6556
rect 4963 6496 5027 6500
rect 1423 6012 1487 6016
rect 1423 5956 1427 6012
rect 1427 5956 1483 6012
rect 1483 5956 1487 6012
rect 1423 5952 1487 5956
rect 1503 6012 1567 6016
rect 1503 5956 1507 6012
rect 1507 5956 1563 6012
rect 1563 5956 1567 6012
rect 1503 5952 1567 5956
rect 1583 6012 1647 6016
rect 1583 5956 1587 6012
rect 1587 5956 1643 6012
rect 1643 5956 1647 6012
rect 1583 5952 1647 5956
rect 1663 6012 1727 6016
rect 1663 5956 1667 6012
rect 1667 5956 1723 6012
rect 1723 5956 1727 6012
rect 1663 5952 1727 5956
rect 2366 6012 2430 6016
rect 2366 5956 2370 6012
rect 2370 5956 2426 6012
rect 2426 5956 2430 6012
rect 2366 5952 2430 5956
rect 2446 6012 2510 6016
rect 2446 5956 2450 6012
rect 2450 5956 2506 6012
rect 2506 5956 2510 6012
rect 2446 5952 2510 5956
rect 2526 6012 2590 6016
rect 2526 5956 2530 6012
rect 2530 5956 2586 6012
rect 2586 5956 2590 6012
rect 2526 5952 2590 5956
rect 2606 6012 2670 6016
rect 2606 5956 2610 6012
rect 2610 5956 2666 6012
rect 2666 5956 2670 6012
rect 2606 5952 2670 5956
rect 3309 6012 3373 6016
rect 3309 5956 3313 6012
rect 3313 5956 3369 6012
rect 3369 5956 3373 6012
rect 3309 5952 3373 5956
rect 3389 6012 3453 6016
rect 3389 5956 3393 6012
rect 3393 5956 3449 6012
rect 3449 5956 3453 6012
rect 3389 5952 3453 5956
rect 3469 6012 3533 6016
rect 3469 5956 3473 6012
rect 3473 5956 3529 6012
rect 3529 5956 3533 6012
rect 3469 5952 3533 5956
rect 3549 6012 3613 6016
rect 3549 5956 3553 6012
rect 3553 5956 3609 6012
rect 3609 5956 3613 6012
rect 3549 5952 3613 5956
rect 4252 6012 4316 6016
rect 4252 5956 4256 6012
rect 4256 5956 4312 6012
rect 4312 5956 4316 6012
rect 4252 5952 4316 5956
rect 4332 6012 4396 6016
rect 4332 5956 4336 6012
rect 4336 5956 4392 6012
rect 4392 5956 4396 6012
rect 4332 5952 4396 5956
rect 4412 6012 4476 6016
rect 4412 5956 4416 6012
rect 4416 5956 4472 6012
rect 4472 5956 4476 6012
rect 4412 5952 4476 5956
rect 4492 6012 4556 6016
rect 4492 5956 4496 6012
rect 4496 5956 4552 6012
rect 4552 5956 4556 6012
rect 4492 5952 4556 5956
rect 1894 5468 1958 5472
rect 1894 5412 1898 5468
rect 1898 5412 1954 5468
rect 1954 5412 1958 5468
rect 1894 5408 1958 5412
rect 1974 5468 2038 5472
rect 1974 5412 1978 5468
rect 1978 5412 2034 5468
rect 2034 5412 2038 5468
rect 1974 5408 2038 5412
rect 2054 5468 2118 5472
rect 2054 5412 2058 5468
rect 2058 5412 2114 5468
rect 2114 5412 2118 5468
rect 2054 5408 2118 5412
rect 2134 5468 2198 5472
rect 2134 5412 2138 5468
rect 2138 5412 2194 5468
rect 2194 5412 2198 5468
rect 2134 5408 2198 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 3077 5468 3141 5472
rect 3077 5412 3081 5468
rect 3081 5412 3137 5468
rect 3137 5412 3141 5468
rect 3077 5408 3141 5412
rect 3780 5468 3844 5472
rect 3780 5412 3784 5468
rect 3784 5412 3840 5468
rect 3840 5412 3844 5468
rect 3780 5408 3844 5412
rect 3860 5468 3924 5472
rect 3860 5412 3864 5468
rect 3864 5412 3920 5468
rect 3920 5412 3924 5468
rect 3860 5408 3924 5412
rect 3940 5468 4004 5472
rect 3940 5412 3944 5468
rect 3944 5412 4000 5468
rect 4000 5412 4004 5468
rect 3940 5408 4004 5412
rect 4020 5468 4084 5472
rect 4020 5412 4024 5468
rect 4024 5412 4080 5468
rect 4080 5412 4084 5468
rect 4020 5408 4084 5412
rect 4723 5468 4787 5472
rect 4723 5412 4727 5468
rect 4727 5412 4783 5468
rect 4783 5412 4787 5468
rect 4723 5408 4787 5412
rect 4803 5468 4867 5472
rect 4803 5412 4807 5468
rect 4807 5412 4863 5468
rect 4863 5412 4867 5468
rect 4803 5408 4867 5412
rect 4883 5468 4947 5472
rect 4883 5412 4887 5468
rect 4887 5412 4943 5468
rect 4943 5412 4947 5468
rect 4883 5408 4947 5412
rect 4963 5468 5027 5472
rect 4963 5412 4967 5468
rect 4967 5412 5023 5468
rect 5023 5412 5027 5468
rect 4963 5408 5027 5412
rect 1423 4924 1487 4928
rect 1423 4868 1427 4924
rect 1427 4868 1483 4924
rect 1483 4868 1487 4924
rect 1423 4864 1487 4868
rect 1503 4924 1567 4928
rect 1503 4868 1507 4924
rect 1507 4868 1563 4924
rect 1563 4868 1567 4924
rect 1503 4864 1567 4868
rect 1583 4924 1647 4928
rect 1583 4868 1587 4924
rect 1587 4868 1643 4924
rect 1643 4868 1647 4924
rect 1583 4864 1647 4868
rect 1663 4924 1727 4928
rect 1663 4868 1667 4924
rect 1667 4868 1723 4924
rect 1723 4868 1727 4924
rect 1663 4864 1727 4868
rect 2366 4924 2430 4928
rect 2366 4868 2370 4924
rect 2370 4868 2426 4924
rect 2426 4868 2430 4924
rect 2366 4864 2430 4868
rect 2446 4924 2510 4928
rect 2446 4868 2450 4924
rect 2450 4868 2506 4924
rect 2506 4868 2510 4924
rect 2446 4864 2510 4868
rect 2526 4924 2590 4928
rect 2526 4868 2530 4924
rect 2530 4868 2586 4924
rect 2586 4868 2590 4924
rect 2526 4864 2590 4868
rect 2606 4924 2670 4928
rect 2606 4868 2610 4924
rect 2610 4868 2666 4924
rect 2666 4868 2670 4924
rect 2606 4864 2670 4868
rect 3309 4924 3373 4928
rect 3309 4868 3313 4924
rect 3313 4868 3369 4924
rect 3369 4868 3373 4924
rect 3309 4864 3373 4868
rect 3389 4924 3453 4928
rect 3389 4868 3393 4924
rect 3393 4868 3449 4924
rect 3449 4868 3453 4924
rect 3389 4864 3453 4868
rect 3469 4924 3533 4928
rect 3469 4868 3473 4924
rect 3473 4868 3529 4924
rect 3529 4868 3533 4924
rect 3469 4864 3533 4868
rect 3549 4924 3613 4928
rect 3549 4868 3553 4924
rect 3553 4868 3609 4924
rect 3609 4868 3613 4924
rect 3549 4864 3613 4868
rect 4252 4924 4316 4928
rect 4252 4868 4256 4924
rect 4256 4868 4312 4924
rect 4312 4868 4316 4924
rect 4252 4864 4316 4868
rect 4332 4924 4396 4928
rect 4332 4868 4336 4924
rect 4336 4868 4392 4924
rect 4392 4868 4396 4924
rect 4332 4864 4396 4868
rect 4412 4924 4476 4928
rect 4412 4868 4416 4924
rect 4416 4868 4472 4924
rect 4472 4868 4476 4924
rect 4412 4864 4476 4868
rect 4492 4924 4556 4928
rect 4492 4868 4496 4924
rect 4496 4868 4552 4924
rect 4552 4868 4556 4924
rect 4492 4864 4556 4868
rect 1894 4380 1958 4384
rect 1894 4324 1898 4380
rect 1898 4324 1954 4380
rect 1954 4324 1958 4380
rect 1894 4320 1958 4324
rect 1974 4380 2038 4384
rect 1974 4324 1978 4380
rect 1978 4324 2034 4380
rect 2034 4324 2038 4380
rect 1974 4320 2038 4324
rect 2054 4380 2118 4384
rect 2054 4324 2058 4380
rect 2058 4324 2114 4380
rect 2114 4324 2118 4380
rect 2054 4320 2118 4324
rect 2134 4380 2198 4384
rect 2134 4324 2138 4380
rect 2138 4324 2194 4380
rect 2194 4324 2198 4380
rect 2134 4320 2198 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 3077 4380 3141 4384
rect 3077 4324 3081 4380
rect 3081 4324 3137 4380
rect 3137 4324 3141 4380
rect 3077 4320 3141 4324
rect 3780 4380 3844 4384
rect 3780 4324 3784 4380
rect 3784 4324 3840 4380
rect 3840 4324 3844 4380
rect 3780 4320 3844 4324
rect 3860 4380 3924 4384
rect 3860 4324 3864 4380
rect 3864 4324 3920 4380
rect 3920 4324 3924 4380
rect 3860 4320 3924 4324
rect 3940 4380 4004 4384
rect 3940 4324 3944 4380
rect 3944 4324 4000 4380
rect 4000 4324 4004 4380
rect 3940 4320 4004 4324
rect 4020 4380 4084 4384
rect 4020 4324 4024 4380
rect 4024 4324 4080 4380
rect 4080 4324 4084 4380
rect 4020 4320 4084 4324
rect 4723 4380 4787 4384
rect 4723 4324 4727 4380
rect 4727 4324 4783 4380
rect 4783 4324 4787 4380
rect 4723 4320 4787 4324
rect 4803 4380 4867 4384
rect 4803 4324 4807 4380
rect 4807 4324 4863 4380
rect 4863 4324 4867 4380
rect 4803 4320 4867 4324
rect 4883 4380 4947 4384
rect 4883 4324 4887 4380
rect 4887 4324 4943 4380
rect 4943 4324 4947 4380
rect 4883 4320 4947 4324
rect 4963 4380 5027 4384
rect 4963 4324 4967 4380
rect 4967 4324 5023 4380
rect 5023 4324 5027 4380
rect 4963 4320 5027 4324
rect 1423 3836 1487 3840
rect 1423 3780 1427 3836
rect 1427 3780 1483 3836
rect 1483 3780 1487 3836
rect 1423 3776 1487 3780
rect 1503 3836 1567 3840
rect 1503 3780 1507 3836
rect 1507 3780 1563 3836
rect 1563 3780 1567 3836
rect 1503 3776 1567 3780
rect 1583 3836 1647 3840
rect 1583 3780 1587 3836
rect 1587 3780 1643 3836
rect 1643 3780 1647 3836
rect 1583 3776 1647 3780
rect 1663 3836 1727 3840
rect 1663 3780 1667 3836
rect 1667 3780 1723 3836
rect 1723 3780 1727 3836
rect 1663 3776 1727 3780
rect 2366 3836 2430 3840
rect 2366 3780 2370 3836
rect 2370 3780 2426 3836
rect 2426 3780 2430 3836
rect 2366 3776 2430 3780
rect 2446 3836 2510 3840
rect 2446 3780 2450 3836
rect 2450 3780 2506 3836
rect 2506 3780 2510 3836
rect 2446 3776 2510 3780
rect 2526 3836 2590 3840
rect 2526 3780 2530 3836
rect 2530 3780 2586 3836
rect 2586 3780 2590 3836
rect 2526 3776 2590 3780
rect 2606 3836 2670 3840
rect 2606 3780 2610 3836
rect 2610 3780 2666 3836
rect 2666 3780 2670 3836
rect 2606 3776 2670 3780
rect 3309 3836 3373 3840
rect 3309 3780 3313 3836
rect 3313 3780 3369 3836
rect 3369 3780 3373 3836
rect 3309 3776 3373 3780
rect 3389 3836 3453 3840
rect 3389 3780 3393 3836
rect 3393 3780 3449 3836
rect 3449 3780 3453 3836
rect 3389 3776 3453 3780
rect 3469 3836 3533 3840
rect 3469 3780 3473 3836
rect 3473 3780 3529 3836
rect 3529 3780 3533 3836
rect 3469 3776 3533 3780
rect 3549 3836 3613 3840
rect 3549 3780 3553 3836
rect 3553 3780 3609 3836
rect 3609 3780 3613 3836
rect 3549 3776 3613 3780
rect 4252 3836 4316 3840
rect 4252 3780 4256 3836
rect 4256 3780 4312 3836
rect 4312 3780 4316 3836
rect 4252 3776 4316 3780
rect 4332 3836 4396 3840
rect 4332 3780 4336 3836
rect 4336 3780 4392 3836
rect 4392 3780 4396 3836
rect 4332 3776 4396 3780
rect 4412 3836 4476 3840
rect 4412 3780 4416 3836
rect 4416 3780 4472 3836
rect 4472 3780 4476 3836
rect 4412 3776 4476 3780
rect 4492 3836 4556 3840
rect 4492 3780 4496 3836
rect 4496 3780 4552 3836
rect 4552 3780 4556 3836
rect 4492 3776 4556 3780
rect 1894 3292 1958 3296
rect 1894 3236 1898 3292
rect 1898 3236 1954 3292
rect 1954 3236 1958 3292
rect 1894 3232 1958 3236
rect 1974 3292 2038 3296
rect 1974 3236 1978 3292
rect 1978 3236 2034 3292
rect 2034 3236 2038 3292
rect 1974 3232 2038 3236
rect 2054 3292 2118 3296
rect 2054 3236 2058 3292
rect 2058 3236 2114 3292
rect 2114 3236 2118 3292
rect 2054 3232 2118 3236
rect 2134 3292 2198 3296
rect 2134 3236 2138 3292
rect 2138 3236 2194 3292
rect 2194 3236 2198 3292
rect 2134 3232 2198 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 3077 3292 3141 3296
rect 3077 3236 3081 3292
rect 3081 3236 3137 3292
rect 3137 3236 3141 3292
rect 3077 3232 3141 3236
rect 3780 3292 3844 3296
rect 3780 3236 3784 3292
rect 3784 3236 3840 3292
rect 3840 3236 3844 3292
rect 3780 3232 3844 3236
rect 3860 3292 3924 3296
rect 3860 3236 3864 3292
rect 3864 3236 3920 3292
rect 3920 3236 3924 3292
rect 3860 3232 3924 3236
rect 3940 3292 4004 3296
rect 3940 3236 3944 3292
rect 3944 3236 4000 3292
rect 4000 3236 4004 3292
rect 3940 3232 4004 3236
rect 4020 3292 4084 3296
rect 4020 3236 4024 3292
rect 4024 3236 4080 3292
rect 4080 3236 4084 3292
rect 4020 3232 4084 3236
rect 4723 3292 4787 3296
rect 4723 3236 4727 3292
rect 4727 3236 4783 3292
rect 4783 3236 4787 3292
rect 4723 3232 4787 3236
rect 4803 3292 4867 3296
rect 4803 3236 4807 3292
rect 4807 3236 4863 3292
rect 4863 3236 4867 3292
rect 4803 3232 4867 3236
rect 4883 3292 4947 3296
rect 4883 3236 4887 3292
rect 4887 3236 4943 3292
rect 4943 3236 4947 3292
rect 4883 3232 4947 3236
rect 4963 3292 5027 3296
rect 4963 3236 4967 3292
rect 4967 3236 5023 3292
rect 5023 3236 5027 3292
rect 4963 3232 5027 3236
rect 1423 2748 1487 2752
rect 1423 2692 1427 2748
rect 1427 2692 1483 2748
rect 1483 2692 1487 2748
rect 1423 2688 1487 2692
rect 1503 2748 1567 2752
rect 1503 2692 1507 2748
rect 1507 2692 1563 2748
rect 1563 2692 1567 2748
rect 1503 2688 1567 2692
rect 1583 2748 1647 2752
rect 1583 2692 1587 2748
rect 1587 2692 1643 2748
rect 1643 2692 1647 2748
rect 1583 2688 1647 2692
rect 1663 2748 1727 2752
rect 1663 2692 1667 2748
rect 1667 2692 1723 2748
rect 1723 2692 1727 2748
rect 1663 2688 1727 2692
rect 2366 2748 2430 2752
rect 2366 2692 2370 2748
rect 2370 2692 2426 2748
rect 2426 2692 2430 2748
rect 2366 2688 2430 2692
rect 2446 2748 2510 2752
rect 2446 2692 2450 2748
rect 2450 2692 2506 2748
rect 2506 2692 2510 2748
rect 2446 2688 2510 2692
rect 2526 2748 2590 2752
rect 2526 2692 2530 2748
rect 2530 2692 2586 2748
rect 2586 2692 2590 2748
rect 2526 2688 2590 2692
rect 2606 2748 2670 2752
rect 2606 2692 2610 2748
rect 2610 2692 2666 2748
rect 2666 2692 2670 2748
rect 2606 2688 2670 2692
rect 3309 2748 3373 2752
rect 3309 2692 3313 2748
rect 3313 2692 3369 2748
rect 3369 2692 3373 2748
rect 3309 2688 3373 2692
rect 3389 2748 3453 2752
rect 3389 2692 3393 2748
rect 3393 2692 3449 2748
rect 3449 2692 3453 2748
rect 3389 2688 3453 2692
rect 3469 2748 3533 2752
rect 3469 2692 3473 2748
rect 3473 2692 3529 2748
rect 3529 2692 3533 2748
rect 3469 2688 3533 2692
rect 3549 2748 3613 2752
rect 3549 2692 3553 2748
rect 3553 2692 3609 2748
rect 3609 2692 3613 2748
rect 3549 2688 3613 2692
rect 4252 2748 4316 2752
rect 4252 2692 4256 2748
rect 4256 2692 4312 2748
rect 4312 2692 4316 2748
rect 4252 2688 4316 2692
rect 4332 2748 4396 2752
rect 4332 2692 4336 2748
rect 4336 2692 4392 2748
rect 4392 2692 4396 2748
rect 4332 2688 4396 2692
rect 4412 2748 4476 2752
rect 4412 2692 4416 2748
rect 4416 2692 4472 2748
rect 4472 2692 4476 2748
rect 4412 2688 4476 2692
rect 4492 2748 4556 2752
rect 4492 2692 4496 2748
rect 4496 2692 4552 2748
rect 4552 2692 4556 2748
rect 4492 2688 4556 2692
rect 1894 2204 1958 2208
rect 1894 2148 1898 2204
rect 1898 2148 1954 2204
rect 1954 2148 1958 2204
rect 1894 2144 1958 2148
rect 1974 2204 2038 2208
rect 1974 2148 1978 2204
rect 1978 2148 2034 2204
rect 2034 2148 2038 2204
rect 1974 2144 2038 2148
rect 2054 2204 2118 2208
rect 2054 2148 2058 2204
rect 2058 2148 2114 2204
rect 2114 2148 2118 2204
rect 2054 2144 2118 2148
rect 2134 2204 2198 2208
rect 2134 2148 2138 2204
rect 2138 2148 2194 2204
rect 2194 2148 2198 2204
rect 2134 2144 2198 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 3077 2204 3141 2208
rect 3077 2148 3081 2204
rect 3081 2148 3137 2204
rect 3137 2148 3141 2204
rect 3077 2144 3141 2148
rect 3780 2204 3844 2208
rect 3780 2148 3784 2204
rect 3784 2148 3840 2204
rect 3840 2148 3844 2204
rect 3780 2144 3844 2148
rect 3860 2204 3924 2208
rect 3860 2148 3864 2204
rect 3864 2148 3920 2204
rect 3920 2148 3924 2204
rect 3860 2144 3924 2148
rect 3940 2204 4004 2208
rect 3940 2148 3944 2204
rect 3944 2148 4000 2204
rect 4000 2148 4004 2204
rect 3940 2144 4004 2148
rect 4020 2204 4084 2208
rect 4020 2148 4024 2204
rect 4024 2148 4080 2204
rect 4080 2148 4084 2204
rect 4020 2144 4084 2148
rect 4723 2204 4787 2208
rect 4723 2148 4727 2204
rect 4727 2148 4783 2204
rect 4783 2148 4787 2204
rect 4723 2144 4787 2148
rect 4803 2204 4867 2208
rect 4803 2148 4807 2204
rect 4807 2148 4863 2204
rect 4863 2148 4867 2204
rect 4803 2144 4867 2148
rect 4883 2204 4947 2208
rect 4883 2148 4887 2204
rect 4887 2148 4943 2204
rect 4943 2148 4947 2204
rect 4883 2144 4947 2148
rect 4963 2204 5027 2208
rect 4963 2148 4967 2204
rect 4967 2148 5023 2204
rect 5023 2148 5027 2204
rect 4963 2144 5027 2148
<< metal4 >>
rect 1415 13632 1735 13648
rect 1415 13568 1423 13632
rect 1487 13568 1503 13632
rect 1567 13568 1583 13632
rect 1647 13568 1663 13632
rect 1727 13568 1735 13632
rect 1415 12544 1735 13568
rect 1415 12480 1423 12544
rect 1487 12480 1503 12544
rect 1567 12480 1583 12544
rect 1647 12480 1663 12544
rect 1727 12480 1735 12544
rect 1415 11456 1735 12480
rect 1415 11392 1423 11456
rect 1487 11392 1503 11456
rect 1567 11392 1583 11456
rect 1647 11392 1663 11456
rect 1727 11392 1735 11456
rect 1415 10368 1735 11392
rect 1415 10304 1423 10368
rect 1487 10304 1503 10368
rect 1567 10304 1583 10368
rect 1647 10304 1663 10368
rect 1727 10304 1735 10368
rect 1415 9280 1735 10304
rect 1415 9216 1423 9280
rect 1487 9216 1503 9280
rect 1567 9216 1583 9280
rect 1647 9216 1663 9280
rect 1727 9216 1735 9280
rect 1415 8192 1735 9216
rect 1415 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1735 8192
rect 1415 7104 1735 8128
rect 1415 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1735 7104
rect 1415 6016 1735 7040
rect 1415 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1735 6016
rect 1415 4928 1735 5952
rect 1415 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1735 4928
rect 1415 3840 1735 4864
rect 1415 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1735 3840
rect 1415 2752 1735 3776
rect 1415 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1735 2752
rect 1415 2128 1735 2688
rect 1886 13088 2206 13648
rect 1886 13024 1894 13088
rect 1958 13024 1974 13088
rect 2038 13024 2054 13088
rect 2118 13024 2134 13088
rect 2198 13024 2206 13088
rect 1886 12000 2206 13024
rect 1886 11936 1894 12000
rect 1958 11936 1974 12000
rect 2038 11936 2054 12000
rect 2118 11936 2134 12000
rect 2198 11936 2206 12000
rect 1886 10912 2206 11936
rect 1886 10848 1894 10912
rect 1958 10848 1974 10912
rect 2038 10848 2054 10912
rect 2118 10848 2134 10912
rect 2198 10848 2206 10912
rect 1886 9824 2206 10848
rect 1886 9760 1894 9824
rect 1958 9760 1974 9824
rect 2038 9760 2054 9824
rect 2118 9760 2134 9824
rect 2198 9760 2206 9824
rect 1886 8736 2206 9760
rect 1886 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2206 8736
rect 1886 7648 2206 8672
rect 1886 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2206 7648
rect 1886 6560 2206 7584
rect 1886 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2206 6560
rect 1886 5472 2206 6496
rect 1886 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2206 5472
rect 1886 4384 2206 5408
rect 1886 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2206 4384
rect 1886 3296 2206 4320
rect 1886 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2206 3296
rect 1886 2208 2206 3232
rect 1886 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2206 2208
rect 1886 2128 2206 2144
rect 2358 13632 2678 13648
rect 2358 13568 2366 13632
rect 2430 13568 2446 13632
rect 2510 13568 2526 13632
rect 2590 13568 2606 13632
rect 2670 13568 2678 13632
rect 2358 12544 2678 13568
rect 2358 12480 2366 12544
rect 2430 12480 2446 12544
rect 2510 12480 2526 12544
rect 2590 12480 2606 12544
rect 2670 12480 2678 12544
rect 2358 11456 2678 12480
rect 2358 11392 2366 11456
rect 2430 11392 2446 11456
rect 2510 11392 2526 11456
rect 2590 11392 2606 11456
rect 2670 11392 2678 11456
rect 2358 10368 2678 11392
rect 2358 10304 2366 10368
rect 2430 10304 2446 10368
rect 2510 10304 2526 10368
rect 2590 10304 2606 10368
rect 2670 10304 2678 10368
rect 2358 9280 2678 10304
rect 2358 9216 2366 9280
rect 2430 9216 2446 9280
rect 2510 9216 2526 9280
rect 2590 9216 2606 9280
rect 2670 9216 2678 9280
rect 2358 8192 2678 9216
rect 2358 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2678 8192
rect 2358 7104 2678 8128
rect 2358 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2678 7104
rect 2358 6016 2678 7040
rect 2358 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2678 6016
rect 2358 4928 2678 5952
rect 2358 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2678 4928
rect 2358 3840 2678 4864
rect 2358 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2678 3840
rect 2358 2752 2678 3776
rect 2358 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2678 2752
rect 2358 2128 2678 2688
rect 2829 13088 3149 13648
rect 2829 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3077 13088
rect 3141 13024 3149 13088
rect 2829 12000 3149 13024
rect 2829 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3077 12000
rect 3141 11936 3149 12000
rect 2829 10912 3149 11936
rect 2829 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3077 10912
rect 3141 10848 3149 10912
rect 2829 9824 3149 10848
rect 2829 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3077 9824
rect 3141 9760 3149 9824
rect 2829 8736 3149 9760
rect 2829 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3149 8736
rect 2829 7648 3149 8672
rect 2829 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3149 7648
rect 2829 6560 3149 7584
rect 2829 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3149 6560
rect 2829 5472 3149 6496
rect 2829 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3149 5472
rect 2829 4384 3149 5408
rect 2829 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3149 4384
rect 2829 3296 3149 4320
rect 2829 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3149 3296
rect 2829 2208 3149 3232
rect 2829 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3149 2208
rect 2829 2128 3149 2144
rect 3301 13632 3621 13648
rect 3301 13568 3309 13632
rect 3373 13568 3389 13632
rect 3453 13568 3469 13632
rect 3533 13568 3549 13632
rect 3613 13568 3621 13632
rect 3301 12544 3621 13568
rect 3301 12480 3309 12544
rect 3373 12480 3389 12544
rect 3453 12480 3469 12544
rect 3533 12480 3549 12544
rect 3613 12480 3621 12544
rect 3301 11456 3621 12480
rect 3301 11392 3309 11456
rect 3373 11392 3389 11456
rect 3453 11392 3469 11456
rect 3533 11392 3549 11456
rect 3613 11392 3621 11456
rect 3301 10368 3621 11392
rect 3301 10304 3309 10368
rect 3373 10304 3389 10368
rect 3453 10304 3469 10368
rect 3533 10304 3549 10368
rect 3613 10304 3621 10368
rect 3301 9280 3621 10304
rect 3301 9216 3309 9280
rect 3373 9216 3389 9280
rect 3453 9216 3469 9280
rect 3533 9216 3549 9280
rect 3613 9216 3621 9280
rect 3301 8192 3621 9216
rect 3301 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3621 8192
rect 3301 7104 3621 8128
rect 3301 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3621 7104
rect 3301 6016 3621 7040
rect 3301 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3621 6016
rect 3301 4928 3621 5952
rect 3301 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3621 4928
rect 3301 3840 3621 4864
rect 3301 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3621 3840
rect 3301 2752 3621 3776
rect 3301 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3621 2752
rect 3301 2128 3621 2688
rect 3772 13088 4092 13648
rect 3772 13024 3780 13088
rect 3844 13024 3860 13088
rect 3924 13024 3940 13088
rect 4004 13024 4020 13088
rect 4084 13024 4092 13088
rect 3772 12000 4092 13024
rect 3772 11936 3780 12000
rect 3844 11936 3860 12000
rect 3924 11936 3940 12000
rect 4004 11936 4020 12000
rect 4084 11936 4092 12000
rect 3772 10912 4092 11936
rect 3772 10848 3780 10912
rect 3844 10848 3860 10912
rect 3924 10848 3940 10912
rect 4004 10848 4020 10912
rect 4084 10848 4092 10912
rect 3772 9824 4092 10848
rect 3772 9760 3780 9824
rect 3844 9760 3860 9824
rect 3924 9760 3940 9824
rect 4004 9760 4020 9824
rect 4084 9760 4092 9824
rect 3772 8736 4092 9760
rect 3772 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4092 8736
rect 3772 7648 4092 8672
rect 3772 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4092 7648
rect 3772 6560 4092 7584
rect 3772 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4092 6560
rect 3772 5472 4092 6496
rect 3772 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4092 5472
rect 3772 4384 4092 5408
rect 3772 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4092 4384
rect 3772 3296 4092 4320
rect 3772 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4092 3296
rect 3772 2208 4092 3232
rect 3772 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4092 2208
rect 3772 2128 4092 2144
rect 4244 13632 4564 13648
rect 4244 13568 4252 13632
rect 4316 13568 4332 13632
rect 4396 13568 4412 13632
rect 4476 13568 4492 13632
rect 4556 13568 4564 13632
rect 4244 12544 4564 13568
rect 4244 12480 4252 12544
rect 4316 12480 4332 12544
rect 4396 12480 4412 12544
rect 4476 12480 4492 12544
rect 4556 12480 4564 12544
rect 4244 11456 4564 12480
rect 4244 11392 4252 11456
rect 4316 11392 4332 11456
rect 4396 11392 4412 11456
rect 4476 11392 4492 11456
rect 4556 11392 4564 11456
rect 4244 10368 4564 11392
rect 4244 10304 4252 10368
rect 4316 10304 4332 10368
rect 4396 10304 4412 10368
rect 4476 10304 4492 10368
rect 4556 10304 4564 10368
rect 4244 9280 4564 10304
rect 4244 9216 4252 9280
rect 4316 9216 4332 9280
rect 4396 9216 4412 9280
rect 4476 9216 4492 9280
rect 4556 9216 4564 9280
rect 4244 8192 4564 9216
rect 4244 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4564 8192
rect 4244 7104 4564 8128
rect 4244 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4564 7104
rect 4244 6016 4564 7040
rect 4244 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4564 6016
rect 4244 4928 4564 5952
rect 4244 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4564 4928
rect 4244 3840 4564 4864
rect 4244 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4564 3840
rect 4244 2752 4564 3776
rect 4244 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4564 2752
rect 4244 2128 4564 2688
rect 4715 13088 5035 13648
rect 4715 13024 4723 13088
rect 4787 13024 4803 13088
rect 4867 13024 4883 13088
rect 4947 13024 4963 13088
rect 5027 13024 5035 13088
rect 4715 12000 5035 13024
rect 4715 11936 4723 12000
rect 4787 11936 4803 12000
rect 4867 11936 4883 12000
rect 4947 11936 4963 12000
rect 5027 11936 5035 12000
rect 4715 10912 5035 11936
rect 4715 10848 4723 10912
rect 4787 10848 4803 10912
rect 4867 10848 4883 10912
rect 4947 10848 4963 10912
rect 5027 10848 5035 10912
rect 4715 9824 5035 10848
rect 4715 9760 4723 9824
rect 4787 9760 4803 9824
rect 4867 9760 4883 9824
rect 4947 9760 4963 9824
rect 5027 9760 5035 9824
rect 4715 8736 5035 9760
rect 4715 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5035 8736
rect 4715 7648 5035 8672
rect 4715 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5035 7648
rect 4715 6560 5035 7584
rect 4715 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5035 6560
rect 4715 5472 5035 6496
rect 4715 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5035 5472
rect 4715 4384 5035 5408
rect 4715 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5035 4384
rect 4715 3296 5035 4320
rect 4715 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5035 3296
rect 4715 2208 5035 3232
rect 4715 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5035 2208
rect 4715 2128 5035 2144
use sky130_fd_sc_hd__dfxtp_1  _0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_35
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_35
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1688980957
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_35
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_37
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_35
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_22
timestamp 1688980957
transform 1 0 3128 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_34
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_21
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  grid_io_left_out_5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
<< labels >>
flabel metal3 s 5200 2184 6000 2304 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 5200 5992 6000 6112 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 gfpga_pad_GPIO_PAD
port 2 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 prog_clk
port 3 nsew signal input
flabel metal3 s 5200 9800 6000 9920 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 4 nsew signal tristate
flabel metal3 s 5200 13608 6000 13728 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_outpad_0_
port 5 nsew signal input
flabel metal4 s 1415 2128 1735 13648 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 2358 2128 2678 13648 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 3301 2128 3621 13648 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 4244 2128 4564 13648 0 FreeSans 1920 90 0 0 vdd
port 6 nsew power bidirectional
flabel metal4 s 1886 2128 2206 13648 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 2829 2128 3149 13648 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 3772 2128 4092 13648 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
flabel metal4 s 4715 2128 5035 13648 0 FreeSans 1920 90 0 0 vss
port 7 nsew ground bidirectional
rlabel metal1 2990 13600 2990 13600 0 vdd
rlabel via1 3069 13056 3069 13056 0 vss
rlabel metal1 4738 2414 4738 2414 0 ccff_head
rlabel metal1 4600 5882 4600 5882 0 ccff_tail
rlabel metal3 1050 13124 1050 13124 0 gfpga_pad_GPIO_PAD
rlabel metal1 4278 2618 4278 2618 0 net1
rlabel metal1 3726 12818 3726 12818 0 net2
rlabel metal1 4600 5678 4600 5678 0 net3
rlabel metal1 2346 12954 2346 12954 0 net4
rlabel metal1 4554 10166 4554 10166 0 net5
rlabel metal3 1234 7956 1234 7956 0 prog_clk
rlabel metal1 4738 13294 4738 13294 0 right_width_0_height_0_subtile_0__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 6000 16000
<< end >>
