magic
tech sky130A
magscale 1 2
timestamp 1707853340
<< obsli1 >>
rect 1104 2159 10856 9809
<< obsm1 >>
rect 566 1980 11118 10124
<< metal2 >>
rect 754 11200 810 12000
rect 2042 11200 2098 12000
rect 3330 11200 3386 12000
rect 4618 11200 4674 12000
rect 5906 11200 5962 12000
rect 7194 11200 7250 12000
rect 8482 11200 8538 12000
rect 9770 11200 9826 12000
rect 11058 11200 11114 12000
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
<< obsm2 >>
rect 572 11144 698 11257
rect 866 11144 1986 11257
rect 2154 11144 3274 11257
rect 3442 11144 4562 11257
rect 4730 11144 5850 11257
rect 6018 11144 7138 11257
rect 7306 11144 8426 11257
rect 8594 11144 9714 11257
rect 9882 11144 11002 11257
rect 572 856 11112 11144
rect 682 800 1710 856
rect 1878 800 2906 856
rect 3074 800 4102 856
rect 4270 800 5298 856
rect 5466 800 6494 856
rect 6662 800 7690 856
rect 7858 800 8886 856
rect 9054 800 10082 856
rect 10250 800 11112 856
<< metal3 >>
rect 0 11160 800 11280
rect 0 10344 800 10464
rect 11200 10344 12000 10464
rect 0 9528 800 9648
rect 11200 9528 12000 9648
rect 0 8712 800 8832
rect 11200 8712 12000 8832
rect 0 7896 800 8016
rect 11200 7896 12000 8016
rect 0 7080 800 7200
rect 11200 7080 12000 7200
rect 0 6264 800 6384
rect 11200 6264 12000 6384
rect 0 5448 800 5568
rect 11200 5448 12000 5568
rect 0 4632 800 4752
rect 11200 4632 12000 4752
rect 0 3816 800 3936
rect 11200 3816 12000 3936
rect 0 3000 800 3120
rect 11200 3000 12000 3120
rect 0 2184 800 2304
rect 11200 2184 12000 2304
rect 0 1368 800 1488
rect 11200 1368 12000 1488
<< obsm3 >>
rect 880 11080 11346 11253
rect 798 10544 11346 11080
rect 880 10264 11120 10544
rect 798 9728 11346 10264
rect 880 9448 11120 9728
rect 798 8912 11346 9448
rect 880 8632 11120 8912
rect 798 8096 11346 8632
rect 880 7816 11120 8096
rect 798 7280 11346 7816
rect 880 7000 11120 7280
rect 798 6464 11346 7000
rect 880 6184 11120 6464
rect 798 5648 11346 6184
rect 880 5368 11120 5648
rect 798 4832 11346 5368
rect 880 4552 11120 4832
rect 798 4016 11346 4552
rect 880 3736 11120 4016
rect 798 3200 11346 3736
rect 880 2920 11120 3200
rect 798 2384 11346 2920
rect 880 2104 11120 2384
rect 798 1568 11346 2104
rect 880 1395 11120 1568
<< metal4 >>
rect 2163 2128 2483 9840
rect 3382 2128 3702 9840
rect 4601 2128 4921 9840
rect 5820 2128 6140 9840
rect 7039 2128 7359 9840
rect 8258 2128 8578 9840
rect 9477 2128 9797 9840
rect 10696 2128 11016 9840
<< labels >>
rlabel metal3 s 11200 9528 12000 9648 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 11200 10344 12000 10464 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 570 0 626 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[1]
port 4 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 chany_bottom_in[2]
port 5 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[3]
port 6 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[4]
port 7 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 chany_bottom_in[5]
port 8 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[6]
port 9 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[7]
port 10 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_in[8]
port 11 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 chany_bottom_out[0]
port 12 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 chany_bottom_out[1]
port 13 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 chany_bottom_out[2]
port 14 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 chany_bottom_out[3]
port 15 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 chany_bottom_out[4]
port 16 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 chany_bottom_out[5]
port 17 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 chany_bottom_out[6]
port 18 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 chany_bottom_out[7]
port 19 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 chany_bottom_out[8]
port 20 nsew signal output
rlabel metal2 s 754 11200 810 12000 6 chany_top_in[0]
port 21 nsew signal input
rlabel metal2 s 2042 11200 2098 12000 6 chany_top_in[1]
port 22 nsew signal input
rlabel metal2 s 3330 11200 3386 12000 6 chany_top_in[2]
port 23 nsew signal input
rlabel metal2 s 4618 11200 4674 12000 6 chany_top_in[3]
port 24 nsew signal input
rlabel metal2 s 5906 11200 5962 12000 6 chany_top_in[4]
port 25 nsew signal input
rlabel metal2 s 7194 11200 7250 12000 6 chany_top_in[5]
port 26 nsew signal input
rlabel metal2 s 8482 11200 8538 12000 6 chany_top_in[6]
port 27 nsew signal input
rlabel metal2 s 9770 11200 9826 12000 6 chany_top_in[7]
port 28 nsew signal input
rlabel metal2 s 11058 11200 11114 12000 6 chany_top_in[8]
port 29 nsew signal input
rlabel metal3 s 11200 1368 12000 1488 6 chany_top_out[0]
port 30 nsew signal output
rlabel metal3 s 11200 2184 12000 2304 6 chany_top_out[1]
port 31 nsew signal output
rlabel metal3 s 11200 3000 12000 3120 6 chany_top_out[2]
port 32 nsew signal output
rlabel metal3 s 11200 3816 12000 3936 6 chany_top_out[3]
port 33 nsew signal output
rlabel metal3 s 11200 4632 12000 4752 6 chany_top_out[4]
port 34 nsew signal output
rlabel metal3 s 11200 5448 12000 5568 6 chany_top_out[5]
port 35 nsew signal output
rlabel metal3 s 11200 6264 12000 6384 6 chany_top_out[6]
port 36 nsew signal output
rlabel metal3 s 11200 7080 12000 7200 6 chany_top_out[7]
port 37 nsew signal output
rlabel metal3 s 11200 7896 12000 8016 6 chany_top_out[8]
port 38 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 39 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 40 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 41 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 prog_clk
port 42 nsew signal input
rlabel metal3 s 11200 8712 12000 8832 6 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
port 43 nsew signal output
rlabel metal4 s 2163 2128 2483 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 9840 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 3382 2128 3702 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 5820 2128 6140 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 8258 2128 8578 9840 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 10696 2128 11016 9840 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 435462
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/cby_8__1_/runs/24_02_13_13_41/results/signoff/cby_8__1_.magic.gds
string GDS_START 102558
<< end >>

