* NGSPICE file created from sb_8__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

.subckt sb_8__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_out[0]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_ prog_clk top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ vdd vss
XFILLER_0_7_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_062_ net20 vss vss vdd vdd mux_left_track_3.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_9_16 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_045_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_106 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_028_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _023_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_62 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput42 net42 vss vss vdd vdd chany_top_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 vss vss vdd vdd chanx_left_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_061_ net19 vss vss vdd vdd mux_left_track_3.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_9_28 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_044_ _005_ vss vss vdd vdd _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_12_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput32 net32 vss vss vdd vdd chanx_left_out[7] sky130_fd_sc_hd__clkbuf_4
X_098__45 vss vss vdd vdd net45 _098__45/LO sky130_fd_sc_hd__conb_1
XFILLER_0_1_110 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_13_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_060_ mux_left_track_3.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net26 sky130_fd_sc_hd__inv_2
XFILLER_0_10_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_043_ mem_left_track_1.DFF_0_.D vss vss vdd vdd _005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_12_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
Xoutput33 net33 vss vss vdd vdd chanx_left_out[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_13_21 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_19_75 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_19_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_042_ _004_ vss vss vdd vdd _013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput34 net34 vss vss vdd vdd chany_top_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_33 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_0_8 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_19_87 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_19_129 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_041_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_21 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_132 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_15_143 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput24 net24 vss vss vdd vdd ccff_tail sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 vss vss vdd vdd chany_top_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_7_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_102 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_13_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_4_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_19_99 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_040_ mem_top_track_2.DFF_0_.Q vss vss vdd vdd _014_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_33 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_66 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput25 net25 vss vss vdd vdd chanx_left_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput36 net36 vss vss vdd vdd chany_top_out[2] sky130_fd_sc_hd__clkbuf_4
XPHY_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_7_21 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_099_ mux_left_track_1.INVTX1_1_.out _017_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_78 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_16_68 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput26 net26 vss vss vdd vdd chanx_left_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput37 net37 vss vss vdd vdd chany_top_out[3] sky130_fd_sc_hd__clkbuf_4
XPHY_1 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_33 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_098_ net45 _016_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
XFILLER_0_1_57 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xoutput27 net27 vss vss vdd vdd chanx_left_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_143 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xoutput38 net38 vss vss vdd vdd chany_top_out[4] sky130_fd_sc_hd__clkbuf_4
XPHY_2 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_097_ mux_top_track_2.mux_l1_in_0_.TGATE_0_.out _015_ vss vss vdd vdd mux_top_track_2.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_11_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput28 net28 vss vss vdd vdd chanx_left_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xoutput39 net39 vss vss vdd vdd chany_top_out[5] sky130_fd_sc_hd__clkbuf_4
XPHY_3 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_094__44 vss vss vdd vdd net44 _094__44/LO sky130_fd_sc_hd__conb_1
X_096_ mux_top_track_2.INVTX1_0_.out _014_ vss vss vdd vdd mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_11_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_38 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput29 net29 vss vss vdd vdd chanx_left_out[4] sky130_fd_sc_hd__clkbuf_4
X_079_ net15 vss vss vdd vdd net30 sky130_fd_sc_hd__clkbuf_1
XPHY_4 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_18_135 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_095_ mux_top_track_2.INVTX1_1_.out _013_ vss vss vdd vdd mux_top_track_2.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_078_ net14 vss vss vdd vdd net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_5 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_4_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_094_ net44 _012_ vss vss vdd vdd mux_top_track_2.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_077_ net13 vss vss vdd vdd net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_6 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_19_29 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_093_ net43 _011_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
Xinput1 ccff_head vss vss vdd vdd net1 sky130_fd_sc_hd__clkbuf_1
XTAP_90 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_prog_clk prog_clk vss vss vdd vdd clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_132 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_076_ net12 vss vss vdd vdd net33 sky130_fd_sc_hd__buf_1
XFILLER_0_2_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_103__46 vss vss vdd vdd net46 _103__46/LO sky130_fd_sc_hd__conb_1
XPHY_7 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_059_ net21 vss vss vdd vdd mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_0_17_73 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_132 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_092_ mux_top_track_0.INVTX1_1_.out _010_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_91 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 chanx_left_in[0] vss vss vdd vdd net2 sky130_fd_sc_hd__buf_1
XTAP_80 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_144 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_7_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_11_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_058_ net11 vss vss vdd vdd mux_left_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XPHY_8 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_0_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_100 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_091_ mux_top_track_0.mux_l1_in_0_.TGATE_0_.out _009_ vss vss vdd vdd mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XTAP_92 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[1] vss vss vdd vdd net3 sky130_fd_sc_hd__clkbuf_1
XTAP_70 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_123 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_9 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_057_ mux_left_track_1.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net25 sky130_fd_sc_hd__inv_2
XFILLER_0_5_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_090_ mux_top_track_0.INVTX1_0_.out _008_ vss vss vdd vdd mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XTAP_93 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 chanx_left_in[2] vss vss vdd vdd net4 sky130_fd_sc_hd__clkbuf_1
XTAP_60 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_113 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_2_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_056_ net10 vss vss vdd vdd mux_top_track_2.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_039_ mem_left_track_1.DFF_0_.D vss vss vdd vdd _015_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_124 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_8_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_22 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_5_53 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xinput5 chanx_left_in[3] vss vss vdd vdd net5 sky130_fd_sc_hd__buf_1
XFILLER_0_11_12 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_94 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_11_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_055_ net23 vss vss vdd vdd mux_top_track_2.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_17_77 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_038_ _003_ vss vss vdd vdd _016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_8 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_18_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_21 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_24 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_95 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 chanx_left_in[4] vss vss vdd vdd net6 sky130_fd_sc_hd__buf_1
XTAP_73 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_071_ clknet_1_0__leaf_prog_clk net47 vss vss vdd vdd mem_left_track_3.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xinput20 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net20 sky130_fd_sc_hd__clkbuf_1
X_054_ mux_top_track_2.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net35 sky130_fd_sc_hd__inv_2
X_037_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_17_121 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_5_33 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_36 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_96 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_left_in[5] vss vss vdd vdd net7 sky130_fd_sc_hd__buf_1
XTAP_74 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ clknet_1_0__leaf_prog_clk net48 vss vss vdd vdd net24 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_6_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_053_ mux_top_track_0.mux_l2_in_0_.TGATE_0_.out vss vss vdd vdd net34 sky130_fd_sc_hd__inv_2
Xinput10 chanx_left_in[8] vss vss vdd vdd net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_ vss vss vdd vdd
+ net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_105_ mux_left_track_3.INVTX1_0_.out _023_ vss vss vdd vdd mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_036_ _002_ vss vss vdd vdd _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_093__43 vss vss vdd vdd net43 _093__43/LO sky130_fd_sc_hd__conb_1
XFILLER_0_5_45 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XTAP_97 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_48 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XTAP_75 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 chanx_left_in[6] vss vss vdd vdd net8 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_052_ net22 vss vss vdd vdd mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_0_17_69 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xinput22 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_ vss vss vdd vdd
+ net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 chany_top_in[0] vss vss vdd vdd net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_104_ mux_left_track_3.mux_l1_in_0_.TGATE_0_.out _022_ vss vss vdd vdd mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
X_035_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_117 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_prog_clk clknet_0_prog_clk vss vss vdd vdd clknet_1_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_17_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XTAP_98 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 chanx_left_in[7] vss vss vdd vdd net9 sky130_fd_sc_hd__buf_1
XTAP_43 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
X_051_ net2 vss vss vdd vdd mux_top_track_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xinput23 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ vss vss vdd
+ vdd net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 chany_top_in[1] vss vss vdd vdd net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_37 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_103_ net46 _021_ vss vss vdd vdd mux_left_track_3.mux_l2_in_0_.TGATE_0_.out sky130_fd_sc_hd__ebufn_2
X_034_ mem_left_track_1.DFF_0_.Q vss vss vdd vdd _018_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_107 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_18_80 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_14_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xhold1 mem_left_track_1.DFF_1_.Q vss vss vdd vdd net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_80 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_1_9 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_88 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_119 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_108 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_2_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_050_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _008_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
Xinput13 chany_top_in[2] vss vss vdd vdd net13 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_102_ mux_left_track_3.INVTX1_1_.out _020_ vss vss vdd vdd mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
X_033_ mem_left_track_1.DFF_1_.Q vss vss vdd vdd _019_ sky130_fd_sc_hd__inv_2
Xhold2 mem_left_track_3.DFF_0_.Q vss vss vdd vdd net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_89 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_40 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput14 chany_top_in[3] vss vss vdd vdd net14 sky130_fd_sc_hd__buf_1
X_032_ _001_ vss vss vdd vdd _020_ sky130_fd_sc_hd__clkbuf_1
X_101_ mux_left_track_1.mux_l1_in_0_.TGATE_0_.out _019_ vss vss vdd vdd mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_3_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xhold3 mem_left_track_1.DFF_0_.Q vss vss vdd vdd net49 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_0_60 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_17_104 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XTAP_46 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_41 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_30 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput15 chany_top_in[4] vss vss vdd vdd net15 sky130_fd_sc_hd__buf_1
X_031_ mem_left_track_3.DFF_0_.Q vss vss vdd vdd _001_ sky130_fd_sc_hd__clkbuf_1
X_100_ mux_left_track_1.INVTX1_0_.out _018_ vss vss vdd vdd mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_3_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xhold4 mem_top_track_0.DFF_1_.Q vss vss vdd vdd net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_94 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_47 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_130 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_20 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_31 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput16 chany_top_in[5] vss vss vdd vdd net16 sky130_fd_sc_hd__buf_1
XFILLER_0_2_141 vss vss vdd vdd sky130_fd_sc_hd__decap_4
X_030_ _000_ vss vss vdd vdd _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_85 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_20_63 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xhold5 mem_top_track_0.DFF_0_.Q vss vss vdd vdd net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_0_73 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_9_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_48 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XTAP_59 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_10 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_21 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_32 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
Xinput17 chany_top_in[6] vss vss vdd vdd net17 sky130_fd_sc_hd__buf_1
XFILLER_0_18_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_089_ net9 vss vss vdd vdd net36 sky130_fd_sc_hd__clkbuf_1
Xhold6 mem_left_track_1.DFF_0_.D vss vss vdd vdd net52 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_49 vss vdd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_11 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XPHY_22 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xinput18 chany_top_in[7] vss vss vdd vdd net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_088_ net8 vss vss vdd vdd net37 sky130_fd_sc_hd__buf_1
Xhold7 mem_top_track_2.DFF_0_.Q vss vss vdd vdd net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_54 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_10 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_42 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_9_40 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_12 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_13_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_34 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_23 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
Xinput19 chany_top_in[8] vss vss vdd vdd net19 sky130_fd_sc_hd__buf_1
XFILLER_0_2_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_087_ net7 vss vss vdd vdd net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_9 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_52 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_35 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_13 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_24 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_2_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_086_ net6 vss vss vdd vdd net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_89 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_20_78 vss vss vdd vdd sky130_fd_sc_hd__decap_6
X_069_ clknet_1_0__leaf_prog_clk net52 vss vss vdd vdd mem_left_track_1.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_66 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_0_22 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_16_110 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_13_124 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_36 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_14 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_25 vss vss vdd vdd sky130_fd_sc_hd__decap_3
X_085_ net5 vss vss vdd vdd net40 sky130_fd_sc_hd__clkbuf_1
X_068_ clknet_1_0__leaf_prog_clk net49 vss vss vdd vdd mem_left_track_1.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XPHY_37 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_6_77 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_15 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XPHY_26 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_3_12 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_084_ net4 vss vss vdd vdd net41 sky130_fd_sc_hd__buf_1
XFILLER_0_20_14 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_067_ clknet_1_1__leaf_prog_clk net50 vss vss vdd vdd mem_top_track_2.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_36 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vss vss vdd vdd sky130_fd_sc_hd__decap_4
XPHY_38 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_16 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_27 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_145 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_24 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_083_ net3 vss vss vdd vdd net42 sky130_fd_sc_hd__buf_1
X_066_ clknet_1_1__leaf_prog_clk net53 vss vss vdd vdd mem_left_track_1.DFF_0_.D sky130_fd_sc_hd__dfxtp_1
X_049_ _007_ vss vss vdd vdd _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_15 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_15_48 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_1_90 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_17 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_28 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_13_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_39 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_36 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_082_ net18 vss vss vdd vdd net27 sky130_fd_sc_hd__buf_1
XFILLER_0_18_59 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_18_26 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_065_ clknet_1_1__leaf_prog_clk net1 vss vss vdd vdd mem_top_track_0.DFF_0_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_38 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_19_111 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_048_ mem_top_track_0.DFF_0_.Q vss vss vdd vdd _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_133 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XPHY_18 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XPHY_29 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_10_109 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_3_48 vss vss vdd vdd sky130_fd_sc_hd__decap_8
XFILLER_0_2_139 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vss vss vdd vdd sky130_ef_sc_hd__decap_12
X_081_ net17 vss vss vdd vdd net28 sky130_fd_sc_hd__clkbuf_1
X_064_ clknet_1_1__leaf_prog_clk net51 vss vss vdd vdd mem_top_track_0.DFF_1_.Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_69 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vss vss vdd vdd sky130_fd_sc_hd__fill_1
X_047_ mem_top_track_0.DFF_1_.Q vss vss vdd vdd _009_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_9 vss vss vdd vdd sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XPHY_19 vss vss vdd vdd sky130_fd_sc_hd__decap_3
XFILLER_0_16_82 vss vss vdd vdd sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput40 net40 vss vss vdd vdd chany_top_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_137 vss vss vdd vdd sky130_fd_sc_hd__decap_8
X_080_ net16 vss vss vdd vdd net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_3 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_063_ net24 vss vss vdd vdd _022_ sky130_fd_sc_hd__inv_2
X_046_ _006_ vss vss vdd vdd _011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_138 vss vss vdd vdd sky130_fd_sc_hd__fill_2
X_029_ net24 vss vss vdd vdd _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_27 vss vss vdd vdd sky130_fd_sc_hd__fill_1
XFILLER_0_16_50 vss vss vdd vdd sky130_ef_sc_hd__decap_12
XFILLER_0_16_94 vss vss vdd vdd sky130_ef_sc_hd__decap_12
Xoutput30 net30 vss vss vdd vdd chanx_left_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 vss vss vdd vdd chany_top_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_105 vss vss vdd vdd sky130_fd_sc_hd__decap_6
.ends

