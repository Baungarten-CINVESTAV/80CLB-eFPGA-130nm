magic
tech sky130A
magscale 1 2
timestamp 1707852211
<< viali >>
rect 2697 9673 2731 9707
rect 10241 9673 10275 9707
rect 1593 9605 1627 9639
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3617 9537 3651 9571
rect 4905 9537 4939 9571
rect 6009 9537 6043 9571
rect 7481 9537 7515 9571
rect 8769 9537 8803 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 3433 9401 3467 9435
rect 2329 9333 2363 9367
rect 2973 9333 3007 9367
rect 4721 9333 4755 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 8585 9333 8619 9367
rect 9597 9333 9631 9367
rect 2145 9129 2179 9163
rect 10425 9129 10459 9163
rect 3617 9061 3651 9095
rect 9965 9061 9999 9095
rect 4261 8993 4295 9027
rect 2329 8925 2363 8959
rect 2605 8925 2639 8959
rect 2881 8925 2915 8959
rect 3433 8925 3467 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 1409 8857 1443 8891
rect 1777 8857 1811 8891
rect 2789 8857 2823 8891
rect 2421 8789 2455 8823
rect 3801 8789 3835 8823
rect 4537 8789 4571 8823
rect 9689 8789 9723 8823
rect 3709 8585 3743 8619
rect 7021 8585 7055 8619
rect 9873 8585 9907 8619
rect 1777 8517 1811 8551
rect 6009 8517 6043 8551
rect 7564 8517 7598 8551
rect 2145 8449 2179 8483
rect 4169 8449 4203 8483
rect 4537 8449 4571 8483
rect 4629 8449 4663 8483
rect 7205 8449 7239 8483
rect 9045 8449 9079 8483
rect 9781 8449 9815 8483
rect 10149 8449 10183 8483
rect 4353 8381 4387 8415
rect 5273 8381 5307 8415
rect 5365 8381 5399 8415
rect 5549 8381 5583 8415
rect 7297 8381 7331 8415
rect 1501 8313 1535 8347
rect 1961 8313 1995 8347
rect 8677 8245 8711 8279
rect 8953 8245 8987 8279
rect 10425 8245 10459 8279
rect 5733 8041 5767 8075
rect 5825 8041 5859 8075
rect 3893 7973 3927 8007
rect 6561 7973 6595 8007
rect 7757 7973 7791 8007
rect 9321 7973 9355 8007
rect 4353 7905 4387 7939
rect 7573 7905 7607 7939
rect 8585 7905 8619 7939
rect 8953 7905 8987 7939
rect 1869 7837 1903 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 4261 7837 4295 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 7389 7837 7423 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 9137 7837 9171 7871
rect 10241 7837 10275 7871
rect 4620 7769 4654 7803
rect 2053 7701 2087 7735
rect 3433 7701 3467 7735
rect 4077 7701 4111 7735
rect 6929 7701 6963 7735
rect 10425 7701 10459 7735
rect 4169 7497 4203 7531
rect 4905 7497 4939 7531
rect 6009 7497 6043 7531
rect 7757 7497 7791 7531
rect 7849 7497 7883 7531
rect 8309 7497 8343 7531
rect 8953 7497 8987 7531
rect 10057 7497 10091 7531
rect 10241 7497 10275 7531
rect 1777 7429 1811 7463
rect 5273 7429 5307 7463
rect 2145 7361 2179 7395
rect 3626 7361 3660 7395
rect 3985 7361 4019 7395
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 8033 7361 8067 7395
rect 8125 7361 8159 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10425 7361 10459 7395
rect 3893 7293 3927 7327
rect 4353 7293 4387 7327
rect 5181 7293 5215 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 8769 7293 8803 7327
rect 9413 7293 9447 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 5733 7225 5767 7259
rect 7021 7225 7055 7259
rect 8401 7225 8435 7259
rect 1501 7157 1535 7191
rect 2329 7157 2363 7191
rect 2513 7157 2547 7191
rect 6377 7157 6411 7191
rect 3617 6953 3651 6987
rect 4721 6953 4755 6987
rect 7113 6953 7147 6987
rect 4629 6885 4663 6919
rect 9689 6885 9723 6919
rect 10149 6885 10183 6919
rect 2053 6817 2087 6851
rect 2237 6817 2271 6851
rect 2421 6817 2455 6851
rect 4169 6817 4203 6851
rect 7481 6817 7515 6851
rect 9045 6817 9079 6851
rect 2145 6749 2179 6783
rect 3065 6749 3099 6783
rect 3985 6749 4019 6783
rect 4905 6749 4939 6783
rect 7021 6749 7055 6783
rect 7573 6749 7607 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 9229 6749 9263 6783
rect 9781 6749 9815 6783
rect 9965 6749 9999 6783
rect 1409 6681 1443 6715
rect 1777 6681 1811 6715
rect 4997 6681 5031 6715
rect 8769 6681 8803 6715
rect 2881 6613 2915 6647
rect 6285 6613 6319 6647
rect 7665 6613 7699 6647
rect 3893 6409 3927 6443
rect 4813 6409 4847 6443
rect 9873 6341 9907 6375
rect 9965 6341 9999 6375
rect 1685 6273 1719 6307
rect 2513 6273 2547 6307
rect 3433 6273 3467 6307
rect 4629 6273 4663 6307
rect 5926 6273 5960 6307
rect 6193 6273 6227 6307
rect 6561 6273 6595 6307
rect 6828 6273 6862 6307
rect 8769 6273 8803 6307
rect 9045 6273 9079 6307
rect 10241 6273 10275 6307
rect 1777 6205 1811 6239
rect 1961 6205 1995 6239
rect 2697 6205 2731 6239
rect 3249 6205 3283 6239
rect 4077 6205 4111 6239
rect 8677 6205 8711 6239
rect 9689 6205 9723 6239
rect 2421 6137 2455 6171
rect 7941 6137 7975 6171
rect 8953 6137 8987 6171
rect 10425 6137 10459 6171
rect 1593 6069 1627 6103
rect 3157 6069 3191 6103
rect 8033 6069 8067 6103
rect 9229 6069 9263 6103
rect 1685 5865 1719 5899
rect 3525 5865 3559 5899
rect 5181 5865 5215 5899
rect 9965 5865 9999 5899
rect 10425 5865 10459 5899
rect 2421 5797 2455 5831
rect 3065 5729 3099 5763
rect 6929 5729 6963 5763
rect 7297 5729 7331 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 2605 5661 2639 5695
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 3801 5661 3835 5695
rect 5273 5661 5307 5695
rect 7564 5661 7598 5695
rect 9781 5661 9815 5695
rect 10241 5661 10275 5695
rect 4068 5593 4102 5627
rect 9045 5593 9079 5627
rect 9137 5593 9171 5627
rect 9689 5593 9723 5627
rect 8677 5525 8711 5559
rect 3065 5321 3099 5355
rect 4445 5321 4479 5355
rect 8953 5321 8987 5355
rect 9689 5321 9723 5355
rect 9965 5321 9999 5355
rect 4353 5253 4387 5287
rect 5457 5253 5491 5287
rect 6009 5253 6043 5287
rect 1593 5185 1627 5219
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 2513 5185 2547 5219
rect 5181 5185 5215 5219
rect 6653 5185 6687 5219
rect 7481 5185 7515 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 4997 5117 5031 5151
rect 5273 5117 5307 5151
rect 6101 5117 6135 5151
rect 7573 5117 7607 5151
rect 7757 5117 7791 5151
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 9045 5117 9079 5151
rect 9229 5117 9263 5151
rect 1409 4981 1443 5015
rect 2329 4981 2363 5015
rect 6469 4981 6503 5015
rect 6837 4981 6871 5015
rect 7941 4981 7975 5015
rect 10425 4981 10459 5015
rect 1501 4777 1535 4811
rect 1961 4777 1995 4811
rect 2421 4777 2455 4811
rect 2973 4777 3007 4811
rect 3801 4777 3835 4811
rect 6285 4777 6319 4811
rect 8309 4777 8343 4811
rect 9321 4777 9355 4811
rect 9965 4777 9999 4811
rect 7941 4709 7975 4743
rect 8401 4709 8435 4743
rect 9689 4709 9723 4743
rect 2789 4641 2823 4675
rect 1777 4573 1811 4607
rect 2145 4573 2179 4607
rect 2513 4573 2547 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3617 4573 3651 4607
rect 5181 4573 5215 4607
rect 5273 4573 5307 4607
rect 5825 4573 5859 4607
rect 6101 4573 6135 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 7113 4573 7147 4607
rect 7297 4573 7331 4607
rect 7849 4573 7883 4607
rect 8125 4573 8159 4607
rect 8585 4573 8619 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 9789 4573 9823 4607
rect 10241 4573 10275 4607
rect 4936 4505 4970 4539
rect 7757 4505 7791 4539
rect 3433 4437 3467 4471
rect 5365 4437 5399 4471
rect 6009 4437 6043 4471
rect 7021 4437 7055 4471
rect 9045 4437 9079 4471
rect 10425 4437 10459 4471
rect 6561 4233 6595 4267
rect 6929 4233 6963 4267
rect 7757 4233 7791 4267
rect 10057 4233 10091 4267
rect 10241 4233 10275 4267
rect 1501 4165 1535 4199
rect 2145 4097 2179 4131
rect 2237 4097 2271 4131
rect 2697 4097 2731 4131
rect 4169 4097 4203 4131
rect 4261 4097 4295 4131
rect 4445 4097 4479 4131
rect 6745 4097 6779 4131
rect 6837 4097 6871 4131
rect 7113 4097 7147 4131
rect 7849 4097 7883 4131
rect 9965 4097 9999 4131
rect 10425 4097 10459 4131
rect 2053 4029 2087 4063
rect 7297 4029 7331 4063
rect 2513 3961 2547 3995
rect 4629 3961 4663 3995
rect 1593 3893 1627 3927
rect 2329 3893 2363 3927
rect 8033 3893 8067 3927
rect 2329 3689 2363 3723
rect 7297 3689 7331 3723
rect 7573 3689 7607 3723
rect 10057 3621 10091 3655
rect 10425 3621 10459 3655
rect 2237 3485 2271 3519
rect 2513 3485 2547 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 9873 3485 9907 3519
rect 10241 3485 10275 3519
rect 1409 3417 1443 3451
rect 1777 3417 1811 3451
rect 2053 3349 2087 3383
rect 3709 3145 3743 3179
rect 10149 3077 10183 3111
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 9597 3009 9631 3043
rect 4353 2805 4387 2839
rect 9781 2805 9815 2839
rect 10425 2805 10459 2839
rect 3249 2601 3283 2635
rect 5641 2601 5675 2635
rect 6837 2601 6871 2635
rect 8033 2601 8067 2635
rect 9229 2601 9263 2635
rect 9597 2601 9631 2635
rect 2053 2533 2087 2567
rect 4445 2533 4479 2567
rect 1409 2397 1443 2431
rect 1869 2397 1903 2431
rect 3065 2397 3099 2431
rect 4261 2397 4295 2431
rect 5457 2397 5491 2431
rect 6653 2397 6687 2431
rect 7849 2397 7883 2431
rect 9045 2397 9079 2431
rect 9413 2397 9447 2431
rect 9689 2397 9723 2431
rect 10149 2397 10183 2431
rect 1593 2261 1627 2295
rect 9873 2261 9907 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 2038 9664 2044 9716
rect 2096 9664 2102 9716
rect 2682 9664 2688 9716
rect 2740 9664 2746 9716
rect 4614 9664 4620 9716
rect 4672 9664 4678 9716
rect 5718 9664 5724 9716
rect 5776 9664 5782 9716
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 8662 9664 8668 9716
rect 8720 9664 8726 9716
rect 9766 9664 9772 9716
rect 9824 9664 9830 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10318 9704 10324 9716
rect 10275 9676 10324 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 2056 9636 2084 9664
rect 2056 9608 3188 9636
rect 750 9528 756 9580
rect 808 9528 814 9580
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 3160 9577 3188 9608
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 2096 9540 2237 9568
rect 2096 9528 2102 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2225 9531 2283 9537
rect 2746 9540 2881 9568
rect 768 9500 796 9528
rect 2746 9500 2774 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9537 3203 9571
rect 3252 9568 3280 9596
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3252 9540 3617 9568
rect 3145 9531 3203 9537
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 4632 9568 4660 9664
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4632 9540 4905 9568
rect 3605 9531 3663 9537
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 5736 9568 5764 9664
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5736 9540 6009 9568
rect 4893 9531 4951 9537
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 7208 9568 7236 9664
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7208 9540 7481 9568
rect 5997 9531 6055 9537
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 8680 9568 8708 9664
rect 9784 9577 9812 9664
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8680 9540 8769 9568
rect 7469 9531 7527 9537
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 768 9472 2774 9500
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 9968 9500 9996 9531
rect 5776 9472 9996 9500
rect 5776 9460 5782 9472
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 1912 9404 2452 9432
rect 1912 9392 1918 9404
rect 1210 9324 1216 9376
rect 1268 9364 1274 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 1268 9336 2329 9364
rect 1268 9324 1274 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2424 9364 2452 9404
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 3421 9435 3479 9441
rect 3421 9432 3433 9435
rect 2556 9404 3433 9432
rect 2556 9392 2562 9404
rect 3421 9401 3433 9404
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 2424 9336 2973 9364
rect 2317 9327 2375 9333
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 2961 9327 3019 9333
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 3936 9336 4721 9364
rect 3936 9324 3942 9336
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6638 9364 6644 9376
rect 6227 9336 6644 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6972 9336 7297 9364
rect 6972 9324 6978 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 8570 9324 8576 9376
rect 8628 9324 8634 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 8720 9336 9597 9364
rect 8720 9324 8726 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 1946 9120 1952 9172
rect 2004 9120 2010 9172
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 2096 9132 2145 9160
rect 2096 9120 2102 9132
rect 2133 9129 2145 9132
rect 2179 9129 2191 9163
rect 8662 9160 8668 9172
rect 2133 9123 2191 9129
rect 2608 9132 8668 9160
rect 1964 9024 1992 9120
rect 1964 8996 2544 9024
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 2516 8888 2544 8996
rect 2608 8965 2636 9132
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 10413 9163 10471 9169
rect 10413 9129 10425 9163
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 3651 9064 4154 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 4126 9024 4154 9064
rect 9048 9064 9965 9092
rect 9048 9036 9076 9064
rect 9953 9061 9965 9064
rect 9999 9061 10011 9095
rect 9953 9055 10011 9061
rect 10428 9036 10456 9123
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4126 8996 4261 9024
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 9030 8984 9036 9036
rect 9088 8984 9094 9036
rect 9876 8996 10364 9024
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3467 8928 4016 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 2777 8891 2835 8897
rect 2777 8888 2789 8891
rect 1811 8860 2452 8888
rect 2516 8860 2789 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 2424 8829 2452 8860
rect 2777 8857 2789 8860
rect 2823 8857 2835 8891
rect 2884 8888 2912 8919
rect 3988 8888 4016 8928
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 5718 8956 5724 8968
rect 4764 8928 5724 8956
rect 4764 8916 4770 8928
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 9876 8965 9904 8996
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10152 8888 10180 8919
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 10336 8956 10364 8996
rect 10410 8984 10416 9036
rect 10468 8984 10474 9036
rect 10594 8956 10600 8968
rect 10336 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11054 8888 11060 8900
rect 2884 8860 3832 8888
rect 3988 8860 4154 8888
rect 10152 8860 11060 8888
rect 2777 8851 2835 8857
rect 3804 8832 3832 8860
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8789 2467 8823
rect 2409 8783 2467 8789
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 4126 8820 4154 8860
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4126 8792 4537 8820
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 9674 8780 9680 8832
rect 9732 8780 9738 8832
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 3786 8616 3792 8628
rect 3743 8588 3792 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 7009 8619 7067 8625
rect 7009 8616 7021 8619
rect 4126 8588 7021 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 4126 8548 4154 8588
rect 7009 8585 7021 8588
rect 7055 8585 7067 8619
rect 7009 8579 7067 8585
rect 9861 8619 9919 8625
rect 9861 8585 9873 8619
rect 9907 8616 9919 8619
rect 10226 8616 10232 8628
rect 9907 8588 10232 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 1811 8520 4154 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 4430 8508 4436 8560
rect 4488 8548 4494 8560
rect 5810 8548 5816 8560
rect 4488 8520 5816 8548
rect 4488 8508 4494 8520
rect 5810 8508 5816 8520
rect 5868 8548 5874 8560
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5868 8520 6009 8548
rect 5868 8508 5874 8520
rect 5997 8517 6009 8520
rect 6043 8517 6055 8551
rect 5997 8511 6055 8517
rect 7552 8551 7610 8557
rect 7552 8517 7564 8551
rect 7598 8548 7610 8551
rect 9674 8548 9680 8560
rect 7598 8520 9680 8548
rect 7598 8517 7610 8520
rect 7552 8511 7610 8517
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 3878 8480 3884 8492
rect 2179 8452 3884 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4203 8452 4537 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4706 8480 4712 8492
rect 4663 8452 4712 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 8662 8480 8668 8492
rect 7239 8452 8668 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9180 8452 9781 8480
rect 9180 8440 9186 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 2314 8372 2320 8424
rect 2372 8372 2378 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8412 4399 8415
rect 4982 8412 4988 8424
rect 4387 8384 4988 8412
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8412 5319 8415
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 5307 8384 5365 8412
rect 5307 8381 5319 8384
rect 5261 8375 5319 8381
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 5353 8375 5411 8381
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 9048 8412 9076 8440
rect 8496 8384 9076 8412
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 1946 8304 1952 8356
rect 2004 8304 2010 8356
rect 2332 8344 2360 8372
rect 2332 8316 4154 8344
rect 4126 8276 4154 8316
rect 8496 8276 8524 8384
rect 4126 8248 8524 8276
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8628 8248 8677 8276
rect 8628 8236 8634 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 8938 8236 8944 8288
rect 8996 8236 9002 8288
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 10502 8276 10508 8288
rect 10459 8248 10508 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1636 8044 5396 8072
rect 1636 8032 1642 8044
rect 3881 8007 3939 8013
rect 3881 7973 3893 8007
rect 3927 8004 3939 8007
rect 4154 8004 4160 8016
rect 3927 7976 4160 8004
rect 3927 7973 3939 7976
rect 3881 7967 3939 7973
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 5368 8004 5396 8044
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 5810 8032 5816 8084
rect 5868 8032 5874 8084
rect 6549 8007 6607 8013
rect 6549 8004 6561 8007
rect 5368 7976 6561 8004
rect 6549 7973 6561 7976
rect 6595 7973 6607 8007
rect 6549 7967 6607 7973
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 7745 8007 7803 8013
rect 7745 8004 7757 8007
rect 6880 7976 7757 8004
rect 6880 7964 6886 7976
rect 7745 7973 7757 7976
rect 7791 7973 7803 8007
rect 7745 7967 7803 7973
rect 9306 7964 9312 8016
rect 9364 7964 9370 8016
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 4028 7908 4353 7936
rect 4028 7896 4034 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 7607 7908 8585 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 8938 7896 8944 7948
rect 8996 7896 9002 7948
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7868 3847 7871
rect 4246 7868 4252 7880
rect 3835 7840 4252 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3620 7800 3648 7831
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 6914 7868 6920 7880
rect 6779 7840 6920 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 4430 7800 4436 7812
rect 3620 7772 4436 7800
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 4608 7803 4666 7809
rect 4608 7769 4620 7803
rect 4654 7800 4666 7803
rect 4890 7800 4896 7812
rect 4654 7772 4896 7800
rect 4654 7769 4666 7772
rect 4608 7763 4666 7769
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 6472 7800 6500 7831
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7834 7868 7840 7880
rect 7423 7840 7840 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7868 8539 7871
rect 8662 7868 8668 7880
rect 8527 7840 8668 7868
rect 8527 7837 8539 7840
rect 8481 7831 8539 7837
rect 8404 7800 8432 7831
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8812 7840 9137 7868
rect 8812 7828 8818 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 8570 7800 8576 7812
rect 6472 7772 6960 7800
rect 8404 7772 8576 7800
rect 2038 7692 2044 7744
rect 2096 7692 2102 7744
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 3421 7735 3479 7741
rect 3421 7732 3433 7735
rect 3292 7704 3433 7732
rect 3292 7692 3298 7704
rect 3421 7701 3433 7704
rect 3467 7701 3479 7735
rect 3421 7695 3479 7701
rect 4062 7692 4068 7744
rect 4120 7692 4126 7744
rect 6932 7741 6960 7772
rect 8570 7760 8576 7772
rect 8628 7800 8634 7812
rect 8628 7772 8708 7800
rect 8628 7760 8634 7772
rect 8680 7744 8708 7772
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7742 7732 7748 7744
rect 6963 7704 7748 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8662 7692 8668 7744
rect 8720 7692 8726 7744
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 1578 7488 1584 7540
rect 1636 7488 1642 7540
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 4062 7488 4068 7540
rect 4120 7488 4126 7540
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 1596 7460 1624 7488
rect 1765 7463 1823 7469
rect 1765 7460 1777 7463
rect 1596 7432 1777 7460
rect 1765 7429 1777 7432
rect 1811 7429 1823 7463
rect 1765 7423 1823 7429
rect 2056 7392 2084 7488
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 2056 7364 2145 7392
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 3602 7352 3608 7404
rect 3660 7401 3666 7404
rect 3660 7355 3672 7401
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4080 7392 4108 7488
rect 4172 7460 4200 7491
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 5534 7528 5540 7540
rect 5000 7500 5540 7528
rect 5000 7460 5028 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6270 7528 6276 7540
rect 6043 7500 6276 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 7834 7488 7840 7540
rect 7892 7488 7898 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8754 7528 8760 7540
rect 8343 7500 8760 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 9306 7528 9312 7540
rect 8987 7500 9312 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10134 7528 10140 7540
rect 10091 7500 10140 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10226 7488 10232 7540
rect 10284 7488 10290 7540
rect 4172 7432 5028 7460
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 5350 7460 5356 7472
rect 5307 7432 5356 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 4019 7364 4108 7392
rect 5905 7395 5963 7401
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 3660 7352 3666 7355
rect 3878 7284 3884 7336
rect 3936 7284 3942 7336
rect 4338 7324 4344 7336
rect 4080 7296 4344 7324
rect 2590 7256 2596 7268
rect 2332 7228 2596 7256
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 2332 7197 2360 7228
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 992 7160 1501 7188
rect 992 7148 998 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7157 2375 7191
rect 2317 7151 2375 7157
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 4080 7188 4108 7296
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4580 7296 5181 7324
rect 4580 7284 4586 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5920 7324 5948 7355
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6144 7364 6561 7392
rect 6144 7352 6150 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6914 7392 6920 7404
rect 6871 7364 6920 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7024 7364 8033 7392
rect 5169 7287 5227 7293
rect 5276 7296 5948 7324
rect 5276 7188 5304 7296
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 7024 7265 7052 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8573 7395 8631 7401
rect 8159 7364 8432 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7466 7324 7472 7336
rect 7331 7296 7472 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5684 7228 5733 7256
rect 5684 7216 5690 7228
rect 5721 7225 5733 7228
rect 5767 7256 5779 7259
rect 7009 7259 7067 7265
rect 5767 7228 6914 7256
rect 5767 7225 5779 7228
rect 5721 7219 5779 7225
rect 2547 7160 5304 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 6362 7148 6368 7200
rect 6420 7148 6426 7200
rect 6886 7188 6914 7228
rect 7009 7225 7021 7259
rect 7055 7225 7067 7259
rect 7116 7256 7144 7287
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 7558 7256 7564 7268
rect 7116 7228 7564 7256
rect 7009 7219 7067 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 8404 7265 8432 7364
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8662 7392 8668 7404
rect 8619 7364 8668 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7225 8447 7259
rect 8680 7256 8708 7352
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 9401 7327 9459 7333
rect 9401 7324 9413 7327
rect 8803 7296 9413 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 9401 7293 9413 7296
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9631 7296 9781 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9876 7324 9904 7355
rect 9950 7352 9956 7404
rect 10008 7352 10014 7404
rect 10413 7395 10471 7401
rect 10413 7392 10425 7395
rect 10336 7364 10425 7392
rect 10336 7324 10364 7364
rect 10413 7361 10425 7364
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 9876 7296 10364 7324
rect 9769 7287 9827 7293
rect 10336 7268 10364 7296
rect 8938 7256 8944 7268
rect 8680 7228 8944 7256
rect 8389 7219 8447 7225
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 9122 7216 9128 7268
rect 9180 7216 9186 7268
rect 10318 7216 10324 7268
rect 10376 7216 10382 7268
rect 9140 7188 9168 7216
rect 6886 7160 9168 7188
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 3602 6944 3608 6996
rect 3660 6944 3666 6996
rect 4430 6944 4436 6996
rect 4488 6984 4494 6996
rect 4709 6987 4767 6993
rect 4709 6984 4721 6987
rect 4488 6956 4721 6984
rect 4488 6944 4494 6956
rect 4709 6953 4721 6956
rect 4755 6953 4767 6987
rect 4709 6947 4767 6953
rect 4982 6944 4988 6996
rect 5040 6944 5046 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 7466 6984 7472 6996
rect 7147 6956 7472 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 7558 6944 7564 6996
rect 7616 6944 7622 6996
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 5000 6916 5028 6944
rect 4672 6888 5028 6916
rect 4672 6876 4678 6888
rect 1670 6808 1676 6860
rect 1728 6848 1734 6860
rect 2041 6851 2099 6857
rect 1728 6820 1900 6848
rect 1728 6808 1734 6820
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1397 6715 1455 6721
rect 1397 6712 1409 6715
rect 992 6684 1409 6712
rect 992 6672 998 6684
rect 1397 6681 1409 6684
rect 1443 6681 1455 6715
rect 1397 6675 1455 6681
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 1765 6715 1823 6721
rect 1765 6712 1777 6715
rect 1728 6684 1777 6712
rect 1728 6672 1734 6684
rect 1765 6681 1777 6684
rect 1811 6681 1823 6715
rect 1872 6712 1900 6820
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 2087 6820 2237 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2590 6848 2596 6860
rect 2455 6820 2596 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 6914 6808 6920 6860
rect 6972 6808 6978 6860
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6848 7527 6851
rect 7576 6848 7604 6944
rect 9677 6919 9735 6925
rect 9677 6885 9689 6919
rect 9723 6916 9735 6919
rect 10042 6916 10048 6928
rect 9723 6888 10048 6916
rect 9723 6885 9735 6888
rect 9677 6879 9735 6885
rect 10042 6876 10048 6888
rect 10100 6916 10106 6928
rect 10137 6919 10195 6925
rect 10137 6916 10149 6919
rect 10100 6888 10149 6916
rect 10100 6876 10106 6888
rect 10137 6885 10149 6888
rect 10183 6885 10195 6919
rect 10137 6879 10195 6885
rect 7515 6820 7604 6848
rect 9033 6851 9091 6857
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9306 6848 9312 6860
rect 9079 6820 9312 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 2498 6780 2504 6792
rect 2179 6752 2504 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3068 6712 3096 6743
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4396 6752 4905 6780
rect 4396 6740 4402 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 6932 6780 6960 6808
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6932 6752 7021 6780
rect 4893 6743 4951 6749
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 8297 6783 8355 6789
rect 7607 6752 8156 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 1872 6684 4154 6712
rect 1765 6675 1823 6681
rect 2516 6656 2544 6684
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2866 6604 2872 6656
rect 2924 6604 2930 6656
rect 4126 6644 4154 6684
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4985 6715 5043 6721
rect 4985 6712 4997 6715
rect 4304 6684 4997 6712
rect 4304 6672 4310 6684
rect 4985 6681 4997 6684
rect 5031 6681 5043 6715
rect 4985 6675 5043 6681
rect 8128 6656 8156 6752
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8435 6752 9229 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 8312 6712 8340 6743
rect 8757 6715 8815 6721
rect 8312 6684 8708 6712
rect 8680 6656 8708 6684
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9784 6712 9812 6743
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 8803 6684 9812 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 4798 6644 4804 6656
rect 4126 6616 4804 6644
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 8110 6604 8116 6656
rect 8168 6604 8174 6656
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 2866 6400 2872 6452
rect 2924 6400 2930 6452
rect 3234 6400 3240 6452
rect 3292 6400 3298 6452
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4614 6440 4620 6452
rect 3927 6412 4620 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 7006 6440 7012 6452
rect 4856 6412 7012 6440
rect 4856 6400 4862 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 10042 6440 10048 6452
rect 9968 6412 10048 6440
rect 1578 6332 1584 6384
rect 1636 6372 1642 6384
rect 1636 6344 1716 6372
rect 1636 6332 1642 6344
rect 1688 6313 1716 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 1673 6267 1731 6273
rect 1780 6276 2513 6304
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 1780 6245 1808 6276
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1544 6208 1777 6236
rect 1544 6196 1550 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 1946 6196 1952 6248
rect 2004 6196 2010 6248
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2774 6236 2780 6248
rect 2731 6208 2780 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 2884 6236 2912 6400
rect 3252 6304 3280 6400
rect 6914 6372 6920 6384
rect 6564 6344 6920 6372
rect 6564 6313 6592 6344
rect 6914 6332 6920 6344
rect 6972 6372 6978 6384
rect 7374 6372 7380 6384
rect 6972 6344 7380 6372
rect 6972 6332 6978 6344
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 9858 6332 9864 6384
rect 9916 6332 9922 6384
rect 9968 6381 9996 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 9953 6375 10011 6381
rect 9953 6341 9965 6375
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 6822 6313 6828 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3252 6276 3433 6304
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 5914 6307 5972 6313
rect 5914 6304 5926 6307
rect 4663 6276 5926 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 5914 6273 5926 6276
rect 5960 6273 5972 6307
rect 5914 6267 5972 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6227 6276 6561 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6816 6304 6828 6313
rect 6783 6276 6828 6304
rect 6549 6267 6607 6273
rect 6816 6267 6828 6276
rect 6822 6264 6828 6267
rect 6880 6264 6886 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 8128 6276 8769 6304
rect 8128 6248 8156 6276
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2884 6208 3249 6236
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 5166 6236 5172 6248
rect 4111 6208 5172 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 8110 6196 8116 6248
rect 8168 6196 8174 6248
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9048 6236 9076 6267
rect 10226 6264 10232 6316
rect 10284 6264 10290 6316
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 8720 6208 9076 6236
rect 9416 6208 9689 6236
rect 8720 6196 8726 6208
rect 2409 6171 2467 6177
rect 2409 6137 2421 6171
rect 2455 6168 2467 6171
rect 3970 6168 3976 6180
rect 2455 6140 3976 6168
rect 2455 6137 2467 6140
rect 2409 6131 2467 6137
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 7929 6171 7987 6177
rect 7929 6137 7941 6171
rect 7975 6168 7987 6171
rect 8680 6168 8708 6196
rect 9416 6180 9444 6208
rect 9677 6205 9689 6208
rect 9723 6236 9735 6239
rect 9766 6236 9772 6248
rect 9723 6208 9772 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 7975 6140 8708 6168
rect 8941 6171 8999 6177
rect 7975 6137 7987 6140
rect 7929 6131 7987 6137
rect 8941 6137 8953 6171
rect 8987 6168 8999 6171
rect 9306 6168 9312 6180
rect 8987 6140 9312 6168
rect 8987 6137 8999 6140
rect 8941 6131 8999 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9398 6128 9404 6180
rect 9456 6128 9462 6180
rect 10410 6128 10416 6180
rect 10468 6128 10474 6180
rect 1578 6060 1584 6112
rect 1636 6060 1642 6112
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 4522 6100 4528 6112
rect 3200 6072 4528 6100
rect 3200 6060 3206 6072
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 8018 6060 8024 6112
rect 8076 6060 8082 6112
rect 9214 6060 9220 6112
rect 9272 6060 9278 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2866 5896 2872 5908
rect 1719 5868 2872 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3142 5856 3148 5908
rect 3200 5856 3206 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 5166 5856 5172 5908
rect 5224 5856 5230 5908
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5865 10471 5899
rect 10413 5859 10471 5865
rect 1596 5760 1624 5856
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 3160 5828 3188 5856
rect 2455 5800 3188 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 6972 5732 7297 5760
rect 6972 5720 6978 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 9232 5760 9260 5856
rect 9324 5828 9352 5856
rect 9324 5800 10272 5828
rect 9232 5732 9812 5760
rect 7285 5723 7343 5729
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2593 5695 2651 5701
rect 2087 5664 2544 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 1872 5624 1900 5655
rect 2406 5624 2412 5636
rect 1872 5596 2412 5624
rect 2406 5584 2412 5596
rect 2464 5584 2470 5636
rect 2516 5556 2544 5664
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2823 5664 2881 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 2869 5661 2881 5664
rect 2915 5692 2927 5695
rect 3789 5695 3847 5701
rect 2915 5664 3372 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2608 5624 2636 5655
rect 3344 5624 3372 5664
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 3878 5692 3884 5704
rect 3835 5664 3884 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4338 5692 4344 5704
rect 3988 5664 4344 5692
rect 3988 5624 4016 5664
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 6270 5692 6276 5704
rect 5316 5664 6276 5692
rect 5316 5652 5322 5664
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 7552 5695 7610 5701
rect 7552 5661 7564 5695
rect 7598 5692 7610 5695
rect 8018 5692 8024 5704
rect 7598 5664 8024 5692
rect 7598 5661 7610 5664
rect 7552 5655 7610 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 9784 5701 9812 5732
rect 10244 5701 10272 5800
rect 10428 5772 10456 5859
rect 10410 5720 10416 5772
rect 10468 5720 10474 5772
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 2608 5596 2912 5624
rect 3344 5596 4016 5624
rect 4056 5627 4114 5633
rect 2774 5556 2780 5568
rect 2516 5528 2780 5556
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 2884 5556 2912 5596
rect 4056 5593 4068 5627
rect 4102 5624 4114 5627
rect 4430 5624 4436 5636
rect 4102 5596 4436 5624
rect 4102 5593 4114 5596
rect 4056 5587 4114 5593
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 9030 5584 9036 5636
rect 9088 5584 9094 5636
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 9456 5596 9689 5624
rect 9456 5584 9462 5596
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9677 5587 9735 5593
rect 4522 5556 4528 5568
rect 2884 5528 4528 5556
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 7524 5528 8677 5556
rect 7524 5516 7530 5528
rect 8665 5525 8677 5528
rect 8711 5556 8723 5559
rect 8846 5556 8852 5568
rect 8711 5528 8852 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1854 5312 1860 5364
rect 1912 5312 1918 5364
rect 2498 5312 2504 5364
rect 2556 5312 2562 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3878 5352 3884 5364
rect 3099 5324 3884 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 4430 5312 4436 5364
rect 4488 5312 4494 5364
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9030 5352 9036 5364
rect 8987 5324 9036 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9030 5312 9036 5324
rect 9088 5352 9094 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9088 5324 9689 5352
rect 9088 5312 9094 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9916 5324 9965 5352
rect 9916 5312 9922 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 1670 5284 1676 5296
rect 1596 5256 1676 5284
rect 1596 5225 1624 5256
rect 1670 5244 1676 5256
rect 1728 5284 1734 5296
rect 1872 5284 1900 5312
rect 1728 5256 1900 5284
rect 1728 5244 1734 5256
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1780 5148 1808 5179
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 2516 5225 2544 5312
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 5258 5284 5264 5296
rect 4387 5256 5264 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5445 5287 5503 5293
rect 5445 5253 5457 5287
rect 5491 5284 5503 5287
rect 5626 5284 5632 5296
rect 5491 5256 5632 5284
rect 5491 5253 5503 5256
rect 5445 5247 5503 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 5997 5287 6055 5293
rect 5997 5253 6009 5287
rect 6043 5284 6055 5287
rect 6362 5284 6368 5296
rect 6043 5256 6368 5284
rect 6043 5253 6055 5256
rect 5997 5247 6055 5253
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 7650 5284 7656 5296
rect 6840 5256 7656 5284
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 1912 5188 2145 5216
rect 1912 5176 1918 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2774 5216 2780 5228
rect 2547 5188 2780 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6512 5188 6653 5216
rect 6512 5176 6518 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 992 5120 1808 5148
rect 992 5108 998 5120
rect 4982 5108 4988 5160
rect 5040 5108 5046 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5350 5148 5356 5160
rect 5307 5120 5356 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6840 5148 6868 5256
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 10134 5176 10140 5228
rect 10192 5176 10198 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 6135 5120 6868 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 7558 5108 7564 5160
rect 7616 5108 7622 5160
rect 7742 5108 7748 5160
rect 7800 5108 7806 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7944 5120 8309 5148
rect 7944 5024 7972 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 8478 5108 8484 5160
rect 8536 5108 8542 5160
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 10244 5148 10272 5179
rect 9916 5120 10272 5148
rect 9916 5108 9922 5120
rect 1394 4972 1400 5024
rect 1452 4972 1458 5024
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2317 5015 2375 5021
rect 2317 5012 2329 5015
rect 2096 4984 2329 5012
rect 2096 4972 2102 4984
rect 2317 4981 2329 4984
rect 2363 4981 2375 5015
rect 2317 4975 2375 4981
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6328 4984 6469 5012
rect 6328 4972 6334 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 6822 4972 6828 5024
rect 6880 4972 6886 5024
rect 7926 4972 7932 5024
rect 7984 4972 7990 5024
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1026 4768 1032 4820
rect 1084 4808 1090 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1084 4780 1501 4808
rect 1084 4768 1090 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 1946 4768 1952 4820
rect 2004 4768 2010 4820
rect 2038 4768 2044 4820
rect 2096 4768 2102 4820
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2498 4808 2504 4820
rect 2455 4780 2504 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2774 4808 2780 4820
rect 2746 4768 2780 4808
rect 2832 4768 2838 4820
rect 2866 4768 2872 4820
rect 2924 4768 2930 4820
rect 2958 4768 2964 4820
rect 3016 4768 3022 4820
rect 3789 4811 3847 4817
rect 3789 4777 3801 4811
rect 3835 4808 3847 4811
rect 4982 4808 4988 4820
rect 3835 4780 4988 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 2056 4604 2084 4768
rect 2746 4740 2774 4768
rect 2516 4712 2774 4740
rect 2516 4613 2544 4712
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 2884 4672 2912 4768
rect 2823 4644 2912 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 2056 4576 2145 4604
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2866 4564 2872 4616
rect 2924 4564 2930 4616
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3605 4607 3663 4613
rect 3191 4576 3464 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3436 4477 3464 4576
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3804 4604 3832 4771
rect 4982 4768 4988 4780
rect 5040 4808 5046 4820
rect 6273 4811 6331 4817
rect 5040 4780 5304 4808
rect 5040 4768 5046 4780
rect 3651 4576 3832 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 5276 4613 5304 4780
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 7742 4808 7748 4820
rect 6319 4780 7748 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8478 4808 8484 4820
rect 8343 4780 8484 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9272 4780 9321 4808
rect 9272 4768 9278 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10134 4808 10140 4820
rect 9999 4780 10140 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10226 4768 10232 4820
rect 10284 4768 10290 4820
rect 6730 4740 6736 4752
rect 6472 4712 6736 4740
rect 6472 4684 6500 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 7929 4743 7987 4749
rect 7929 4740 7941 4743
rect 7616 4712 7941 4740
rect 7616 4700 7622 4712
rect 7929 4709 7941 4712
rect 7975 4709 7987 4743
rect 7929 4703 7987 4709
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 10244 4740 10272 4768
rect 9723 4712 10272 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 6454 4672 6460 4684
rect 5828 4644 6460 4672
rect 5828 4613 5856 4644
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6656 4644 7880 4672
rect 6656 4616 6684 4644
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 3936 4576 5181 4604
rect 3936 4564 3942 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6270 4604 6276 4616
rect 6135 4576 6276 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 6546 4564 6552 4616
rect 6604 4564 6610 4616
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7852 4613 7880 4644
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8404 4604 8432 4703
rect 8662 4672 8668 4684
rect 8588 4644 8668 4672
rect 8588 4613 8616 4644
rect 8662 4632 8668 4644
rect 8720 4672 8726 4684
rect 8720 4644 9260 4672
rect 8720 4632 8726 4644
rect 8159 4576 8432 4604
rect 8573 4607 8631 4613
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 4522 4496 4528 4548
rect 4580 4496 4586 4548
rect 4924 4539 4982 4545
rect 4924 4505 4936 4539
rect 4970 4536 4982 4539
rect 6840 4536 6868 4564
rect 4970 4508 6868 4536
rect 4970 4505 4982 4508
rect 4924 4499 4982 4505
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4437 3479 4471
rect 4540 4468 4568 4496
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 4540 4440 5365 4468
rect 3421 4431 3479 4437
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6178 4468 6184 4480
rect 6043 4440 6184 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 7009 4471 7067 4477
rect 7009 4437 7021 4471
rect 7055 4468 7067 4471
rect 7190 4468 7196 4480
rect 7055 4440 7196 4468
rect 7055 4437 7067 4440
rect 7009 4431 7067 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7300 4468 7328 4567
rect 8938 4564 8944 4616
rect 8996 4564 9002 4616
rect 9232 4613 9260 4644
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9490 4564 9496 4616
rect 9548 4564 9554 4616
rect 9766 4564 9772 4616
rect 9824 4613 9830 4616
rect 9824 4604 9835 4613
rect 9824 4576 9869 4604
rect 9824 4567 9835 4576
rect 9824 4564 9830 4567
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 7745 4539 7803 4545
rect 7745 4505 7757 4539
rect 7791 4536 7803 4539
rect 7926 4536 7932 4548
rect 7791 4508 7932 4536
rect 7791 4505 7803 4508
rect 7745 4499 7803 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 7300 4440 9045 4468
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1452 4236 1532 4264
rect 1452 4224 1458 4236
rect 1504 4205 1532 4236
rect 1670 4224 1676 4276
rect 1728 4224 1734 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 6178 4224 6184 4276
rect 6236 4224 6242 4276
rect 6546 4224 6552 4276
rect 6604 4224 6610 4276
rect 6917 4267 6975 4273
rect 6917 4233 6929 4267
rect 6963 4264 6975 4267
rect 7098 4264 7104 4276
rect 6963 4236 7104 4264
rect 6963 4233 6975 4236
rect 6917 4227 6975 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7248 4236 7757 4264
rect 7248 4224 7254 4236
rect 7745 4233 7757 4236
rect 7791 4264 7803 4267
rect 9030 4264 9036 4276
rect 7791 4236 9036 4264
rect 7791 4233 7803 4236
rect 7745 4227 7803 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 9180 4236 10057 4264
rect 9180 4224 9186 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 10045 4227 10103 4233
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4165 1547 4199
rect 1489 4159 1547 4165
rect 1688 4128 1716 4224
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 1688 4100 2145 4128
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4097 2283 4131
rect 2225 4091 2283 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2731 4100 4108 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1544 4032 2053 4060
rect 1544 4020 1550 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2240 4060 2268 4091
rect 4080 4060 4108 4100
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4338 4128 4344 4140
rect 4295 4100 4344 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 5184 4128 5212 4224
rect 4479 4100 5212 4128
rect 6196 4128 6224 4224
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6512 4168 10456 4196
rect 6512 4156 6518 4168
rect 6840 4137 6868 4168
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6196 4100 6745 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 7101 4131 7159 4137
rect 6871 4100 6905 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7558 4128 7564 4140
rect 7147 4100 7564 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 9766 4128 9772 4140
rect 8904 4100 9772 4128
rect 8904 4088 8910 4100
rect 9766 4088 9772 4100
rect 9824 4128 9830 4140
rect 10428 4137 10456 4168
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9824 4100 9965 4128
rect 9824 4088 9830 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 6638 4060 6644 4072
rect 2240 4032 2728 4060
rect 4080 4032 6644 4060
rect 2041 4023 2099 4029
rect 2700 4004 2728 4032
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7374 4060 7380 4072
rect 7331 4032 7380 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 1728 3964 2513 3992
rect 1728 3952 1734 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 2682 3952 2688 4004
rect 2740 3952 2746 4004
rect 4617 3995 4675 4001
rect 4617 3961 4629 3995
rect 4663 3992 4675 3995
rect 5718 3992 5724 4004
rect 4663 3964 5724 3992
rect 4663 3961 4675 3964
rect 4617 3955 4675 3961
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 992 3896 1593 3924
rect 992 3884 998 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 6362 3924 6368 3936
rect 2363 3896 6368 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 9858 3924 9864 3936
rect 8067 3896 9864 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1912 3692 2329 3720
rect 1912 3680 1918 3692
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 2317 3683 2375 3689
rect 2682 3680 2688 3732
rect 2740 3680 2746 3732
rect 7285 3723 7343 3729
rect 7285 3689 7297 3723
rect 7331 3720 7343 3723
rect 7374 3720 7380 3732
rect 7331 3692 7380 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 7558 3680 7564 3732
rect 7616 3680 7622 3732
rect 2700 3584 2728 3680
rect 10045 3655 10103 3661
rect 10045 3621 10057 3655
rect 10091 3621 10103 3655
rect 10045 3615 10103 3621
rect 2240 3556 2728 3584
rect 2240 3525 2268 3556
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2590 3516 2596 3528
rect 2547 3488 2596 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6788 3488 7389 3516
rect 6788 3476 6794 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 992 3420 1409 3448
rect 992 3408 998 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 1397 3411 1455 3417
rect 1765 3451 1823 3457
rect 1765 3417 1777 3451
rect 1811 3417 1823 3451
rect 7668 3448 7696 3479
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 7984 3488 9873 3516
rect 7984 3476 7990 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 10060 3516 10088 3615
rect 10410 3612 10416 3664
rect 10468 3612 10474 3664
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 10060 3488 10241 3516
rect 9861 3479 9919 3485
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 1765 3411 1823 3417
rect 6932 3420 7696 3448
rect 1780 3380 1808 3411
rect 6932 3392 6960 3420
rect 2041 3383 2099 3389
rect 2041 3380 2053 3383
rect 1780 3352 2053 3380
rect 2041 3349 2053 3352
rect 2087 3349 2099 3383
rect 2041 3343 2099 3349
rect 6914 3340 6920 3392
rect 6972 3340 6978 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 3743 3148 4154 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 2884 3040 2912 3136
rect 4126 3108 4154 3148
rect 10137 3111 10195 3117
rect 10137 3108 10149 3111
rect 4126 3080 10149 3108
rect 10137 3077 10149 3080
rect 10183 3077 10195 3111
rect 10137 3071 10195 3077
rect 3234 3040 3240 3052
rect 2884 3012 3240 3040
rect 3234 3000 3240 3012
rect 3292 3040 3298 3052
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3292 3012 3525 3040
rect 3292 3000 3298 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 6972 3012 9597 3040
rect 6972 3000 6978 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 4338 2796 4344 2848
rect 4396 2796 4402 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 9950 2836 9956 2848
rect 9815 2808 9956 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 3234 2592 3240 2644
rect 3292 2592 3298 2644
rect 4338 2592 4344 2644
rect 4396 2592 4402 2644
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 6454 2632 6460 2644
rect 5675 2604 6460 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7834 2632 7840 2644
rect 6871 2604 7840 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 7926 2592 7932 2644
rect 7984 2592 7990 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8110 2632 8116 2644
rect 8067 2604 8116 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9217 2635 9275 2641
rect 9217 2601 9229 2635
rect 9263 2632 9275 2635
rect 9306 2632 9312 2644
rect 9263 2604 9312 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10318 2632 10324 2644
rect 9631 2604 10324 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 4154 2564 4160 2576
rect 2087 2536 4160 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 4356 2496 4384 2592
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2564 4491 2567
rect 7944 2564 7972 2592
rect 4479 2536 7972 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 4356 2468 9720 2496
rect 566 2388 572 2440
rect 624 2428 630 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 624 2400 1409 2428
rect 624 2388 630 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1854 2388 1860 2440
rect 1912 2388 1918 2440
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4338 2428 4344 2440
rect 4295 2400 4344 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9692 2437 9720 2468
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 6914 2360 6920 2372
rect 1596 2332 6920 2360
rect 1596 2301 1624 2332
rect 6914 2320 6920 2332
rect 6972 2320 6978 2372
rect 9416 2360 9444 2391
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 10008 2400 10149 2428
rect 10008 2388 10014 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10042 2360 10048 2372
rect 9416 2332 10048 2360
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 9858 2252 9864 2304
rect 9916 2252 9922 2304
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 10502 2292 10508 2304
rect 10459 2264 10508 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 2044 9664 2096 9716
rect 2688 9707 2740 9716
rect 2688 9673 2697 9707
rect 2697 9673 2731 9707
rect 2731 9673 2740 9707
rect 2688 9664 2740 9673
rect 4620 9664 4672 9716
rect 5724 9664 5776 9716
rect 7196 9664 7248 9716
rect 8668 9664 8720 9716
rect 9772 9664 9824 9716
rect 10324 9664 10376 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 756 9528 808 9580
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2044 9528 2096 9580
rect 3240 9596 3292 9648
rect 5724 9460 5776 9512
rect 1860 9392 1912 9444
rect 1216 9324 1268 9376
rect 2504 9392 2556 9444
rect 3884 9324 3936 9376
rect 6644 9324 6696 9376
rect 6920 9324 6972 9376
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 8668 9324 8720 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 1952 9120 2004 9172
rect 2044 9120 2096 9172
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 940 8848 992 8900
rect 8668 9120 8720 9172
rect 9036 8984 9088 9036
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5724 8916 5776 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10416 8984 10468 9036
rect 10600 8916 10652 8968
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 11060 8848 11112 8900
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 3792 8576 3844 8628
rect 10232 8576 10284 8628
rect 4436 8508 4488 8560
rect 5816 8508 5868 8560
rect 9680 8508 9732 8560
rect 3884 8440 3936 8492
rect 4712 8440 4764 8492
rect 8668 8440 8720 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9128 8440 9180 8492
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 2320 8372 2372 8424
rect 4988 8372 5040 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 8576 8236 8628 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 10508 8236 10560 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 1584 8032 1636 8084
rect 4160 7964 4212 8016
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 6828 7964 6880 8016
rect 9312 8007 9364 8016
rect 9312 7973 9321 8007
rect 9321 7973 9355 8007
rect 9355 7973 9364 8007
rect 9312 7964 9364 7973
rect 3976 7896 4028 7948
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 4436 7760 4488 7812
rect 4896 7760 4948 7812
rect 6920 7828 6972 7880
rect 7840 7828 7892 7880
rect 8668 7828 8720 7880
rect 8760 7828 8812 7880
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 3240 7692 3292 7744
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 8576 7760 8628 7812
rect 7748 7692 7800 7744
rect 8668 7692 8720 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 1584 7488 1636 7540
rect 2044 7488 2096 7540
rect 4068 7488 4120 7540
rect 3608 7395 3660 7404
rect 3608 7361 3626 7395
rect 3626 7361 3660 7395
rect 3608 7352 3660 7361
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 5540 7488 5592 7540
rect 6276 7488 6328 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 8760 7488 8812 7540
rect 9312 7488 9364 7540
rect 10140 7488 10192 7540
rect 10232 7531 10284 7540
rect 10232 7497 10241 7531
rect 10241 7497 10275 7531
rect 10275 7497 10284 7531
rect 10232 7488 10284 7497
rect 5356 7420 5408 7472
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 4344 7327 4396 7336
rect 940 7148 992 7200
rect 2596 7216 2648 7268
rect 4344 7293 4353 7327
rect 4353 7293 4387 7327
rect 4387 7293 4396 7327
rect 4344 7284 4396 7293
rect 4528 7284 4580 7336
rect 6092 7352 6144 7404
rect 6920 7352 6972 7404
rect 5632 7216 5684 7268
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 7472 7284 7524 7336
rect 7564 7216 7616 7268
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 8944 7216 8996 7268
rect 9128 7216 9180 7268
rect 10324 7216 10376 7268
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 4436 6944 4488 6996
rect 4988 6944 5040 6996
rect 7472 6944 7524 6996
rect 7564 6944 7616 6996
rect 4620 6919 4672 6928
rect 4620 6885 4629 6919
rect 4629 6885 4663 6919
rect 4663 6885 4672 6919
rect 4620 6876 4672 6885
rect 1676 6808 1728 6860
rect 940 6672 992 6724
rect 1676 6672 1728 6724
rect 2596 6808 2648 6860
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 6920 6808 6972 6860
rect 10048 6876 10100 6928
rect 9312 6808 9364 6860
rect 2504 6740 2556 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4344 6740 4396 6792
rect 2504 6604 2556 6656
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 4252 6672 4304 6724
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 4804 6604 4856 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 8116 6604 8168 6656
rect 8668 6604 8720 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 2872 6400 2924 6452
rect 3240 6400 3292 6452
rect 4620 6400 4672 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 7012 6400 7064 6452
rect 1584 6332 1636 6384
rect 1492 6196 1544 6248
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 2780 6196 2832 6248
rect 6920 6332 6972 6384
rect 7380 6332 7432 6384
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 10048 6400 10100 6452
rect 6828 6307 6880 6316
rect 6828 6273 6862 6307
rect 6862 6273 6880 6307
rect 6828 6264 6880 6273
rect 5172 6196 5224 6248
rect 8116 6196 8168 6248
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 8668 6196 8720 6205
rect 3976 6128 4028 6180
rect 9772 6196 9824 6248
rect 9312 6128 9364 6180
rect 9404 6128 9456 6180
rect 10416 6171 10468 6180
rect 10416 6137 10425 6171
rect 10425 6137 10459 6171
rect 10459 6137 10468 6171
rect 10416 6128 10468 6137
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 4528 6060 4580 6112
rect 8024 6103 8076 6112
rect 8024 6069 8033 6103
rect 8033 6069 8067 6103
rect 8067 6069 8076 6103
rect 8024 6060 8076 6069
rect 9220 6103 9272 6112
rect 9220 6069 9229 6103
rect 9229 6069 9263 6103
rect 9263 6069 9272 6103
rect 9220 6060 9272 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1584 5856 1636 5908
rect 2872 5856 2924 5908
rect 3148 5856 3200 5908
rect 3976 5856 4028 5908
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 9220 5856 9272 5908
rect 9312 5856 9364 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 2412 5584 2464 5636
rect 3884 5652 3936 5704
rect 4344 5652 4396 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6276 5652 6328 5704
rect 8024 5652 8076 5704
rect 10416 5720 10468 5772
rect 2780 5516 2832 5568
rect 4436 5584 4488 5636
rect 9036 5627 9088 5636
rect 9036 5593 9045 5627
rect 9045 5593 9079 5627
rect 9079 5593 9088 5627
rect 9036 5584 9088 5593
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 9404 5584 9456 5636
rect 4528 5516 4580 5568
rect 7472 5516 7524 5568
rect 8852 5516 8904 5568
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 1860 5312 1912 5364
rect 2504 5312 2556 5364
rect 3884 5312 3936 5364
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 9036 5312 9088 5364
rect 9864 5312 9916 5364
rect 1676 5244 1728 5296
rect 940 5108 992 5160
rect 1860 5176 1912 5228
rect 5264 5244 5316 5296
rect 5632 5244 5684 5296
rect 6368 5244 6420 5296
rect 2780 5176 2832 5228
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 6460 5176 6512 5228
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5356 5108 5408 5160
rect 7656 5244 7708 5296
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 7564 5151 7616 5160
rect 7564 5117 7573 5151
rect 7573 5117 7607 5151
rect 7607 5117 7616 5151
rect 7564 5108 7616 5117
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 9864 5108 9916 5160
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 2044 4972 2096 5024
rect 6276 4972 6328 5024
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 1032 4768 1084 4820
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2044 4768 2096 4820
rect 2504 4768 2556 4820
rect 2780 4768 2832 4820
rect 2872 4768 2924 4820
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 4988 4768 5040 4820
rect 3884 4564 3936 4616
rect 7748 4768 7800 4820
rect 8484 4768 8536 4820
rect 9220 4768 9272 4820
rect 10140 4768 10192 4820
rect 10232 4768 10284 4820
rect 6736 4700 6788 4752
rect 7564 4700 7616 4752
rect 6460 4632 6512 4684
rect 6276 4564 6328 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 6644 4564 6696 4616
rect 6828 4564 6880 4616
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 8668 4632 8720 4684
rect 4528 4496 4580 4548
rect 6184 4428 6236 4480
rect 7196 4428 7248 4480
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9772 4607 9824 4616
rect 9772 4573 9789 4607
rect 9789 4573 9823 4607
rect 9823 4573 9824 4607
rect 9772 4564 9824 4573
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 7932 4496 7984 4548
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1400 4224 1452 4276
rect 1676 4224 1728 4276
rect 5172 4224 5224 4276
rect 6184 4224 6236 4276
rect 6552 4267 6604 4276
rect 6552 4233 6561 4267
rect 6561 4233 6595 4267
rect 6595 4233 6604 4267
rect 6552 4224 6604 4233
rect 7104 4224 7156 4276
rect 7196 4224 7248 4276
rect 9036 4224 9088 4276
rect 9128 4224 9180 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 1492 4020 1544 4072
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4344 4088 4396 4140
rect 6460 4156 6512 4208
rect 7564 4088 7616 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 8852 4088 8904 4140
rect 9772 4088 9824 4140
rect 6644 4020 6696 4072
rect 7380 4020 7432 4072
rect 1676 3952 1728 4004
rect 2688 3952 2740 4004
rect 5724 3952 5776 4004
rect 940 3884 992 3936
rect 6368 3884 6420 3936
rect 9864 3884 9916 3936
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 1860 3680 1912 3732
rect 2688 3680 2740 3732
rect 7380 3680 7432 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 2596 3476 2648 3528
rect 6736 3476 6788 3528
rect 940 3408 992 3460
rect 7932 3476 7984 3528
rect 10416 3655 10468 3664
rect 10416 3621 10425 3655
rect 10425 3621 10459 3655
rect 10459 3621 10468 3655
rect 10416 3612 10468 3621
rect 6920 3340 6972 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 2872 3136 2924 3188
rect 3240 3000 3292 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 6920 3000 6972 3052
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 9956 2796 10008 2848
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 4344 2592 4396 2644
rect 6460 2592 6512 2644
rect 7840 2592 7892 2644
rect 7932 2592 7984 2644
rect 8116 2592 8168 2644
rect 9312 2592 9364 2644
rect 10324 2592 10376 2644
rect 4160 2524 4212 2576
rect 572 2388 624 2440
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4344 2388 4396 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 6920 2320 6972 2372
rect 9956 2388 10008 2440
rect 10048 2320 10100 2372
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 10508 2252 10560 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
<< metal2 >>
rect 754 11200 810 12000
rect 2042 11200 2098 12000
rect 3330 11200 3386 12000
rect 4618 11200 4674 12000
rect 5906 11200 5962 12000
rect 7194 11200 7250 12000
rect 8482 11200 8538 12000
rect 9770 11200 9826 12000
rect 11058 11200 11114 12000
rect 768 9586 796 11200
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1596 9654 1624 10231
rect 2056 9722 2084 11200
rect 3344 10010 3372 11200
rect 3252 9982 3372 10010
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 1584 9648 1636 9654
rect 1214 9616 1270 9625
rect 756 9580 808 9586
rect 1584 9590 1636 9596
rect 1214 9551 1270 9560
rect 1952 9580 2004 9586
rect 756 9522 808 9528
rect 1228 9382 1256 9551
rect 1952 9522 2004 9528
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1216 9376 1268 9382
rect 1216 9318 1268 9324
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8809 980 8842
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 1872 8514 1900 9386
rect 1964 9178 1992 9522
rect 2056 9178 2084 9522
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1872 8486 2084 8514
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1596 7546 1624 8026
rect 1860 7880 1912 7886
rect 1688 7840 1860 7868
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 940 7200 992 7206
rect 938 7168 940 7177
rect 992 7168 994 7177
rect 938 7103 994 7112
rect 1688 6882 1716 7840
rect 1860 7822 1912 7828
rect 1964 7562 1992 8298
rect 2056 7834 2084 8486
rect 2332 8430 2360 8910
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2056 7806 2176 7834
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1596 6866 1716 6882
rect 1780 7534 1992 7562
rect 2056 7546 2084 7686
rect 2044 7540 2096 7546
rect 1596 6860 1728 6866
rect 1596 6854 1676 6860
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6361 980 6666
rect 1596 6390 1624 6854
rect 1676 6802 1728 6808
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1584 6384 1636 6390
rect 938 6352 994 6361
rect 1584 6326 1636 6332
rect 938 6287 994 6296
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 1044 4826 1072 5471
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1032 4820 1084 4826
rect 1032 4762 1084 4768
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1412 4282 1440 4966
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1504 4078 1532 6190
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1688 5386 1716 6666
rect 1596 5358 1716 5386
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1596 4026 1624 5358
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1688 4282 1716 5238
rect 1780 4622 1808 7534
rect 2044 7482 2096 7488
rect 2148 7426 2176 7806
rect 1872 7398 2176 7426
rect 1872 5370 1900 7398
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2516 6798 2544 9386
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2608 6866 2636 7210
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2504 6792 2556 6798
rect 2556 6740 2636 6746
rect 2504 6734 2636 6740
rect 2516 6718 2636 6734
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1596 4010 1716 4026
rect 1596 4004 1728 4010
rect 1596 3998 1676 4004
rect 1676 3946 1728 3952
rect 940 3936 992 3942
rect 938 3904 940 3913
rect 992 3904 994 3913
rect 938 3839 994 3848
rect 1872 3738 1900 5170
rect 1964 4826 1992 6190
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2424 5114 2452 5578
rect 2516 5370 2544 6598
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2424 5086 2544 5114
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4826 2084 4966
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2516 4826 2544 5086
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2608 3534 2636 6718
rect 2700 4010 2728 9658
rect 3252 9654 3280 9982
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 4632 9722 4660 11200
rect 5920 10146 5948 11200
rect 5736 10118 5948 10146
rect 5736 9722 5764 10118
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 7208 9722 7236 11200
rect 8496 10282 8524 11200
rect 8496 10254 8708 10282
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8680 9722 8708 10254
rect 9784 9722 9812 11200
rect 10322 10704 10378 10713
rect 10322 10639 10378 10648
rect 10336 9722 10364 10639
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 10598 9616 10654 9625
rect 10598 9551 10654 9560
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3804 8634 3832 8774
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3896 8498 3924 9318
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 5736 8974 5764 9454
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 4448 8566 4476 8910
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4724 8498 4752 8910
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3988 7834 4016 7890
rect 3896 7806 4016 7834
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 6458 2912 6598
rect 3252 6458 3280 7686
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7002 3648 7346
rect 3896 7342 3924 7806
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7546 4108 7686
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2792 5658 2820 6190
rect 2884 5914 2912 6394
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5914 3188 6054
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3896 5710 3924 7278
rect 4172 6866 4200 7958
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4264 7324 4292 7822
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4344 7336 4396 7342
rect 4264 7296 4344 7324
rect 4344 7278 4396 7284
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4356 6798 4384 7278
rect 4448 7002 4476 7754
rect 4908 7546 4936 7754
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 3988 6186 4016 6734
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5914 4016 6122
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3884 5704 3936 5710
rect 2792 5630 3004 5658
rect 3884 5646 3936 5652
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5352 2820 5510
rect 2792 5324 2912 5352
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2792 4826 2820 5170
rect 2884 4826 2912 5324
rect 2976 4826 3004 5630
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3896 5370 3924 5646
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3896 4622 3924 5306
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2700 3738 2728 3946
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 2884 3194 2912 4558
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 938 3088 994 3097
rect 4172 3058 4200 4082
rect 938 3023 994 3032
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 3252 2650 3280 2994
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 4172 2582 4200 2994
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 4066 2408 4122 2417
rect 584 800 612 2382
rect 1872 1306 1900 2382
rect 3068 1306 3096 2382
rect 4264 2394 4292 6666
rect 4540 6118 4568 7278
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5000 7002 5028 8366
rect 5552 7546 5580 8366
rect 5736 8090 5764 8910
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5828 8090 5856 8502
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 6288 7546 6316 7822
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4632 6458 4660 6870
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 6458 4844 6598
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5184 5914 5212 6190
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 4146 4384 5646
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4448 5370 4476 5578
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4540 4554 4568 5510
rect 5184 5234 5212 5850
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5276 5302 5304 5646
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 5000 4826 5028 5102
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 5184 4282 5212 5170
rect 5368 5166 5396 7414
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5644 5302 5672 7210
rect 6104 6746 6132 7346
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 5736 6718 6132 6746
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 5736 4010 5764 6718
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 6288 5710 6316 6598
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6380 5302 6408 7142
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4622 6316 4966
rect 6472 4690 6500 5170
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6656 4622 6684 9318
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6840 6322 6868 7958
rect 6932 7886 6960 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 8588 8922 8616 9318
rect 8680 9178 8708 9318
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 10414 9072 10470 9081
rect 9036 9036 9088 9042
rect 10414 9007 10416 9016
rect 9036 8978 9088 8984
rect 10468 9007 10470 9016
rect 10416 8978 10468 8984
rect 8588 8894 8708 8922
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8680 8498 8708 8894
rect 9048 8498 9076 8978
rect 10612 8974 10640 9551
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8566 9720 8774
rect 10244 8634 10272 8910
rect 11072 8906 11100 11200
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 7288 8424 7340 8430
rect 7340 8372 7420 8378
rect 7288 8366 7420 8372
rect 7300 8350 7420 8366
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 6866 6960 7346
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 6474 6960 6802
rect 6932 6458 7052 6474
rect 6932 6452 7064 6458
rect 6932 6446 7012 6452
rect 7012 6394 7064 6400
rect 7392 6390 7420 8350
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7546 7788 7686
rect 7852 7546 7880 7822
rect 8588 7818 8616 8230
rect 8680 7886 8708 8434
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 7954 8984 8230
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8680 7410 8708 7686
rect 8772 7546 8800 7822
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7484 7002 7512 7278
rect 9140 7274 9168 8434
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9324 7546 9352 7958
rect 10152 7546 10180 8434
rect 10508 8288 10560 8294
rect 10506 8256 10508 8265
rect 10560 8256 10562 8265
rect 10506 8191 10562 8200
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 7546 10272 7822
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 7576 7002 7604 7210
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6932 5778 6960 6326
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5234 7512 5510
rect 7668 5302 7696 6598
rect 8128 6254 8156 6598
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8680 6254 8708 6598
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5710 8064 6054
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6644 4616 6696 4622
rect 6748 4593 6776 4694
rect 6840 4622 6868 4966
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7576 4758 7604 5102
rect 7760 4826 7788 5102
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 6828 4616 6880 4622
rect 6644 4558 6696 4564
rect 6734 4584 6790 4593
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 6196 4282 6224 4422
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 6380 3942 6408 4558
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2650 4384 2790
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 6472 2650 6500 4150
rect 6656 4078 6684 4558
rect 6828 4558 6880 4564
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6734 4519 6790 4528
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6748 3534 6776 4519
rect 7116 4282 7144 4558
rect 7944 4554 7972 4966
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4282 7236 4422
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7392 3738 7420 4014
rect 7576 3738 7604 4082
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3058 6960 3334
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 4122 2366 4292 2394
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 4066 2343 4122 2352
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 4356 1306 4384 2382
rect 5460 1306 5488 2382
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6656 1306 6684 2382
rect 6932 2378 6960 2994
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7852 2650 7880 4082
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 2650 7972 3470
rect 8128 2650 8156 6190
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8496 4826 8524 5102
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8680 4690 8708 6190
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8864 4146 8892 5510
rect 8956 4622 8984 7210
rect 9324 6866 9352 7482
rect 10428 7449 10456 7686
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10414 7440 10470 7449
rect 9956 7404 10008 7410
rect 10414 7375 10470 7384
rect 9956 7346 10008 7352
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9968 6914 9996 7346
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 9784 6886 9996 6914
rect 10048 6928 10100 6934
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9784 6254 9812 6886
rect 10048 6870 10100 6876
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5914 9260 6054
rect 9324 5914 9352 6122
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5642 9444 6122
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9048 5370 9076 5578
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8944 4616 8996 4622
rect 8942 4584 8944 4593
rect 8996 4584 8998 4593
rect 8942 4519 8998 4528
rect 9048 4282 9076 5102
rect 9140 4282 9168 5578
rect 9876 5370 9904 6326
rect 9968 5914 9996 6734
rect 10060 6458 10088 6870
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9232 4826 9260 5102
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9496 4616 9548 4622
rect 9324 4576 9496 4604
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 9324 2650 9352 4576
rect 9496 4558 9548 4564
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4146 9812 4558
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9876 3942 9904 5102
rect 10152 4826 10180 5170
rect 10244 4826 10272 6258
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4282 10272 4558
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9968 2446 9996 2790
rect 10336 2650 10364 7210
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10414 6352 10470 6361
rect 10414 6287 10470 6296
rect 10428 6186 10456 6287
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10414 5808 10470 5817
rect 10414 5743 10416 5752
rect 10468 5743 10470 5752
rect 10416 5714 10468 5720
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10416 5024 10468 5030
rect 10414 4992 10416 5001
rect 10468 4992 10470 5001
rect 10414 4927 10470 4936
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4185 10456 4422
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10414 4176 10470 4185
rect 10414 4111 10470 4120
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10428 3505 10456 3606
rect 10414 3496 10470 3505
rect 10414 3431 10470 3440
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10416 2848 10468 2854
rect 10468 2796 10548 2802
rect 10416 2790 10548 2796
rect 10428 2774 10548 2790
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10520 2553 10548 2774
rect 10506 2544 10562 2553
rect 10506 2479 10562 2488
rect 7840 2440 7892 2446
rect 9036 2440 9088 2446
rect 7840 2382 7892 2388
rect 8956 2400 9036 2428
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7852 1306 7880 2382
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 1780 1278 1900 1306
rect 2976 1278 3096 1306
rect 4172 1278 4384 1306
rect 5368 1278 5488 1306
rect 6564 1278 6684 1306
rect 7760 1278 7880 1306
rect 1780 800 1808 1278
rect 2976 800 3004 1278
rect 4172 800 4200 1278
rect 5368 800 5396 1278
rect 6564 800 6592 1278
rect 7760 800 7788 1278
rect 8956 800 8984 2400
rect 9036 2382 9088 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9876 1737 9904 2246
rect 9862 1728 9918 1737
rect 9862 1663 9918 1672
rect 10060 1306 10088 2314
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10060 1278 10180 1306
rect 10152 800 10180 1278
rect 10520 921 10548 2246
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 10506 912 10562 921
rect 10506 847 10562 856
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
<< via2 >>
rect 1582 10240 1638 10296
rect 1214 9560 1270 9616
rect 938 8744 994 8800
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 1490 8200 1546 8256
rect 938 7148 940 7168
rect 940 7148 992 7168
rect 992 7148 994 7168
rect 938 7112 994 7148
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 938 6296 994 6352
rect 1030 5480 1086 5536
rect 938 4664 994 4720
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 938 3884 940 3904
rect 940 3884 992 3904
rect 992 3884 994 3904
rect 938 3848 994 3884
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 10322 10648 10378 10704
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10598 9560 10654 9616
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 938 3032 994 3088
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 4066 2352 4122 2408
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10414 9036 10470 9072
rect 10414 9016 10416 9036
rect 10416 9016 10468 9036
rect 10468 9016 10470 9036
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10506 8236 10508 8256
rect 10508 8236 10560 8256
rect 10560 8236 10562 8256
rect 10506 8200 10562 8236
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 6734 4528 6790 4584
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10414 7384 10470 7440
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 8942 4564 8944 4584
rect 8944 4564 8996 4584
rect 8996 4564 8998 4584
rect 8942 4528 8998 4564
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10414 6296 10470 6352
rect 10414 5772 10470 5808
rect 10414 5752 10416 5772
rect 10416 5752 10468 5772
rect 10468 5752 10470 5772
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10414 4972 10416 4992
rect 10416 4972 10468 4992
rect 10468 4972 10470 4992
rect 10414 4936 10470 4972
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10414 4120 10470 4176
rect 10414 3440 10470 3496
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 10506 2488 10562 2544
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 9862 1672 9918 1728
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 10506 856 10562 912
<< metal3 >>
rect 10317 10706 10383 10709
rect 11200 10706 12000 10736
rect 10317 10704 12000 10706
rect 10317 10648 10322 10704
rect 10378 10648 12000 10704
rect 10317 10646 12000 10648
rect 10317 10643 10383 10646
rect 11200 10616 12000 10646
rect 0 10434 800 10464
rect 0 10374 1042 10434
rect 0 10344 800 10374
rect 982 10298 1042 10374
rect 1577 10298 1643 10301
rect 982 10296 1643 10298
rect 982 10240 1582 10296
rect 1638 10240 1643 10296
rect 982 10238 1643 10240
rect 1577 10235 1643 10238
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 11200 9800 12000 9920
rect 10698 9759 11014 9760
rect 11470 9690 11530 9800
rect 0 9618 800 9648
rect 11102 9630 11530 9690
rect 1209 9618 1275 9621
rect 0 9616 1275 9618
rect 0 9560 1214 9616
rect 1270 9560 1275 9616
rect 0 9558 1275 9560
rect 0 9528 800 9558
rect 1209 9555 1275 9558
rect 10593 9618 10659 9621
rect 11102 9618 11162 9630
rect 10593 9616 11162 9618
rect 10593 9560 10598 9616
rect 10654 9560 11162 9616
rect 10593 9558 11162 9560
rect 10593 9555 10659 9558
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 10409 9074 10475 9077
rect 11200 9074 12000 9104
rect 10409 9072 12000 9074
rect 10409 9016 10414 9072
rect 10470 9016 12000 9072
rect 10409 9014 12000 9016
rect 10409 9011 10475 9014
rect 11200 8984 12000 9014
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 1485 8258 1551 8261
rect 798 8256 1551 8258
rect 798 8200 1490 8256
rect 1546 8200 1551 8256
rect 798 8198 1551 8200
rect 798 8016 858 8198
rect 1485 8195 1551 8198
rect 10501 8258 10567 8261
rect 11200 8258 12000 8288
rect 10501 8256 12000 8258
rect 10501 8200 10506 8256
rect 10562 8200 12000 8256
rect 10501 8198 12000 8200
rect 10501 8195 10567 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 11200 8168 12000 8198
rect 9479 8127 9795 8128
rect 0 7926 858 8016
rect 0 7896 800 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 10409 7442 10475 7445
rect 11200 7442 12000 7472
rect 10409 7440 12000 7442
rect 10409 7384 10414 7440
rect 10470 7384 12000 7440
rect 10409 7382 12000 7384
rect 10409 7379 10475 7382
rect 11200 7352 12000 7382
rect 0 7170 800 7200
rect 933 7170 999 7173
rect 0 7168 999 7170
rect 0 7112 938 7168
rect 994 7112 999 7168
rect 0 7110 999 7112
rect 0 7080 800 7110
rect 933 7107 999 7110
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 11200 6536 12000 6656
rect 10698 6495 11014 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 10409 6354 10475 6357
rect 11286 6354 11346 6536
rect 10409 6352 11346 6354
rect 10409 6296 10414 6352
rect 10470 6296 11346 6352
rect 10409 6294 11346 6296
rect 10409 6291 10475 6294
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 10409 5810 10475 5813
rect 11200 5810 12000 5840
rect 10409 5808 12000 5810
rect 10409 5752 10414 5808
rect 10470 5752 12000 5808
rect 10409 5750 12000 5752
rect 10409 5747 10475 5750
rect 11200 5720 12000 5750
rect 0 5538 800 5568
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 0 5478 1091 5480
rect 0 5448 800 5478
rect 1025 5475 1091 5478
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 10409 4994 10475 4997
rect 11200 4994 12000 5024
rect 10409 4992 12000 4994
rect 10409 4936 10414 4992
rect 10470 4936 12000 4992
rect 10409 4934 12000 4936
rect 10409 4931 10475 4934
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 11200 4904 12000 4934
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 6729 4586 6795 4589
rect 8937 4586 9003 4589
rect 6729 4584 9003 4586
rect 6729 4528 6734 4584
rect 6790 4528 8942 4584
rect 8998 4528 9003 4584
rect 6729 4526 9003 4528
rect 6729 4523 6795 4526
rect 8937 4523 9003 4526
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 10409 4178 10475 4181
rect 11200 4178 12000 4208
rect 10409 4176 12000 4178
rect 10409 4120 10414 4176
rect 10470 4120 12000 4176
rect 10409 4118 12000 4120
rect 10409 4115 10475 4118
rect 11200 4088 12000 4118
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 10409 3498 10475 3501
rect 10409 3496 11162 3498
rect 10409 3440 10414 3496
rect 10470 3440 11162 3496
rect 10409 3438 11162 3440
rect 10409 3435 10475 3438
rect 11102 3396 11162 3438
rect 11102 3392 11346 3396
rect 11102 3336 12000 3392
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 11200 3272 12000 3336
rect 10698 3231 11014 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 10501 2546 10567 2549
rect 11200 2546 12000 2576
rect 10501 2544 12000 2546
rect 10501 2488 10506 2544
rect 10562 2488 12000 2544
rect 10501 2486 12000 2488
rect 10501 2483 10567 2486
rect 11200 2456 12000 2486
rect 4061 2410 4127 2413
rect 2454 2408 4127 2410
rect 2454 2352 4066 2408
rect 4122 2352 4127 2408
rect 2454 2350 4127 2352
rect 0 2274 800 2304
rect 2454 2274 2514 2350
rect 4061 2347 4127 2350
rect 0 2214 2514 2274
rect 0 2184 800 2214
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 9857 1730 9923 1733
rect 11200 1730 12000 1760
rect 9857 1728 12000 1730
rect 9857 1672 9862 1728
rect 9918 1672 12000 1728
rect 9857 1670 12000 1672
rect 9857 1667 9923 1670
rect 11200 1640 12000 1670
rect 10501 914 10567 917
rect 11200 914 12000 944
rect 10501 912 12000 914
rect 10501 856 10506 912
rect 10562 856 12000 912
rect 10501 854 12000 856
rect 10501 851 10567 854
rect 11200 824 12000 854
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform -1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform -1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform -1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1688980957
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform -1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform -1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1688980957
transform 1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform -1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform -1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform -1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform -1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1688980957
transform -1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1688980957
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1688980957
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1688980957
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1688980957
transform -1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1688980957
transform -1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1688980957
transform -1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1688980957
transform -1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1688980957
transform -1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1688980957
transform -1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _102_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _103_
timestamp 1688980957
transform 1 0 6532 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _104_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp 1688980957
transform -1 0 3956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _107_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp 1688980957
transform -1 0 5244 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform -1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform -1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1688980957
transform -1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform -1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _131__42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _132_
timestamp 1688980957
transform 1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _133_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10120 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _134_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _135_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _136_
timestamp 1688980957
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _137_
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _138_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _139_
timestamp 1688980957
transform -1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _140_
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _141_
timestamp 1688980957
transform 1 0 9016 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _142_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _143_
timestamp 1688980957
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _144__43
timestamp 1688980957
transform -1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _144_
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _145_
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _146_
timestamp 1688980957
transform -1 0 7636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _147_
timestamp 1688980957
transform 1 0 2208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _148_
timestamp 1688980957
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _149_
timestamp 1688980957
transform -1 0 4416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _150_
timestamp 1688980957
transform -1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _151_
timestamp 1688980957
transform 1 0 3956 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _152_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _153_
timestamp 1688980957
transform -1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _154_
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _155__44
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _155_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _156_
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _157_
timestamp 1688980957
transform 1 0 5060 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _158_
timestamp 1688980957
transform -1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_19
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_23
timestamp 1688980957
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_29
timestamp 1688980957
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_36
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_89
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_95
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_16
timestamp 1688980957
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1688980957
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_98
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_30
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_76
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_88
timestamp 1688980957
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_102
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_12
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_16
timestamp 1688980957
transform 1 0 2576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_23
timestamp 1688980957
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_48
timestamp 1688980957
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1688980957
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_62
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_67
timestamp 1688980957
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_74
timestamp 1688980957
transform 1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_14
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1688980957
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_11
timestamp 1688980957
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_23
timestamp 1688980957
transform 1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_62
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_20
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_24
timestamp 1688980957
transform 1 0 3312 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_40
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_64
timestamp 1688980957
transform 1 0 6992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_42
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_70
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_78
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_91
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 4232 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 8464 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 10212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 1932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1688980957
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1688980957
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1688980957
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal3 s 11200 9800 12000 9920 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 11200 10616 12000 10736 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 3 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 4 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 5 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 6 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 7 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 8 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 9 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 10 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 11 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 12 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 13 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 14 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 15 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 16 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 17 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 18 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 19 nsew signal tristate
flabel metal2 s 754 11200 810 12000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 20 nsew signal input
flabel metal2 s 2042 11200 2098 12000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 21 nsew signal input
flabel metal2 s 3330 11200 3386 12000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 22 nsew signal input
flabel metal2 s 4618 11200 4674 12000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 23 nsew signal input
flabel metal2 s 5906 11200 5962 12000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 24 nsew signal input
flabel metal2 s 7194 11200 7250 12000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 25 nsew signal input
flabel metal2 s 8482 11200 8538 12000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 26 nsew signal input
flabel metal2 s 9770 11200 9826 12000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 27 nsew signal input
flabel metal2 s 11058 11200 11114 12000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 28 nsew signal input
flabel metal3 s 11200 824 12000 944 0 FreeSans 480 0 0 0 chany_top_out[0]
port 29 nsew signal tristate
flabel metal3 s 11200 1640 12000 1760 0 FreeSans 480 0 0 0 chany_top_out[1]
port 30 nsew signal tristate
flabel metal3 s 11200 2456 12000 2576 0 FreeSans 480 0 0 0 chany_top_out[2]
port 31 nsew signal tristate
flabel metal3 s 11200 3272 12000 3392 0 FreeSans 480 0 0 0 chany_top_out[3]
port 32 nsew signal tristate
flabel metal3 s 11200 4088 12000 4208 0 FreeSans 480 0 0 0 chany_top_out[4]
port 33 nsew signal tristate
flabel metal3 s 11200 4904 12000 5024 0 FreeSans 480 0 0 0 chany_top_out[5]
port 34 nsew signal tristate
flabel metal3 s 11200 5720 12000 5840 0 FreeSans 480 0 0 0 chany_top_out[6]
port 35 nsew signal tristate
flabel metal3 s 11200 6536 12000 6656 0 FreeSans 480 0 0 0 chany_top_out[7]
port 36 nsew signal tristate
flabel metal3 s 11200 7352 12000 7472 0 FreeSans 480 0 0 0 chany_top_out[8]
port 37 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
port 38 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 prog_clk
port 39 nsew signal input
flabel metal3 s 11200 8168 12000 8288 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 40 nsew signal tristate
flabel metal3 s 11200 8984 12000 9104 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 41 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 43 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 8280 7378 8280 7378 0 _000_
rlabel metal1 6486 4114 6486 4114 0 _001_
rlabel metal1 9798 5712 9798 5712 0 _002_
rlabel metal1 3312 4590 3312 4590 0 _003_
rlabel metal1 5198 3978 5198 3978 0 _004_
rlabel metal1 2116 4590 2116 4590 0 _005_
rlabel metal1 3634 7820 3634 7820 0 _006_
rlabel metal1 2116 7378 2116 7378 0 _007_
rlabel metal1 3726 8942 3726 8942 0 _008_
rlabel metal1 7544 7378 7544 7378 0 _009_
rlabel metal1 4048 7378 4048 7378 0 _010_
rlabel metal1 8280 4590 8280 4590 0 _011_
rlabel metal1 6210 4590 6210 4590 0 _012_
rlabel metal1 10074 4794 10074 4794 0 _013_
rlabel metal2 9982 6324 9982 6324 0 _014_
rlabel metal2 6578 4420 6578 4420 0 _015_
rlabel metal1 9936 5338 9936 5338 0 _016_
rlabel metal2 7774 4964 7774 4964 0 _017_
rlabel metal1 8556 7514 8556 7514 0 _018_
rlabel metal1 8418 4794 8418 4794 0 _019_
rlabel metal1 7360 3706 7360 3706 0 _020_
rlabel metal1 7314 4522 7314 4522 0 _021_
rlabel metal1 9108 7310 9108 7310 0 _022_
rlabel metal1 9292 4794 9292 4794 0 _023_
rlabel metal1 8832 6766 8832 6766 0 _024_
rlabel metal1 9614 4250 9614 4250 0 _025_
rlabel metal1 3887 9078 3887 9078 0 _026_
rlabel metal1 4186 7480 4186 7480 0 _027_
rlabel metal1 3358 6290 3358 6290 0 _028_
rlabel metal2 7866 7684 7866 7684 0 _029_
rlabel metal1 2530 6834 2530 6834 0 _030_
rlabel metal2 1978 5508 1978 5508 0 _031_
rlabel metal1 4370 8466 4370 8466 0 _032_
rlabel metal1 6164 7514 6164 7514 0 _033_
rlabel metal2 4186 7412 4186 7412 0 _034_
rlabel metal1 7314 6970 7314 6970 0 _035_
rlabel metal1 2484 4794 2484 4794 0 _036_
rlabel metal1 1610 5814 1610 5814 0 _037_
rlabel metal1 6210 5270 6210 5270 0 _038_
rlabel metal2 2990 5219 2990 5219 0 _039_
rlabel metal1 5336 5134 5336 5134 0 _040_
rlabel metal1 2622 5644 2622 5644 0 _041_
rlabel metal1 9890 8976 9890 8976 0 ccff_head
rlabel metal1 10304 9690 10304 9690 0 ccff_tail
rlabel metal2 598 1588 598 1588 0 chany_bottom_in[0]
rlabel metal2 1794 1027 1794 1027 0 chany_bottom_in[1]
rlabel metal2 2990 1027 2990 1027 0 chany_bottom_in[2]
rlabel metal2 4186 1027 4186 1027 0 chany_bottom_in[3]
rlabel metal2 5382 1027 5382 1027 0 chany_bottom_in[4]
rlabel metal2 6578 1027 6578 1027 0 chany_bottom_in[5]
rlabel metal2 7774 1027 7774 1027 0 chany_bottom_in[6]
rlabel metal2 8970 1588 8970 1588 0 chany_bottom_in[7]
rlabel metal2 10166 1027 10166 1027 0 chany_bottom_in[8]
rlabel metal3 820 3060 820 3060 0 chany_bottom_out[0]
rlabel metal3 820 3876 820 3876 0 chany_bottom_out[1]
rlabel metal3 820 4692 820 4692 0 chany_bottom_out[2]
rlabel metal3 866 5508 866 5508 0 chany_bottom_out[3]
rlabel metal3 820 6324 820 6324 0 chany_bottom_out[4]
rlabel metal3 820 7140 820 7140 0 chany_bottom_out[5]
rlabel metal3 751 7956 751 7956 0 chany_bottom_out[6]
rlabel metal3 820 8772 820 8772 0 chany_bottom_out[7]
rlabel metal3 958 9588 958 9588 0 chany_bottom_out[8]
rlabel metal1 782 9520 782 9520 0 chany_top_in[0]
rlabel metal1 2070 9656 2070 9656 0 chany_top_in[1]
rlabel metal1 3450 9554 3450 9554 0 chany_top_in[2]
rlabel metal1 4784 9554 4784 9554 0 chany_top_in[3]
rlabel metal1 5888 9554 5888 9554 0 chany_top_in[4]
rlabel metal1 7360 9554 7360 9554 0 chany_top_in[5]
rlabel metal1 8740 9554 8740 9554 0 chany_top_in[6]
rlabel metal1 9798 9622 9798 9622 0 chany_top_in[7]
rlabel metal1 10166 8908 10166 8908 0 chany_top_in[8]
rlabel metal1 10488 2278 10488 2278 0 chany_top_out[0]
rlabel metal2 9890 1989 9890 1989 0 chany_top_out[1]
rlabel metal3 10910 2516 10910 2516 0 chany_top_out[2]
rlabel metal2 10442 3553 10442 3553 0 chany_top_out[3]
rlabel metal2 10442 4301 10442 4301 0 chany_top_out[4]
rlabel via2 10442 4981 10442 4981 0 chany_top_out[5]
rlabel metal1 10442 5814 10442 5814 0 chany_top_out[6]
rlabel metal2 10442 6239 10442 6239 0 chany_top_out[7]
rlabel metal2 10442 7565 10442 7565 0 chany_top_out[8]
rlabel metal1 5796 5678 5796 5678 0 clknet_0_prog_clk
rlabel metal1 3864 5678 3864 5678 0 clknet_1_0__leaf_prog_clk
rlabel metal1 6578 6324 6578 6324 0 clknet_1_1__leaf_prog_clk
rlabel metal3 843 10404 843 10404 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 6578 5202 6578 5202 0 mem_left_ipin_0.DFF_0_.Q
rlabel metal1 8602 4624 8602 4624 0 mem_left_ipin_0.DFF_1_.Q
rlabel metal1 8096 5542 8096 5542 0 mem_left_ipin_0.DFF_2_.Q
rlabel metal1 3726 4590 3726 4590 0 mem_left_ipin_1.DFF_0_.Q
rlabel metal1 4830 4114 4830 4114 0 mem_left_ipin_1.DFF_1_.Q
rlabel metal1 1794 6834 1794 6834 0 mem_right_ipin_0.DFF_0_.Q
rlabel metal1 4094 7242 4094 7242 0 mem_right_ipin_0.DFF_1_.Q
rlabel metal2 7590 3910 7590 3910 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 4370 3910 4370 3910 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 7038 4250 7038 4250 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal1 7774 4726 7774 4726 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 9706 7310 9706 7310 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal2 8970 8092 8970 8092 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 8418 4250 8418 4250 0 mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 7958 4760 7958 4760 0 mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 9154 7514 9154 7514 0 mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 9016 5338 9016 5338 0 mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9936 6902 9936 6902 0 mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 9982 7139 9982 7139 0 mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 3128 5678 3128 5678 0 mux_left_ipin_1.INVTX1_0_.out
rlabel metal1 1656 6222 1656 6222 0 mux_left_ipin_1.INVTX1_1_.out
rlabel metal1 3174 5848 3174 5848 0 mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5566 5270 5566 5270 0 mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2530 5610 2530 5610 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal1 2162 6834 2162 6834 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal2 7590 7106 7590 7106 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal1 8096 7922 8096 7922 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 3772 5882 3772 5882 0 mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3082 6222 3082 6222 0 mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 6486 7820 6486 7820 0 mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 4830 6902 4830 6902 0 mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5244 8534 5244 8534 0 mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 3772 8602 3772 8602 0 mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 8643 8534 8643 8534 0 net1
rlabel metal1 9982 2618 9982 2618 0 net10
rlabel metal1 2254 4080 2254 4080 0 net11
rlabel metal1 1610 5236 1610 5236 0 net12
rlabel metal2 2576 6732 2576 6732 0 net13
rlabel metal2 3910 8908 3910 8908 0 net14
rlabel metal1 4094 4080 4094 4080 0 net15
rlabel metal2 6946 8602 6946 8602 0 net16
rlabel metal1 8602 7854 8602 7854 0 net17
rlabel metal1 2622 9044 2622 9044 0 net18
rlabel metal1 2346 8364 2346 8364 0 net19
rlabel metal1 1610 2312 1610 2312 0 net2
rlabel metal2 5750 8772 5750 8772 0 net20
rlabel metal1 1794 3400 1794 3400 0 net21
rlabel metal1 1518 4216 1518 4216 0 net22
rlabel metal1 2116 3706 2116 3706 0 net23
rlabel metal2 1886 7548 1886 7548 0 net24
rlabel metal1 2116 3978 2116 3978 0 net25
rlabel metal1 1702 7446 1702 7446 0 net26
rlabel metal1 2967 8534 2967 8534 0 net27
rlabel metal1 2116 8874 2116 8874 0 net28
rlabel metal1 2116 9146 2116 9146 0 net29
rlabel metal2 4186 3570 4186 3570 0 net3
rlabel metal1 10074 2414 10074 2414 0 net30
rlabel metal1 4370 2550 4370 2550 0 net31
rlabel metal1 3933 3162 3933 3162 0 net32
rlabel metal1 10166 3502 10166 3502 0 net33
rlabel metal2 10258 4420 10258 4420 0 net34
rlabel metal1 8970 3910 8970 3910 0 net35
rlabel metal1 10258 5746 10258 5746 0 net36
rlabel metal1 9982 4726 9982 4726 0 net37
rlabel metal2 10258 7684 10258 7684 0 net38
rlabel metal1 2530 8942 2530 8942 0 net39
rlabel metal1 3220 3026 3220 3026 0 net4
rlabel metal1 10120 7514 10120 7514 0 net40
rlabel metal1 10074 8602 10074 8602 0 net41
rlabel metal1 9292 6698 9292 6698 0 net42
rlabel metal1 5336 8398 5336 8398 0 net43
rlabel metal1 6486 5134 6486 5134 0 net44
rlabel metal1 5294 6290 5294 6290 0 net45
rlabel metal1 5903 4522 5903 4522 0 net46
rlabel metal2 4462 5474 4462 5474 0 net47
rlabel metal2 3634 7174 3634 7174 0 net48
rlabel metal1 7815 5678 7815 5678 0 net49
rlabel metal1 6210 2550 6210 2550 0 net5
rlabel metal2 4922 7650 4922 7650 0 net50
rlabel via1 6849 6290 6849 6290 0 net51
rlabel metal1 6072 2618 6072 2618 0 net6
rlabel metal1 7360 2618 7360 2618 0 net7
rlabel metal1 8096 2618 8096 2618 0 net8
rlabel metal1 9292 2618 9292 2618 0 net9
rlabel metal3 1579 2244 1579 2244 0 prog_clk
rlabel metal1 10488 8262 10488 8262 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel metal1 10442 9078 10442 9078 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
