VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.570 -38.270 26.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 -38.270 206.670 326.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 416.820 206.670 640.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 730.820 206.670 954.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 1044.820 206.670 1268.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 1358.820 206.670 1582.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 1672.820 206.670 1896.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 1986.820 206.670 2210.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 2300.820 206.670 2524.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 2614.820 206.670 2838.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 2928.820 206.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 -38.270 386.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 552.965 386.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 866.965 386.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 1180.965 386.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 1494.965 386.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 1808.965 386.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 2122.965 386.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 2436.965 386.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 2750.965 386.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 3064.965 386.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 3378.965 386.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 -38.270 566.670 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 277.980 566.670 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 446.740 566.670 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 589.900 566.670 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 760.740 566.670 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 870.900 566.670 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1074.740 566.670 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1184.900 566.670 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1388.740 566.670 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1498.900 566.670 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1702.740 566.670 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 1812.900 566.670 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2016.740 566.670 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2126.900 566.670 2209.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2330.740 566.670 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2440.900 566.670 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2644.740 566.670 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2754.900 566.670 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 2958.740 566.670 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 3068.900 566.670 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 3250.980 566.670 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 3382.900 566.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 63.900 746.670 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 239.900 746.670 351.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 411.900 746.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 601.660 746.670 665.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 725.900 746.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 915.660 746.670 979.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1039.900 746.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1229.660 746.670 1293.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1353.900 746.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1543.660 746.670 1607.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1667.900 746.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1857.660 746.670 1921.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 1981.900 746.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2171.660 746.670 2235.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2295.900 746.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2485.660 746.670 2549.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2609.900 746.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2799.660 746.670 2857.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 2917.900 746.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 3113.660 746.670 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 3237.900 746.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 3427.660 746.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.570 -38.270 926.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 -38.270 1106.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 552.965 1106.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 866.965 1106.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 1180.965 1106.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 1494.965 1106.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 1808.965 1106.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 2122.965 1106.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 2436.965 1106.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 2750.965 1106.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 3064.965 1106.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 3378.965 1106.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.570 -38.270 1286.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 -38.270 1466.670 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 441.565 1466.670 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 755.565 1466.670 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 1069.565 1466.670 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 1383.565 1466.670 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 1697.565 1466.670 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 2011.565 1466.670 2209.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 2325.565 1466.670 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 2639.565 1466.670 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 2953.565 1466.670 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 3236.285 1466.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 -38.270 1646.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 552.965 1646.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 866.965 1646.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 1180.965 1646.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 1494.965 1646.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 1808.965 1646.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 2122.965 1646.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 2436.965 1646.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 2750.965 1646.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 3064.965 1646.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 3378.965 1646.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 -38.270 1826.670 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 441.565 1826.670 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 589.900 1826.670 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 755.565 1826.670 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 870.900 1826.670 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1069.565 1826.670 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1184.900 1826.670 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1383.565 1826.670 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1498.900 1826.670 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1697.565 1826.670 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 1812.900 1826.670 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2011.565 1826.670 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2126.900 1826.670 2209.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2325.565 1826.670 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2440.900 1826.670 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2639.565 1826.670 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2754.900 1826.670 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 2953.565 1826.670 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 3068.900 1826.670 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 3236.285 1826.670 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 3382.900 1826.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 -38.270 2006.670 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 239.900 2006.670 342.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 411.900 2006.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 601.660 2006.670 656.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 725.900 2006.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 915.660 2006.670 970.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1039.900 2006.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1229.660 2006.670 1284.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1353.900 2006.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1543.660 2006.670 1598.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1667.900 2006.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1857.660 2006.670 1912.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 1981.900 2006.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2171.660 2006.670 2226.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2295.900 2006.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2485.660 2006.670 2540.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2609.900 2006.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2799.660 2006.670 2848.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 2917.900 2006.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 3113.660 2006.670 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 3237.900 2006.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 3499.460 2006.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2183.570 -38.270 2186.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 -38.270 2366.670 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 239.900 2366.670 351.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 411.900 2366.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 601.660 2366.670 665.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 725.900 2366.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 915.660 2366.670 979.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1039.900 2366.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1229.660 2366.670 1293.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1353.900 2366.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1543.660 2366.670 1607.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1667.900 2366.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1857.660 2366.670 1921.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 1981.900 2366.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2171.660 2366.670 2235.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2295.900 2366.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2485.660 2366.670 2549.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2609.900 2366.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2799.660 2366.670 2857.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 2917.900 2366.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 3113.660 2366.670 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 3237.900 2366.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 3427.660 2366.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2543.570 -38.270 2546.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 -38.270 2726.670 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 552.965 2726.670 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 866.965 2726.670 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 1180.965 2726.670 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 1494.965 2726.670 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 1808.965 2726.670 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 2122.965 2726.670 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 2436.965 2726.670 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 2750.965 2726.670 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 3064.965 2726.670 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.570 3378.965 2726.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2903.570 -38.270 2906.670 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 16.530 2963.250 19.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 46.530 2963.250 49.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 76.530 2963.250 79.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 106.530 2963.250 109.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 136.530 2963.250 139.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 166.530 2963.250 169.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 196.530 2963.250 199.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 226.530 2963.250 229.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 256.530 2963.250 259.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 286.530 2963.250 289.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 316.530 2963.250 319.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 346.530 2963.250 349.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 376.530 2963.250 379.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 406.530 2963.250 409.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 436.530 2963.250 439.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 466.530 2963.250 469.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 496.530 2963.250 499.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 526.530 2963.250 529.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 556.530 2963.250 559.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 586.530 2963.250 589.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 616.530 2963.250 619.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 646.530 2963.250 649.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 676.530 2963.250 679.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 706.530 2963.250 709.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 736.530 2963.250 739.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 766.530 2963.250 769.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 796.530 2963.250 799.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 826.530 2963.250 829.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 856.530 2963.250 859.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 886.530 2963.250 889.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 916.530 2963.250 919.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 946.530 2963.250 949.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 976.530 2963.250 979.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1006.530 2963.250 1009.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1036.530 2963.250 1039.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1066.530 2963.250 1069.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1096.530 2963.250 1099.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1126.530 2963.250 1129.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1156.530 2963.250 1159.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1186.530 2963.250 1189.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1216.530 2963.250 1219.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1246.530 2963.250 1249.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1276.530 2963.250 1279.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1306.530 2963.250 1309.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1336.530 2963.250 1339.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1366.530 2963.250 1369.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1396.530 2963.250 1399.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1426.530 2963.250 1429.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1456.530 2963.250 1459.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1486.530 2963.250 1489.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1516.530 2963.250 1519.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1546.530 2963.250 1549.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1576.530 2963.250 1579.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1606.530 2963.250 1609.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1636.530 2963.250 1639.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1666.530 2963.250 1669.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1696.530 2963.250 1699.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1726.530 2963.250 1729.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1756.530 2963.250 1759.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1786.530 2963.250 1789.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1816.530 2963.250 1819.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1846.530 2963.250 1849.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1876.530 2963.250 1879.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1906.530 2963.250 1909.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1936.530 2963.250 1939.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1966.530 2963.250 1969.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1996.530 2963.250 1999.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2026.530 2963.250 2029.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2056.530 2963.250 2059.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2086.530 2963.250 2089.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2116.530 2963.250 2119.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2146.530 2963.250 2149.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2176.530 2963.250 2179.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2206.530 2963.250 2209.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2236.530 2963.250 2239.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2266.530 2963.250 2269.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2296.530 2963.250 2299.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2326.530 2963.250 2329.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2356.530 2963.250 2359.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2386.530 2963.250 2389.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2416.530 2963.250 2419.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2446.530 2963.250 2449.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2476.530 2963.250 2479.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2506.530 2963.250 2509.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2536.530 2963.250 2539.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2566.530 2963.250 2569.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2596.530 2963.250 2599.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2626.530 2963.250 2629.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2656.530 2963.250 2659.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2686.530 2963.250 2689.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2716.530 2963.250 2719.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2746.530 2963.250 2749.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2776.530 2963.250 2779.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2806.530 2963.250 2809.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2836.530 2963.250 2839.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2866.530 2963.250 2869.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2896.530 2963.250 2899.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2926.530 2963.250 2929.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2956.530 2963.250 2959.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2986.530 2963.250 2989.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3016.530 2963.250 3019.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3046.530 2963.250 3049.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3076.530 2963.250 3079.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3106.530 2963.250 3109.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3136.530 2963.250 3139.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3166.530 2963.250 3169.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3196.530 2963.250 3199.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3226.530 2963.250 3229.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3256.530 2963.250 3259.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3286.530 2963.250 3289.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3316.530 2963.250 3319.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3346.530 2963.250 3349.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3376.530 2963.250 3379.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3406.530 2963.250 3409.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3436.530 2963.250 3439.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3466.530 2963.250 3469.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3496.530 2963.250 3499.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 516.560 109.650 536.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 165.680 469.370 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 611.630 1079.600 614.730 1090.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 337.040 789.530 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.510 976.240 1110.610 1042.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 655.280 1439.050 737.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 595.440 1574.290 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 1280.880 1750.010 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.350 2678.960 1894.450 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 1593.680 2070.170 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.510 3073.360 2214.610 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 1906.480 2389.410 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 1378.800 2832.850 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 796.720 109.650 851.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 326.160 469.370 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 611.630 875.600 614.730 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 165.680 789.530 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.510 1917.360 1110.610 1983.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 965.360 1439.050 1052.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1079.600 1574.290 1118.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 652.560 1750.010 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.350 3073.360 1894.450 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 1280.880 2070.170 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.510 3307.280 2214.610 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 1593.680 2389.410 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2810.430 1694.320 2813.530 1746.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 1109.520 109.650 1164.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 652.560 469.370 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 611.630 3073.360 614.730 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 965.360 789.530 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.510 176.560 1110.610 242.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 339.760 1439.050 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 454.000 1574.290 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 1593.680 1750.010 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.350 875.600 1894.450 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 1906.480 2070.170 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 796.720 2215.530 875.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 1280.880 2389.410 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 2007.120 2832.850 2062.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 1425.040 109.650 1477.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 965.360 469.370 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 516.560 615.650 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 652.560 789.530 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.510 3174.000 1110.610 3239.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 165.680 1439.050 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 766.800 1574.290 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 337.040 1750.010 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.350 1079.600 1894.450 1090.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 2222.000 2070.170 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2188.510 875.600 2191.610 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 2534.800 2389.410 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2810.430 2322.640 2813.530 2374.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 1737.840 109.650 1792.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 1280.880 469.370 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 796.720 615.650 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 1593.680 789.530 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 1906.480 1439.050 1994.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1191.120 1574.290 1243.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 965.360 1750.010 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.350 3307.280 1894.450 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 337.040 2070.170 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 1425.040 2215.530 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 652.560 2389.410 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 437.680 2832.850 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 2053.360 109.650 2105.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 1593.680 469.370 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 1109.520 615.650 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 1289.520 789.530 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 2222.000 1439.050 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 875.600 1574.290 930.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 1906.480 1750.010 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 516.560 1895.370 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 652.560 2070.170 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 2366.160 2215.530 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 337.040 2389.410 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 750.480 2832.850 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 2366.160 109.650 2421.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 1906.480 469.370 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 1425.040 615.650 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 2222.000 789.530 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 1280.880 1439.050 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1707.920 1574.290 1746.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 2534.800 1750.010 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 796.720 1895.370 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 965.360 2070.170 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 516.560 2215.530 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 2844.880 2389.410 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2810.430 1066.000 2813.530 1118.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 2681.680 109.650 2733.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 2222.000 469.370 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 1737.840 615.650 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 1906.480 789.530 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 1596.400 1439.050 1678.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1395.120 1574.290 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 165.680 1750.010 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 1109.520 1895.370 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 2534.800 2070.170 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 2053.360 2215.530 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 965.360 2389.410 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 2950.960 2832.850 3003.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 2994.480 109.650 3049.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 2534.800 469.370 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 2053.360 615.650 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 2853.520 789.530 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 3163.120 1439.050 3250.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1503.920 1574.290 1558.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 2222.000 1750.010 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 1737.840 1895.370 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 165.680 2070.170 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 1109.520 2215.530 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 2635.440 2832.850 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 106.550 3310.000 109.650 3362.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 2844.880 469.370 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 2366.160 615.650 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 2534.800 789.530 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 1819.440 1574.290 1871.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 3163.120 1750.010 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 1425.040 1895.370 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 2681.680 2215.530 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 165.680 2389.410 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 525.600 2835.610 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.590 981.680 304.690 1042.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 466.270 3163.120 469.370 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 2681.680 615.650 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 2537.520 1439.050 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2023.440 1574.290 2062.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.910 2844.880 1750.010 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 2366.160 1895.370 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 2994.480 2215.530 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 2222.000 2389.410 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 3263.760 2832.850 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.590 1922.800 304.690 1983.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 2994.480 615.650 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.430 3163.120 789.530 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.950 2847.600 1439.050 2929.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2132.240 1574.290 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 2690.720 1895.370 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 3319.040 2215.530 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 805.760 2835.610 859.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.950 182.000 335.050 242.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.550 3310.000 615.650 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2336.240 1574.290 2374.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 2994.480 1895.370 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 2853.520 2070.170 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.430 1737.840 2215.530 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.310 3163.120 2389.410 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2837.110 1112.240 2840.210 1175.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 165.680 639.570 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.390 2447.760 1537.490 2499.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 3319.040 1895.370 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2067.070 3163.120 2070.170 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 337.040 2239.450 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 1434.080 2835.610 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 337.040 639.570 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2651.760 1574.290 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 165.680 1920.210 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 437.680 2217.370 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2837.110 1737.840 2840.210 1803.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 437.680 617.490 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2760.560 1574.290 2815.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.270 2053.360 1895.370 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 165.680 2239.450 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 2690.720 2835.610 2744.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 652.560 639.570 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 2964.560 1574.290 3003.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 337.040 1920.210 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 750.480 2217.370 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 2062.400 2835.610 2116.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 750.480 617.490 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 3073.360 1574.290 3128.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 437.680 1897.210 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 652.560 2239.450 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 3003.520 2835.610 3057.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 965.360 639.570 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 3263.760 1574.290 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 652.560 1920.210 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 1066.000 2217.370 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2837.110 2368.880 2840.210 2429.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 1066.000 617.490 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.190 3388.880 1574.290 3441.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 750.480 1897.210 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 965.360 2239.450 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2832.510 3319.040 2835.610 3373.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.630 1278.160 637.730 1289.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 525.600 1576.130 595.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 965.360 1920.210 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 1378.800 2217.370 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 1289.920 639.570 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 805.760 1576.130 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 1066.000 1897.210 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 1593.680 2239.450 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 1378.800 617.490 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 793.790 1280.880 796.890 1294.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 1118.560 1576.130 1190.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 1593.680 1920.210 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.910 1672.560 2210.010 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 1593.680 639.570 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 1434.080 1576.130 1503.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 1280.880 1920.210 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 1694.320 2217.370 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 607.030 1672.560 610.130 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 1746.880 1576.130 1819.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 1378.800 1897.210 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 1280.880 2239.450 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 1694.320 617.490 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 793.790 1667.120 796.890 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 2062.400 1576.130 2131.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 1906.480 1920.210 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 2007.120 2217.370 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 1906.480 639.570 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 2375.200 1576.130 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1886.750 1672.560 1889.850 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 2222.000 2239.450 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 2007.120 617.490 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 2690.720 1576.130 2760.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 1694.320 1897.210 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.430 1667.120 2077.530 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 1906.480 2239.450 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 2222.000 639.570 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 3003.520 1576.130 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 2007.120 1897.210 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 2322.640 2217.370 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.590 1667.120 2397.690 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 2322.640 617.490 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.030 3319.040 1576.130 3388.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 2222.000 1920.210 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 2534.800 2239.450 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 2534.800 639.570 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 437.680 1577.050 453.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 2322.640 1897.210 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 2635.440 2217.370 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 2635.440 617.490 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 750.480 1577.050 766.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 2534.800 1920.210 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 2844.880 2239.450 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.630 2842.160 637.730 2853.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 1066.000 1577.050 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 2635.440 1897.210 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.270 2950.960 2217.370 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 2853.920 639.570 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 1378.800 1577.050 1394.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.110 2950.960 1897.210 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.350 3163.120 2239.450 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.630 2948.240 637.730 2959.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 1694.320 1577.050 1707.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1914.350 2842.160 1917.450 2853.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.390 2956.400 617.490 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 793.790 2844.880 796.890 2858.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 2007.120 1577.050 2023.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 3163.120 1920.210 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.470 3163.120 639.570 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 2322.640 1577.050 2335.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.110 2853.920 1920.210 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 2635.440 1577.050 2651.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.430 2844.880 2077.530 2858.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1573.950 2950.960 1577.050 2964.160 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.970 -38.270 8.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 -38.270 188.070 326.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 416.820 188.070 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 589.900 188.070 640.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 730.820 188.070 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 870.900 188.070 954.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1044.820 188.070 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1184.900 188.070 1268.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1358.820 188.070 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1498.900 188.070 1582.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1672.820 188.070 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1812.900 188.070 1896.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 1986.820 188.070 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2126.900 188.070 2210.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2300.820 188.070 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2440.900 188.070 2524.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2614.820 188.070 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2754.900 188.070 2838.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 2928.820 188.070 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 3068.900 188.070 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.970 3382.900 188.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 -38.270 368.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 552.965 368.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 866.965 368.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 1180.965 368.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 1494.965 368.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 1808.965 368.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 2122.965 368.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 2436.965 368.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 2750.965 368.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 3064.965 368.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.970 3378.965 368.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 -38.270 548.070 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 277.980 548.070 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 446.740 548.070 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 589.900 548.070 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 760.740 548.070 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 870.900 548.070 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1074.740 548.070 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1184.900 548.070 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1388.740 548.070 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1498.900 548.070 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1702.740 548.070 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 1812.900 548.070 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2016.740 548.070 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2126.900 548.070 2209.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2330.740 548.070 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2440.900 548.070 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2644.740 548.070 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2754.900 548.070 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 2958.740 548.070 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 3068.900 548.070 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 3250.980 548.070 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.970 3382.900 548.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 -38.270 728.070 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 239.900 728.070 342.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 411.900 728.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 601.660 728.070 656.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 725.900 728.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 915.660 728.070 970.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1039.900 728.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1229.660 728.070 1284.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1353.900 728.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1543.660 728.070 1598.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1667.900 728.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1857.660 728.070 1912.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 1981.900 728.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2171.660 728.070 2226.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2295.900 728.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2485.660 728.070 2540.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2609.900 728.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2799.660 728.070 2848.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 2917.900 728.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 3113.660 728.070 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.970 3237.900 728.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.970 -38.270 908.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 -38.270 1088.070 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 239.900 1088.070 351.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 411.900 1088.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 552.965 1088.070 665.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 725.900 1088.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 866.965 1088.070 979.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1039.900 1088.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1180.965 1088.070 1293.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1353.900 1088.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1494.965 1088.070 1607.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1667.900 1088.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1808.965 1088.070 1921.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 1981.900 1088.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2122.965 1088.070 2235.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2295.900 1088.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2436.965 1088.070 2549.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2609.900 1088.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2750.965 1088.070 2857.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 2917.900 1088.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 3064.965 1088.070 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 3237.900 1088.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.970 3378.965 1088.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.970 -38.270 1268.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 -38.270 1448.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 552.965 1448.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 866.965 1448.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 1180.965 1448.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 1494.965 1448.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 1808.965 1448.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 2122.965 1448.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 2436.965 1448.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 2750.965 1448.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 3064.965 1448.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.970 3378.965 1448.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.970 -38.270 1628.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 -38.270 1808.070 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 441.565 1808.070 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 589.900 1808.070 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 755.565 1808.070 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 870.900 1808.070 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1069.565 1808.070 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1184.900 1808.070 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1383.565 1808.070 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1498.900 1808.070 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1697.565 1808.070 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 1812.900 1808.070 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2011.565 1808.070 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2126.900 1808.070 2209.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2325.565 1808.070 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2440.900 1808.070 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2639.565 1808.070 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2754.900 1808.070 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 2953.565 1808.070 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 3068.900 1808.070 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 3236.285 1808.070 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.970 3382.900 1808.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 -38.270 1988.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 552.965 1988.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 866.965 1988.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 1180.965 1988.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 1494.965 1988.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 1808.965 1988.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 2122.965 1988.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 2436.965 1988.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 2750.965 1988.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 3064.965 1988.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.970 3378.965 1988.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 -38.270 2168.070 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 277.980 2168.070 325.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 446.740 2168.070 529.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 589.900 2168.070 639.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 760.740 2168.070 810.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 870.900 2168.070 953.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1074.740 2168.070 1124.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1184.900 2168.070 1267.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1388.740 2168.070 1438.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1498.900 2168.070 1581.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1702.740 2168.070 1752.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 1812.900 2168.070 1895.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2016.740 2168.070 2066.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2126.900 2168.070 2209.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2330.740 2168.070 2380.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2440.900 2168.070 2523.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2644.740 2168.070 2694.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2754.900 2168.070 2837.315 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 2958.740 2168.070 3008.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 3068.900 2168.070 3145.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 3250.980 2168.070 3322.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.970 3382.900 2168.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 63.900 2348.070 179.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 239.900 2348.070 351.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 411.900 2348.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 601.660 2348.070 665.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 725.900 2348.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 915.660 2348.070 979.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1039.900 2348.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1229.660 2348.070 1293.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1353.900 2348.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1543.660 2348.070 1607.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1667.900 2348.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1857.660 2348.070 1921.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 1981.900 2348.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2171.660 2348.070 2235.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2295.900 2348.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2485.660 2348.070 2549.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2609.900 2348.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2799.660 2348.070 2857.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 2917.900 2348.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 3113.660 2348.070 3177.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 3237.900 2348.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.970 3427.660 2348.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2524.970 -38.270 2528.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 -38.270 2708.070 450.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 552.965 2708.070 764.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 866.965 2708.070 1078.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 1180.965 2708.070 1392.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 1494.965 2708.070 1706.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 1808.965 2708.070 2020.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 2122.965 2708.070 2334.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 2436.965 2708.070 2648.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 2750.965 2708.070 2962.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 3064.965 2708.070 3276.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.970 3378.965 2708.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2884.970 -38.270 2888.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 10.330 2963.250 13.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 40.330 2963.250 43.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.330 2963.250 73.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 100.330 2963.250 103.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 130.330 2963.250 133.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.330 2963.250 163.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 190.330 2963.250 193.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 220.330 2963.250 223.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.330 2963.250 253.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 280.330 2963.250 283.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 310.330 2963.250 313.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.330 2963.250 343.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 370.330 2963.250 373.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 400.330 2963.250 403.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.330 2963.250 433.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 460.330 2963.250 463.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 490.330 2963.250 493.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.330 2963.250 523.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 550.330 2963.250 553.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 580.330 2963.250 583.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.330 2963.250 613.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 640.330 2963.250 643.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 670.330 2963.250 673.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.330 2963.250 703.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 730.330 2963.250 733.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 760.330 2963.250 763.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.330 2963.250 793.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 820.330 2963.250 823.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 850.330 2963.250 853.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.330 2963.250 883.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 910.330 2963.250 913.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 940.330 2963.250 943.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.330 2963.250 973.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1000.330 2963.250 1003.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1030.330 2963.250 1033.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.330 2963.250 1063.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1090.330 2963.250 1093.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1120.330 2963.250 1123.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.330 2963.250 1153.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1180.330 2963.250 1183.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1210.330 2963.250 1213.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.330 2963.250 1243.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1270.330 2963.250 1273.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1300.330 2963.250 1303.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.330 2963.250 1333.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1360.330 2963.250 1363.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1390.330 2963.250 1393.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.330 2963.250 1423.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1450.330 2963.250 1453.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1480.330 2963.250 1483.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.330 2963.250 1513.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1540.330 2963.250 1543.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1570.330 2963.250 1573.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.330 2963.250 1603.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1630.330 2963.250 1633.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1660.330 2963.250 1663.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.330 2963.250 1693.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1720.330 2963.250 1723.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1750.330 2963.250 1753.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.330 2963.250 1783.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1810.330 2963.250 1813.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1840.330 2963.250 1843.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.330 2963.250 1873.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1900.330 2963.250 1903.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1930.330 2963.250 1933.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.330 2963.250 1963.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1990.330 2963.250 1993.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2020.330 2963.250 2023.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.330 2963.250 2053.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2080.330 2963.250 2083.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2110.330 2963.250 2113.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.330 2963.250 2143.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2170.330 2963.250 2173.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2200.330 2963.250 2203.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.330 2963.250 2233.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2260.330 2963.250 2263.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2290.330 2963.250 2293.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.330 2963.250 2323.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2350.330 2963.250 2353.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2380.330 2963.250 2383.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.330 2963.250 2413.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2440.330 2963.250 2443.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2470.330 2963.250 2473.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.330 2963.250 2503.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2530.330 2963.250 2533.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2560.330 2963.250 2563.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.330 2963.250 2593.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2620.330 2963.250 2623.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2650.330 2963.250 2653.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.330 2963.250 2683.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2710.330 2963.250 2713.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2740.330 2963.250 2743.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.330 2963.250 2773.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2800.330 2963.250 2803.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2830.330 2963.250 2833.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.330 2963.250 2863.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2890.330 2963.250 2893.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2920.330 2963.250 2923.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.330 2963.250 2953.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2980.330 2963.250 2983.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3010.330 2963.250 3013.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.330 2963.250 3043.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3070.330 2963.250 3073.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3100.330 2963.250 3103.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.330 2963.250 3133.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3160.330 2963.250 3163.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3190.330 2963.250 3193.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.330 2963.250 3223.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3250.330 2963.250 3253.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3280.330 2963.250 3283.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.330 2963.250 3313.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3340.330 2963.250 3343.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3370.330 2963.250 3373.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.330 2963.250 3403.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3430.330 2963.250 3433.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3460.330 2963.250 3463.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.330 2963.250 3493.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 516.560 113.330 536.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 799.440 271.570 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 165.680 488.690 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.950 1079.600 634.050 1090.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 337.040 808.850 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 549.200 945.010 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.830 976.240 1129.930 1042.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 595.440 1593.610 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 1280.880 1769.330 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1910.670 2678.960 1913.770 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 1593.680 2089.490 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2230.830 3073.360 2233.930 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 1906.480 2408.730 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2715.670 2545.680 2718.770 2611.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 1378.800 2836.530 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 1697.040 2901.850 1800.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 796.720 113.330 851.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 516.560 271.570 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 326.160 488.690 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.950 875.600 634.050 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 165.680 808.850 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1131.280 945.010 1180.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.830 1917.360 1129.930 1983.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1079.600 1593.610 1118.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 652.560 1769.330 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1910.670 3073.360 1913.770 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 1280.880 2089.490 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2230.830 3307.280 2233.930 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 1593.680 2408.730 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 1694.320 2832.850 1746.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 1381.520 2901.850 1485.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 1109.520 113.330 1164.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 1425.040 271.570 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 652.560 488.690 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.950 3073.360 634.050 3084.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 965.360 808.850 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 532.880 945.010 544.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.830 176.560 1129.930 242.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 454.000 1593.610 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 1593.680 1769.330 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1910.670 875.600 1913.770 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 1906.480 2089.490 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 796.720 2234.850 875.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 1280.880 2408.730 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 2007.120 2836.530 2062.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 2322.640 2901.850 2426.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 1425.040 113.330 1477.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 1109.520 271.570 1197.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 965.360 488.690 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 516.560 634.970 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 652.560 808.850 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 810.320 945.010 870.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.830 3174.000 1129.930 3239.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 766.800 1593.610 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 337.040 1769.330 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1910.670 1079.600 1913.770 1090.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 2222.000 2089.490 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2207.830 875.600 2210.930 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 2534.800 2408.730 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2715.670 1604.560 2718.770 1670.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 2322.640 2832.850 2374.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 2007.120 2901.850 2116.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 1737.840 113.330 1792.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 2056.080 271.570 2138.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 1280.880 488.690 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 796.720 634.970 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 1593.680 808.850 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 565.520 945.010 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 168.400 1118.890 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1191.120 1593.610 1243.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 965.360 1769.330 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1910.670 3307.280 1913.770 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 337.040 2089.490 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 1425.040 2234.850 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 652.560 2408.730 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 437.680 2836.530 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 1066.000 2901.850 1175.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 2053.360 113.330 2105.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 1740.560 271.570 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 1593.680 488.690 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 1109.520 634.970 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 1289.520 808.850 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1441.360 945.010 1452.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 190.160 1118.890 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 875.600 1593.610 930.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 1906.480 1769.330 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 516.560 1914.690 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 652.560 2089.490 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 2366.160 2234.850 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 337.040 2408.730 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 750.480 2836.530 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 2638.160 2901.850 2742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 2366.160 113.330 2421.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 2681.680 271.570 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 1906.480 488.690 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 1425.040 634.970 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 2222.000 808.850 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1751.440 945.010 1762.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 217.360 1118.890 234.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1707.920 1593.610 1746.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 2534.800 1769.330 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 796.720 1914.690 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 965.360 2089.490 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 516.560 2234.850 604.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 2844.880 2408.730 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2715.670 347.920 2718.770 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.750 1066.000 2832.850 1118.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 2953.680 2901.850 3057.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 2681.680 113.330 2733.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 2366.160 271.570 2453.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 2222.000 488.690 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 1737.840 634.970 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 1906.480 808.850 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1457.680 945.010 1469.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 337.040 1118.890 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1395.120 1593.610 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 165.680 1769.330 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 1109.520 1914.690 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 2534.800 2089.490 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 2053.360 2234.850 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 965.360 2408.730 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 2950.960 2836.530 3003.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 440.400 2901.850 544.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 2994.480 113.330 3049.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 3312.720 271.570 3394.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 2534.800 488.690 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 2053.360 634.970 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 2853.520 808.850 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1474.000 945.010 1485.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 652.560 1118.890 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1503.920 1593.610 1558.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 2222.000 1769.330 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 1737.840 1914.690 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 165.680 2089.490 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 1109.520 2234.850 1199.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 2635.440 2836.530 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 750.480 2901.850 859.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 3310.000 113.330 3362.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.470 2997.200 271.570 3079.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 2844.880 488.690 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 2366.160 634.970 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 2534.800 808.850 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1767.760 945.010 1779.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 968.080 1118.890 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 1819.440 1593.610 1871.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 3163.120 1769.330 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 1425.040 1914.690 1512.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 2681.680 2234.850 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 165.680 2408.730 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 525.600 2839.290 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.590 3163.120 488.690 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 2681.680 634.970 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1784.080 945.010 1795.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 1289.520 1118.890 1365.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2023.440 1593.610 2062.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.230 2844.880 1769.330 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 2366.160 1914.690 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 2994.480 2234.850 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 2222.000 2408.730 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.430 3263.760 2836.530 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 2994.480 634.970 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.750 3163.120 808.850 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 1800.400 945.010 1811.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 1593.680 1118.890 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2132.240 1593.610 2187.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 2690.720 1914.690 2769.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 3319.040 2234.850 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 805.760 2839.290 859.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.870 3310.000 634.970 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2077.840 945.010 2089.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 1909.200 1118.890 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2336.240 1593.610 2374.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 2994.480 1914.690 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 2853.520 2089.490 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.750 1737.840 2234.850 1828.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2405.630 3163.120 2408.730 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.790 1112.240 2843.890 1175.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 165.680 658.890 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2094.160 945.010 2105.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 2224.720 1118.890 2306.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.710 2447.760 1556.810 2499.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 3319.040 1914.690 3397.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.390 3163.120 2089.490 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 337.040 2258.770 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 1434.080 2839.290 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 337.040 658.890 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2110.480 945.010 2121.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 2534.800 1118.890 2622.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2651.760 1593.610 2690.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 165.680 1939.530 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 437.680 2236.690 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.790 1737.840 2843.890 1803.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2898.750 3263.760 2901.850 3373.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 437.680 636.810 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2387.920 945.010 2399.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 2844.880 1118.890 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2760.560 1593.610 2815.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.590 2053.360 1914.690 2140.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 165.680 2258.770 253.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 2690.720 2839.290 2744.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 652.560 658.890 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2404.240 945.010 2415.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 3165.840 1118.890 3182.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 2964.560 1593.610 3003.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 337.040 1939.530 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 750.480 2236.690 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 2062.400 2839.290 2116.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 750.480 636.810 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2420.560 945.010 2431.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 3187.600 1118.890 3198.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 3073.360 1593.610 3128.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 437.680 1916.530 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 652.560 2258.770 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 3003.520 2839.290 3057.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 965.360 658.890 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2698.000 945.010 2709.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 3203.920 1118.890 3215.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 3263.760 1593.610 3318.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 652.560 1939.530 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 1066.000 2236.690 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.790 2368.880 2843.890 2429.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 1066.000 636.810 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2714.320 945.010 2725.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 3220.240 1118.890 3231.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.510 3388.880 1593.610 3441.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 750.480 1916.530 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 965.360 2258.770 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.190 3319.040 2839.290 3373.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.950 1278.160 657.050 1289.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 2730.640 945.010 2742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 3236.560 1118.890 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 525.600 1595.450 595.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 965.360 1939.530 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 1378.800 2236.690 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 1289.920 658.890 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3008.080 945.010 3019.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 805.760 1595.450 875.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 1066.000 1916.530 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 1593.680 2258.770 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 1378.800 636.810 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.470 1280.880 800.570 1294.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3024.400 945.010 3035.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 1118.560 1595.450 1190.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 1593.680 1939.530 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2226.230 1672.560 2229.330 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 1593.680 658.890 1672.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3040.720 945.010 3052.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 1434.080 1595.450 1503.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 1280.880 1939.530 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 1694.320 2236.690 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 626.350 1672.560 629.450 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3057.040 945.010 3068.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 1746.880 1595.450 1819.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 1378.800 1916.530 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 1280.880 2258.770 1368.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 1694.320 636.810 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.470 1667.120 800.570 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3334.480 945.010 3345.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 2062.400 1595.450 2131.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 1906.480 1939.530 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 2007.120 2236.690 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 1906.480 658.890 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3350.800 945.010 3362.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 2375.200 1595.450 2456.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1906.070 1672.560 1909.170 1683.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 2222.000 2258.770 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 2007.120 636.810 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.910 3367.120 945.010 3378.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 2690.720 1595.450 2760.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 1694.320 1916.530 1716.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.110 1667.120 2081.210 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 1906.480 2258.770 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 2222.000 658.890 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 168.400 968.930 244.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 3003.520 1595.450 3072.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 2007.120 1916.530 2032.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 2322.640 2236.690 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2398.270 1667.120 2401.370 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 2322.640 636.810 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1018.270 244.560 1021.370 255.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1592.350 3319.040 1595.450 3388.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 2222.000 1939.530 2309.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 2534.800 2258.770 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 2534.800 658.890 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 337.040 968.930 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.790 239.120 1118.890 250.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 437.680 1596.370 453.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 2322.640 1916.530 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 2635.440 2236.690 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 2635.440 636.810 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 440.400 946.850 462.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 750.480 1596.370 766.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 2534.800 1939.530 2625.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 2844.880 2258.770 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.950 2842.160 657.050 2853.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 652.560 968.930 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 1066.000 1596.370 1079.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 2635.440 1916.530 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2233.590 2950.960 2236.690 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 2853.920 658.890 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 750.480 946.850 772.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 1378.800 1596.370 1394.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.430 2950.960 1916.530 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.670 3163.120 2258.770 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.950 2948.240 657.050 2959.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 968.080 968.930 1055.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 1694.320 1596.370 1707.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.670 2842.160 1936.770 2853.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 633.710 2960.000 636.810 2973.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.470 2844.880 800.570 2858.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 1066.000 946.850 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 2007.120 1596.370 2023.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 3163.120 1939.530 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.790 3163.120 658.890 3253.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1018.270 1278.160 1021.370 1289.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 2322.640 1596.370 2335.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.430 2853.920 1939.530 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 1289.040 968.930 1365.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 2635.440 1596.370 2651.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.110 2844.880 2081.210 2858.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 1381.520 946.850 1403.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1110.270 1283.600 1113.370 1294.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.270 2950.960 1596.370 2964.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 1593.680 968.930 1681.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 1697.040 946.850 1713.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 1909.200 968.930 1996.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 2007.120 946.850 2029.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 2224.720 968.930 2306.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 2322.640 946.850 2344.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 2534.800 968.930 2622.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 2638.160 946.850 2660.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 2844.880 968.930 2932.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 943.750 2953.680 946.850 2970.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 965.830 3165.840 968.930 3253.360 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 3.750 10.640 2917.250 3509.040 ;
      LAYER met2 ;
        RECT 3.770 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.220 3518.050 ;
        RECT 3.770 2.680 2917.220 3517.320 ;
        RECT 3.770 1.630 7.950 2.680 ;
        RECT 9.070 1.630 13.930 2.680 ;
        RECT 15.050 1.630 19.910 2.680 ;
        RECT 21.030 1.630 25.890 2.680 ;
        RECT 27.010 1.630 31.870 2.680 ;
        RECT 32.990 1.630 37.850 2.680 ;
        RECT 38.970 1.630 43.370 2.680 ;
        RECT 44.490 1.630 49.350 2.680 ;
        RECT 50.470 1.630 55.330 2.680 ;
        RECT 56.450 1.630 61.310 2.680 ;
        RECT 62.430 1.630 67.290 2.680 ;
        RECT 68.410 1.630 73.270 2.680 ;
        RECT 74.390 1.630 79.250 2.680 ;
        RECT 80.370 1.630 84.770 2.680 ;
        RECT 85.890 1.630 90.750 2.680 ;
        RECT 91.870 1.630 96.730 2.680 ;
        RECT 97.850 1.630 102.710 2.680 ;
        RECT 103.830 1.630 108.690 2.680 ;
        RECT 109.810 1.630 114.670 2.680 ;
        RECT 115.790 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 132.150 2.680 ;
        RECT 133.270 1.630 138.130 2.680 ;
        RECT 139.250 1.630 144.110 2.680 ;
        RECT 145.230 1.630 150.090 2.680 ;
        RECT 151.210 1.630 156.070 2.680 ;
        RECT 157.190 1.630 161.590 2.680 ;
        RECT 162.710 1.630 167.570 2.680 ;
        RECT 168.690 1.630 173.550 2.680 ;
        RECT 174.670 1.630 179.530 2.680 ;
        RECT 180.650 1.630 185.510 2.680 ;
        RECT 186.630 1.630 191.490 2.680 ;
        RECT 192.610 1.630 197.470 2.680 ;
        RECT 198.590 1.630 202.990 2.680 ;
        RECT 204.110 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.950 2.680 ;
        RECT 216.070 1.630 220.930 2.680 ;
        RECT 222.050 1.630 226.910 2.680 ;
        RECT 228.030 1.630 232.890 2.680 ;
        RECT 234.010 1.630 238.870 2.680 ;
        RECT 239.990 1.630 244.390 2.680 ;
        RECT 245.510 1.630 250.370 2.680 ;
        RECT 251.490 1.630 256.350 2.680 ;
        RECT 257.470 1.630 262.330 2.680 ;
        RECT 263.450 1.630 268.310 2.680 ;
        RECT 269.430 1.630 274.290 2.680 ;
        RECT 275.410 1.630 279.810 2.680 ;
        RECT 280.930 1.630 285.790 2.680 ;
        RECT 286.910 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.750 2.680 ;
        RECT 298.870 1.630 303.730 2.680 ;
        RECT 304.850 1.630 309.710 2.680 ;
        RECT 310.830 1.630 315.690 2.680 ;
        RECT 316.810 1.630 321.210 2.680 ;
        RECT 322.330 1.630 327.190 2.680 ;
        RECT 328.310 1.630 333.170 2.680 ;
        RECT 334.290 1.630 339.150 2.680 ;
        RECT 340.270 1.630 345.130 2.680 ;
        RECT 346.250 1.630 351.110 2.680 ;
        RECT 352.230 1.630 357.090 2.680 ;
        RECT 358.210 1.630 362.610 2.680 ;
        RECT 363.730 1.630 368.590 2.680 ;
        RECT 369.710 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.550 2.680 ;
        RECT 381.670 1.630 386.530 2.680 ;
        RECT 387.650 1.630 392.510 2.680 ;
        RECT 393.630 1.630 398.030 2.680 ;
        RECT 399.150 1.630 404.010 2.680 ;
        RECT 405.130 1.630 409.990 2.680 ;
        RECT 411.110 1.630 415.970 2.680 ;
        RECT 417.090 1.630 421.950 2.680 ;
        RECT 423.070 1.630 427.930 2.680 ;
        RECT 429.050 1.630 433.910 2.680 ;
        RECT 435.030 1.630 439.430 2.680 ;
        RECT 440.550 1.630 445.410 2.680 ;
        RECT 446.530 1.630 451.390 2.680 ;
        RECT 452.510 1.630 457.370 2.680 ;
        RECT 458.490 1.630 463.350 2.680 ;
        RECT 464.470 1.630 469.330 2.680 ;
        RECT 470.450 1.630 475.310 2.680 ;
        RECT 476.430 1.630 480.830 2.680 ;
        RECT 481.950 1.630 486.810 2.680 ;
        RECT 487.930 1.630 492.790 2.680 ;
        RECT 493.910 1.630 498.770 2.680 ;
        RECT 499.890 1.630 504.750 2.680 ;
        RECT 505.870 1.630 510.730 2.680 ;
        RECT 511.850 1.630 516.250 2.680 ;
        RECT 517.370 1.630 522.230 2.680 ;
        RECT 523.350 1.630 528.210 2.680 ;
        RECT 529.330 1.630 534.190 2.680 ;
        RECT 535.310 1.630 540.170 2.680 ;
        RECT 541.290 1.630 546.150 2.680 ;
        RECT 547.270 1.630 552.130 2.680 ;
        RECT 553.250 1.630 557.650 2.680 ;
        RECT 558.770 1.630 563.630 2.680 ;
        RECT 564.750 1.630 569.610 2.680 ;
        RECT 570.730 1.630 575.590 2.680 ;
        RECT 576.710 1.630 581.570 2.680 ;
        RECT 582.690 1.630 587.550 2.680 ;
        RECT 588.670 1.630 593.530 2.680 ;
        RECT 594.650 1.630 599.050 2.680 ;
        RECT 600.170 1.630 605.030 2.680 ;
        RECT 606.150 1.630 611.010 2.680 ;
        RECT 612.130 1.630 616.990 2.680 ;
        RECT 618.110 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.950 2.680 ;
        RECT 630.070 1.630 634.470 2.680 ;
        RECT 635.590 1.630 640.450 2.680 ;
        RECT 641.570 1.630 646.430 2.680 ;
        RECT 647.550 1.630 652.410 2.680 ;
        RECT 653.530 1.630 658.390 2.680 ;
        RECT 659.510 1.630 664.370 2.680 ;
        RECT 665.490 1.630 670.350 2.680 ;
        RECT 671.470 1.630 675.870 2.680 ;
        RECT 676.990 1.630 681.850 2.680 ;
        RECT 682.970 1.630 687.830 2.680 ;
        RECT 688.950 1.630 693.810 2.680 ;
        RECT 694.930 1.630 699.790 2.680 ;
        RECT 700.910 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.750 2.680 ;
        RECT 712.870 1.630 717.270 2.680 ;
        RECT 718.390 1.630 723.250 2.680 ;
        RECT 724.370 1.630 729.230 2.680 ;
        RECT 730.350 1.630 735.210 2.680 ;
        RECT 736.330 1.630 741.190 2.680 ;
        RECT 742.310 1.630 747.170 2.680 ;
        RECT 748.290 1.630 752.690 2.680 ;
        RECT 753.810 1.630 758.670 2.680 ;
        RECT 759.790 1.630 764.650 2.680 ;
        RECT 765.770 1.630 770.630 2.680 ;
        RECT 771.750 1.630 776.610 2.680 ;
        RECT 777.730 1.630 782.590 2.680 ;
        RECT 783.710 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 800.070 2.680 ;
        RECT 801.190 1.630 806.050 2.680 ;
        RECT 807.170 1.630 812.030 2.680 ;
        RECT 813.150 1.630 818.010 2.680 ;
        RECT 819.130 1.630 823.990 2.680 ;
        RECT 825.110 1.630 829.970 2.680 ;
        RECT 831.090 1.630 835.490 2.680 ;
        RECT 836.610 1.630 841.470 2.680 ;
        RECT 842.590 1.630 847.450 2.680 ;
        RECT 848.570 1.630 853.430 2.680 ;
        RECT 854.550 1.630 859.410 2.680 ;
        RECT 860.530 1.630 865.390 2.680 ;
        RECT 866.510 1.630 870.910 2.680 ;
        RECT 872.030 1.630 876.890 2.680 ;
        RECT 878.010 1.630 882.870 2.680 ;
        RECT 883.990 1.630 888.850 2.680 ;
        RECT 889.970 1.630 894.830 2.680 ;
        RECT 895.950 1.630 900.810 2.680 ;
        RECT 901.930 1.630 906.790 2.680 ;
        RECT 907.910 1.630 912.310 2.680 ;
        RECT 913.430 1.630 918.290 2.680 ;
        RECT 919.410 1.630 924.270 2.680 ;
        RECT 925.390 1.630 930.250 2.680 ;
        RECT 931.370 1.630 936.230 2.680 ;
        RECT 937.350 1.630 942.210 2.680 ;
        RECT 943.330 1.630 948.190 2.680 ;
        RECT 949.310 1.630 953.710 2.680 ;
        RECT 954.830 1.630 959.690 2.680 ;
        RECT 960.810 1.630 965.670 2.680 ;
        RECT 966.790 1.630 971.650 2.680 ;
        RECT 972.770 1.630 977.630 2.680 ;
        RECT 978.750 1.630 983.610 2.680 ;
        RECT 984.730 1.630 989.130 2.680 ;
        RECT 990.250 1.630 995.110 2.680 ;
        RECT 996.230 1.630 1001.090 2.680 ;
        RECT 1002.210 1.630 1007.070 2.680 ;
        RECT 1008.190 1.630 1013.050 2.680 ;
        RECT 1014.170 1.630 1019.030 2.680 ;
        RECT 1020.150 1.630 1025.010 2.680 ;
        RECT 1026.130 1.630 1030.530 2.680 ;
        RECT 1031.650 1.630 1036.510 2.680 ;
        RECT 1037.630 1.630 1042.490 2.680 ;
        RECT 1043.610 1.630 1048.470 2.680 ;
        RECT 1049.590 1.630 1054.450 2.680 ;
        RECT 1055.570 1.630 1060.430 2.680 ;
        RECT 1061.550 1.630 1066.410 2.680 ;
        RECT 1067.530 1.630 1071.930 2.680 ;
        RECT 1073.050 1.630 1077.910 2.680 ;
        RECT 1079.030 1.630 1083.890 2.680 ;
        RECT 1085.010 1.630 1089.870 2.680 ;
        RECT 1090.990 1.630 1095.850 2.680 ;
        RECT 1096.970 1.630 1101.830 2.680 ;
        RECT 1102.950 1.630 1107.350 2.680 ;
        RECT 1108.470 1.630 1113.330 2.680 ;
        RECT 1114.450 1.630 1119.310 2.680 ;
        RECT 1120.430 1.630 1125.290 2.680 ;
        RECT 1126.410 1.630 1131.270 2.680 ;
        RECT 1132.390 1.630 1137.250 2.680 ;
        RECT 1138.370 1.630 1143.230 2.680 ;
        RECT 1144.350 1.630 1148.750 2.680 ;
        RECT 1149.870 1.630 1154.730 2.680 ;
        RECT 1155.850 1.630 1160.710 2.680 ;
        RECT 1161.830 1.630 1166.690 2.680 ;
        RECT 1167.810 1.630 1172.670 2.680 ;
        RECT 1173.790 1.630 1178.650 2.680 ;
        RECT 1179.770 1.630 1184.630 2.680 ;
        RECT 1185.750 1.630 1190.150 2.680 ;
        RECT 1191.270 1.630 1196.130 2.680 ;
        RECT 1197.250 1.630 1202.110 2.680 ;
        RECT 1203.230 1.630 1208.090 2.680 ;
        RECT 1209.210 1.630 1214.070 2.680 ;
        RECT 1215.190 1.630 1220.050 2.680 ;
        RECT 1221.170 1.630 1225.570 2.680 ;
        RECT 1226.690 1.630 1231.550 2.680 ;
        RECT 1232.670 1.630 1237.530 2.680 ;
        RECT 1238.650 1.630 1243.510 2.680 ;
        RECT 1244.630 1.630 1249.490 2.680 ;
        RECT 1250.610 1.630 1255.470 2.680 ;
        RECT 1256.590 1.630 1261.450 2.680 ;
        RECT 1262.570 1.630 1266.970 2.680 ;
        RECT 1268.090 1.630 1272.950 2.680 ;
        RECT 1274.070 1.630 1278.930 2.680 ;
        RECT 1280.050 1.630 1284.910 2.680 ;
        RECT 1286.030 1.630 1290.890 2.680 ;
        RECT 1292.010 1.630 1296.870 2.680 ;
        RECT 1297.990 1.630 1302.850 2.680 ;
        RECT 1303.970 1.630 1308.370 2.680 ;
        RECT 1309.490 1.630 1314.350 2.680 ;
        RECT 1315.470 1.630 1320.330 2.680 ;
        RECT 1321.450 1.630 1326.310 2.680 ;
        RECT 1327.430 1.630 1332.290 2.680 ;
        RECT 1333.410 1.630 1338.270 2.680 ;
        RECT 1339.390 1.630 1343.790 2.680 ;
        RECT 1344.910 1.630 1349.770 2.680 ;
        RECT 1350.890 1.630 1355.750 2.680 ;
        RECT 1356.870 1.630 1361.730 2.680 ;
        RECT 1362.850 1.630 1367.710 2.680 ;
        RECT 1368.830 1.630 1373.690 2.680 ;
        RECT 1374.810 1.630 1379.670 2.680 ;
        RECT 1380.790 1.630 1385.190 2.680 ;
        RECT 1386.310 1.630 1391.170 2.680 ;
        RECT 1392.290 1.630 1397.150 2.680 ;
        RECT 1398.270 1.630 1403.130 2.680 ;
        RECT 1404.250 1.630 1409.110 2.680 ;
        RECT 1410.230 1.630 1415.090 2.680 ;
        RECT 1416.210 1.630 1421.070 2.680 ;
        RECT 1422.190 1.630 1426.590 2.680 ;
        RECT 1427.710 1.630 1432.570 2.680 ;
        RECT 1433.690 1.630 1438.550 2.680 ;
        RECT 1439.670 1.630 1444.530 2.680 ;
        RECT 1445.650 1.630 1450.510 2.680 ;
        RECT 1451.630 1.630 1456.490 2.680 ;
        RECT 1457.610 1.630 1462.470 2.680 ;
        RECT 1463.590 1.630 1467.990 2.680 ;
        RECT 1469.110 1.630 1473.970 2.680 ;
        RECT 1475.090 1.630 1479.950 2.680 ;
        RECT 1481.070 1.630 1485.930 2.680 ;
        RECT 1487.050 1.630 1491.910 2.680 ;
        RECT 1493.030 1.630 1497.890 2.680 ;
        RECT 1499.010 1.630 1503.410 2.680 ;
        RECT 1504.530 1.630 1509.390 2.680 ;
        RECT 1510.510 1.630 1515.370 2.680 ;
        RECT 1516.490 1.630 1521.350 2.680 ;
        RECT 1522.470 1.630 1527.330 2.680 ;
        RECT 1528.450 1.630 1533.310 2.680 ;
        RECT 1534.430 1.630 1539.290 2.680 ;
        RECT 1540.410 1.630 1544.810 2.680 ;
        RECT 1545.930 1.630 1550.790 2.680 ;
        RECT 1551.910 1.630 1556.770 2.680 ;
        RECT 1557.890 1.630 1562.750 2.680 ;
        RECT 1563.870 1.630 1568.730 2.680 ;
        RECT 1569.850 1.630 1574.710 2.680 ;
        RECT 1575.830 1.630 1580.690 2.680 ;
        RECT 1581.810 1.630 1586.210 2.680 ;
        RECT 1587.330 1.630 1592.190 2.680 ;
        RECT 1593.310 1.630 1598.170 2.680 ;
        RECT 1599.290 1.630 1604.150 2.680 ;
        RECT 1605.270 1.630 1610.130 2.680 ;
        RECT 1611.250 1.630 1616.110 2.680 ;
        RECT 1617.230 1.630 1621.630 2.680 ;
        RECT 1622.750 1.630 1627.610 2.680 ;
        RECT 1628.730 1.630 1633.590 2.680 ;
        RECT 1634.710 1.630 1639.570 2.680 ;
        RECT 1640.690 1.630 1645.550 2.680 ;
        RECT 1646.670 1.630 1651.530 2.680 ;
        RECT 1652.650 1.630 1657.510 2.680 ;
        RECT 1658.630 1.630 1663.030 2.680 ;
        RECT 1664.150 1.630 1669.010 2.680 ;
        RECT 1670.130 1.630 1674.990 2.680 ;
        RECT 1676.110 1.630 1680.970 2.680 ;
        RECT 1682.090 1.630 1686.950 2.680 ;
        RECT 1688.070 1.630 1692.930 2.680 ;
        RECT 1694.050 1.630 1698.910 2.680 ;
        RECT 1700.030 1.630 1704.430 2.680 ;
        RECT 1705.550 1.630 1710.410 2.680 ;
        RECT 1711.530 1.630 1716.390 2.680 ;
        RECT 1717.510 1.630 1722.370 2.680 ;
        RECT 1723.490 1.630 1728.350 2.680 ;
        RECT 1729.470 1.630 1734.330 2.680 ;
        RECT 1735.450 1.630 1739.850 2.680 ;
        RECT 1740.970 1.630 1745.830 2.680 ;
        RECT 1746.950 1.630 1751.810 2.680 ;
        RECT 1752.930 1.630 1757.790 2.680 ;
        RECT 1758.910 1.630 1763.770 2.680 ;
        RECT 1764.890 1.630 1769.750 2.680 ;
        RECT 1770.870 1.630 1775.730 2.680 ;
        RECT 1776.850 1.630 1781.250 2.680 ;
        RECT 1782.370 1.630 1787.230 2.680 ;
        RECT 1788.350 1.630 1793.210 2.680 ;
        RECT 1794.330 1.630 1799.190 2.680 ;
        RECT 1800.310 1.630 1805.170 2.680 ;
        RECT 1806.290 1.630 1811.150 2.680 ;
        RECT 1812.270 1.630 1817.130 2.680 ;
        RECT 1818.250 1.630 1822.650 2.680 ;
        RECT 1823.770 1.630 1828.630 2.680 ;
        RECT 1829.750 1.630 1834.610 2.680 ;
        RECT 1835.730 1.630 1840.590 2.680 ;
        RECT 1841.710 1.630 1846.570 2.680 ;
        RECT 1847.690 1.630 1852.550 2.680 ;
        RECT 1853.670 1.630 1858.070 2.680 ;
        RECT 1859.190 1.630 1864.050 2.680 ;
        RECT 1865.170 1.630 1870.030 2.680 ;
        RECT 1871.150 1.630 1876.010 2.680 ;
        RECT 1877.130 1.630 1881.990 2.680 ;
        RECT 1883.110 1.630 1887.970 2.680 ;
        RECT 1889.090 1.630 1893.950 2.680 ;
        RECT 1895.070 1.630 1899.470 2.680 ;
        RECT 1900.590 1.630 1905.450 2.680 ;
        RECT 1906.570 1.630 1911.430 2.680 ;
        RECT 1912.550 1.630 1917.410 2.680 ;
        RECT 1918.530 1.630 1923.390 2.680 ;
        RECT 1924.510 1.630 1929.370 2.680 ;
        RECT 1930.490 1.630 1935.350 2.680 ;
        RECT 1936.470 1.630 1940.870 2.680 ;
        RECT 1941.990 1.630 1946.850 2.680 ;
        RECT 1947.970 1.630 1952.830 2.680 ;
        RECT 1953.950 1.630 1958.810 2.680 ;
        RECT 1959.930 1.630 1964.790 2.680 ;
        RECT 1965.910 1.630 1970.770 2.680 ;
        RECT 1971.890 1.630 1976.290 2.680 ;
        RECT 1977.410 1.630 1982.270 2.680 ;
        RECT 1983.390 1.630 1988.250 2.680 ;
        RECT 1989.370 1.630 1994.230 2.680 ;
        RECT 1995.350 1.630 2000.210 2.680 ;
        RECT 2001.330 1.630 2006.190 2.680 ;
        RECT 2007.310 1.630 2012.170 2.680 ;
        RECT 2013.290 1.630 2017.690 2.680 ;
        RECT 2018.810 1.630 2023.670 2.680 ;
        RECT 2024.790 1.630 2029.650 2.680 ;
        RECT 2030.770 1.630 2035.630 2.680 ;
        RECT 2036.750 1.630 2041.610 2.680 ;
        RECT 2042.730 1.630 2047.590 2.680 ;
        RECT 2048.710 1.630 2053.570 2.680 ;
        RECT 2054.690 1.630 2059.090 2.680 ;
        RECT 2060.210 1.630 2065.070 2.680 ;
        RECT 2066.190 1.630 2071.050 2.680 ;
        RECT 2072.170 1.630 2077.030 2.680 ;
        RECT 2078.150 1.630 2083.010 2.680 ;
        RECT 2084.130 1.630 2088.990 2.680 ;
        RECT 2090.110 1.630 2094.510 2.680 ;
        RECT 2095.630 1.630 2100.490 2.680 ;
        RECT 2101.610 1.630 2106.470 2.680 ;
        RECT 2107.590 1.630 2112.450 2.680 ;
        RECT 2113.570 1.630 2118.430 2.680 ;
        RECT 2119.550 1.630 2124.410 2.680 ;
        RECT 2125.530 1.630 2130.390 2.680 ;
        RECT 2131.510 1.630 2135.910 2.680 ;
        RECT 2137.030 1.630 2141.890 2.680 ;
        RECT 2143.010 1.630 2147.870 2.680 ;
        RECT 2148.990 1.630 2153.850 2.680 ;
        RECT 2154.970 1.630 2159.830 2.680 ;
        RECT 2160.950 1.630 2165.810 2.680 ;
        RECT 2166.930 1.630 2171.790 2.680 ;
        RECT 2172.910 1.630 2177.310 2.680 ;
        RECT 2178.430 1.630 2183.290 2.680 ;
        RECT 2184.410 1.630 2189.270 2.680 ;
        RECT 2190.390 1.630 2195.250 2.680 ;
        RECT 2196.370 1.630 2201.230 2.680 ;
        RECT 2202.350 1.630 2207.210 2.680 ;
        RECT 2208.330 1.630 2212.730 2.680 ;
        RECT 2213.850 1.630 2218.710 2.680 ;
        RECT 2219.830 1.630 2224.690 2.680 ;
        RECT 2225.810 1.630 2230.670 2.680 ;
        RECT 2231.790 1.630 2236.650 2.680 ;
        RECT 2237.770 1.630 2242.630 2.680 ;
        RECT 2243.750 1.630 2248.610 2.680 ;
        RECT 2249.730 1.630 2254.130 2.680 ;
        RECT 2255.250 1.630 2260.110 2.680 ;
        RECT 2261.230 1.630 2266.090 2.680 ;
        RECT 2267.210 1.630 2272.070 2.680 ;
        RECT 2273.190 1.630 2278.050 2.680 ;
        RECT 2279.170 1.630 2284.030 2.680 ;
        RECT 2285.150 1.630 2290.010 2.680 ;
        RECT 2291.130 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2301.510 2.680 ;
        RECT 2302.630 1.630 2307.490 2.680 ;
        RECT 2308.610 1.630 2313.470 2.680 ;
        RECT 2314.590 1.630 2319.450 2.680 ;
        RECT 2320.570 1.630 2325.430 2.680 ;
        RECT 2326.550 1.630 2330.950 2.680 ;
        RECT 2332.070 1.630 2336.930 2.680 ;
        RECT 2338.050 1.630 2342.910 2.680 ;
        RECT 2344.030 1.630 2348.890 2.680 ;
        RECT 2350.010 1.630 2354.870 2.680 ;
        RECT 2355.990 1.630 2360.850 2.680 ;
        RECT 2361.970 1.630 2366.830 2.680 ;
        RECT 2367.950 1.630 2372.350 2.680 ;
        RECT 2373.470 1.630 2378.330 2.680 ;
        RECT 2379.450 1.630 2384.310 2.680 ;
        RECT 2385.430 1.630 2390.290 2.680 ;
        RECT 2391.410 1.630 2396.270 2.680 ;
        RECT 2397.390 1.630 2402.250 2.680 ;
        RECT 2403.370 1.630 2408.230 2.680 ;
        RECT 2409.350 1.630 2413.750 2.680 ;
        RECT 2414.870 1.630 2419.730 2.680 ;
        RECT 2420.850 1.630 2425.710 2.680 ;
        RECT 2426.830 1.630 2431.690 2.680 ;
        RECT 2432.810 1.630 2437.670 2.680 ;
        RECT 2438.790 1.630 2443.650 2.680 ;
        RECT 2444.770 1.630 2449.170 2.680 ;
        RECT 2450.290 1.630 2455.150 2.680 ;
        RECT 2456.270 1.630 2461.130 2.680 ;
        RECT 2462.250 1.630 2467.110 2.680 ;
        RECT 2468.230 1.630 2473.090 2.680 ;
        RECT 2474.210 1.630 2479.070 2.680 ;
        RECT 2480.190 1.630 2485.050 2.680 ;
        RECT 2486.170 1.630 2490.570 2.680 ;
        RECT 2491.690 1.630 2496.550 2.680 ;
        RECT 2497.670 1.630 2502.530 2.680 ;
        RECT 2503.650 1.630 2508.510 2.680 ;
        RECT 2509.630 1.630 2514.490 2.680 ;
        RECT 2515.610 1.630 2520.470 2.680 ;
        RECT 2521.590 1.630 2526.450 2.680 ;
        RECT 2527.570 1.630 2531.970 2.680 ;
        RECT 2533.090 1.630 2537.950 2.680 ;
        RECT 2539.070 1.630 2543.930 2.680 ;
        RECT 2545.050 1.630 2549.910 2.680 ;
        RECT 2551.030 1.630 2555.890 2.680 ;
        RECT 2557.010 1.630 2561.870 2.680 ;
        RECT 2562.990 1.630 2567.390 2.680 ;
        RECT 2568.510 1.630 2573.370 2.680 ;
        RECT 2574.490 1.630 2579.350 2.680 ;
        RECT 2580.470 1.630 2585.330 2.680 ;
        RECT 2586.450 1.630 2591.310 2.680 ;
        RECT 2592.430 1.630 2597.290 2.680 ;
        RECT 2598.410 1.630 2603.270 2.680 ;
        RECT 2604.390 1.630 2608.790 2.680 ;
        RECT 2609.910 1.630 2614.770 2.680 ;
        RECT 2615.890 1.630 2620.750 2.680 ;
        RECT 2621.870 1.630 2626.730 2.680 ;
        RECT 2627.850 1.630 2632.710 2.680 ;
        RECT 2633.830 1.630 2638.690 2.680 ;
        RECT 2639.810 1.630 2644.670 2.680 ;
        RECT 2645.790 1.630 2650.190 2.680 ;
        RECT 2651.310 1.630 2656.170 2.680 ;
        RECT 2657.290 1.630 2662.150 2.680 ;
        RECT 2663.270 1.630 2668.130 2.680 ;
        RECT 2669.250 1.630 2674.110 2.680 ;
        RECT 2675.230 1.630 2680.090 2.680 ;
        RECT 2681.210 1.630 2685.610 2.680 ;
        RECT 2686.730 1.630 2691.590 2.680 ;
        RECT 2692.710 1.630 2697.570 2.680 ;
        RECT 2698.690 1.630 2703.550 2.680 ;
        RECT 2704.670 1.630 2709.530 2.680 ;
        RECT 2710.650 1.630 2715.510 2.680 ;
        RECT 2716.630 1.630 2721.490 2.680 ;
        RECT 2722.610 1.630 2727.010 2.680 ;
        RECT 2728.130 1.630 2732.990 2.680 ;
        RECT 2734.110 1.630 2738.970 2.680 ;
        RECT 2740.090 1.630 2744.950 2.680 ;
        RECT 2746.070 1.630 2750.930 2.680 ;
        RECT 2752.050 1.630 2756.910 2.680 ;
        RECT 2758.030 1.630 2762.890 2.680 ;
        RECT 2764.010 1.630 2768.410 2.680 ;
        RECT 2769.530 1.630 2774.390 2.680 ;
        RECT 2775.510 1.630 2780.370 2.680 ;
        RECT 2781.490 1.630 2786.350 2.680 ;
        RECT 2787.470 1.630 2792.330 2.680 ;
        RECT 2793.450 1.630 2798.310 2.680 ;
        RECT 2799.430 1.630 2803.830 2.680 ;
        RECT 2804.950 1.630 2809.810 2.680 ;
        RECT 2810.930 1.630 2815.790 2.680 ;
        RECT 2816.910 1.630 2821.770 2.680 ;
        RECT 2822.890 1.630 2827.750 2.680 ;
        RECT 2828.870 1.630 2833.730 2.680 ;
        RECT 2834.850 1.630 2839.710 2.680 ;
        RECT 2840.830 1.630 2845.230 2.680 ;
        RECT 2846.350 1.630 2851.210 2.680 ;
        RECT 2852.330 1.630 2857.190 2.680 ;
        RECT 2858.310 1.630 2863.170 2.680 ;
        RECT 2864.290 1.630 2869.150 2.680 ;
        RECT 2870.270 1.630 2875.130 2.680 ;
        RECT 2876.250 1.630 2881.110 2.680 ;
        RECT 2882.230 1.630 2886.630 2.680 ;
        RECT 2887.750 1.630 2892.610 2.680 ;
        RECT 2893.730 1.630 2898.590 2.680 ;
        RECT 2899.710 1.630 2904.570 2.680 ;
        RECT 2905.690 1.630 2910.550 2.680 ;
        RECT 2911.670 1.630 2916.530 2.680 ;
      LAYER met3 ;
        RECT 2.400 3487.700 2917.600 3508.965 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.400 3420.380 2917.600 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.400 3354.420 2917.600 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.400 3287.780 2917.600 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.400 3221.140 2917.600 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.400 3155.180 2917.600 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.400 3088.540 2917.600 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.400 3021.900 2917.600 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.400 2955.940 2917.600 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.400 2889.300 2917.600 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.400 2822.660 2917.600 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.400 2756.700 2917.600 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.400 2690.060 2917.600 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.400 2623.420 2917.600 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.400 2557.460 2917.600 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.400 2490.820 2917.600 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.400 2424.180 2917.600 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.400 2358.220 2917.600 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.400 2291.580 2917.600 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.400 2224.940 2917.600 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.400 2158.980 2917.600 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.400 2092.340 2917.600 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.400 2025.700 2917.600 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1959.740 2917.600 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.400 1893.100 2917.600 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.400 1693.860 2917.600 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.400 1627.220 2917.600 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.400 1561.260 2917.600 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.400 1494.620 2917.600 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.400 1427.980 2917.600 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.400 1362.020 2917.600 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.400 1295.380 2917.600 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.400 1228.740 2917.600 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.400 1162.780 2917.600 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.400 1096.140 2917.600 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.400 1029.500 2917.600 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.400 963.540 2917.600 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.400 896.900 2917.600 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.400 830.260 2917.600 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.400 764.300 2917.600 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.400 697.660 2917.600 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.400 631.020 2917.600 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.400 565.060 2917.600 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.400 498.420 2917.600 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.400 431.780 2917.600 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.400 365.820 2917.600 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.400 299.180 2917.600 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.400 232.540 2917.600 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.400 166.580 2917.600 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.400 99.940 2917.600 161.180 ;
        RECT 2.400 97.940 2917.200 99.940 ;
        RECT 2.400 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 2.400 33.980 2917.600 95.900 ;
        RECT 2.400 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 2.400 10.715 2917.600 31.300 ;
      LAYER met4 ;
        RECT 67.075 3382.500 184.570 3488.760 ;
        RECT 188.470 3382.500 203.170 3488.760 ;
        RECT 67.075 3362.560 203.170 3382.500 ;
        RECT 67.075 3309.600 106.150 3362.560 ;
        RECT 113.730 3323.340 203.170 3362.560 ;
        RECT 113.730 3309.600 184.570 3323.340 ;
        RECT 67.075 3068.500 184.570 3309.600 ;
        RECT 188.470 3068.500 203.170 3323.340 ;
        RECT 67.075 3049.760 203.170 3068.500 ;
        RECT 67.075 2994.080 106.150 3049.760 ;
        RECT 113.730 3009.340 203.170 3049.760 ;
        RECT 113.730 2994.080 184.570 3009.340 ;
        RECT 67.075 2928.420 184.570 2994.080 ;
        RECT 188.470 2928.420 203.170 3009.340 ;
        RECT 207.070 3395.200 364.570 3488.760 ;
        RECT 207.070 3312.320 268.070 3395.200 ;
        RECT 271.970 3378.565 364.570 3395.200 ;
        RECT 368.470 3378.565 383.170 3488.760 ;
        RECT 387.070 3382.500 544.570 3488.760 ;
        RECT 548.470 3382.500 563.170 3488.760 ;
        RECT 567.070 3427.260 743.170 3488.760 ;
        RECT 747.070 3427.260 904.570 3488.760 ;
        RECT 567.070 3397.920 904.570 3427.260 ;
        RECT 567.070 3382.500 612.150 3397.920 ;
        RECT 387.070 3378.565 612.150 3382.500 ;
        RECT 271.970 3323.340 612.150 3378.565 ;
        RECT 271.970 3312.320 544.570 3323.340 ;
        RECT 207.070 3277.395 544.570 3312.320 ;
        RECT 207.070 3079.680 364.570 3277.395 ;
        RECT 207.070 2996.800 268.070 3079.680 ;
        RECT 271.970 3064.565 364.570 3079.680 ;
        RECT 368.470 3064.565 383.170 3277.395 ;
        RECT 387.070 3253.760 544.570 3277.395 ;
        RECT 387.070 3162.720 465.870 3253.760 ;
        RECT 469.770 3162.720 485.190 3253.760 ;
        RECT 489.090 3250.580 544.570 3253.760 ;
        RECT 548.470 3250.580 563.170 3323.340 ;
        RECT 567.070 3309.600 612.150 3323.340 ;
        RECT 616.050 3309.600 631.470 3397.920 ;
        RECT 635.370 3309.600 904.570 3397.920 ;
        RECT 567.070 3277.395 904.570 3309.600 ;
        RECT 567.070 3253.760 724.570 3277.395 ;
        RECT 567.070 3250.580 636.070 3253.760 ;
        RECT 489.090 3162.720 636.070 3250.580 ;
        RECT 639.970 3162.720 655.390 3253.760 ;
        RECT 659.290 3237.500 724.570 3253.760 ;
        RECT 728.470 3237.500 743.170 3277.395 ;
        RECT 747.070 3253.760 904.570 3277.395 ;
        RECT 747.070 3237.500 786.030 3253.760 ;
        RECT 659.290 3178.340 786.030 3237.500 ;
        RECT 659.290 3162.720 724.570 3178.340 ;
        RECT 387.070 3146.275 724.570 3162.720 ;
        RECT 387.070 3068.500 544.570 3146.275 ;
        RECT 548.470 3068.500 563.170 3146.275 ;
        RECT 567.070 3113.260 724.570 3146.275 ;
        RECT 728.470 3113.260 743.170 3178.340 ;
        RECT 747.070 3162.720 786.030 3178.340 ;
        RECT 789.930 3162.720 805.350 3253.760 ;
        RECT 809.250 3162.720 904.570 3253.760 ;
        RECT 747.070 3113.260 904.570 3162.720 ;
        RECT 567.070 3085.120 904.570 3113.260 ;
        RECT 567.070 3072.960 611.230 3085.120 ;
        RECT 615.130 3073.360 630.550 3085.120 ;
        RECT 634.450 3073.360 904.570 3085.120 ;
        RECT 616.050 3072.960 630.550 3073.360 ;
        RECT 567.070 3068.500 612.150 3072.960 ;
        RECT 387.070 3064.565 612.150 3068.500 ;
        RECT 271.970 3009.340 612.150 3064.565 ;
        RECT 271.970 2996.800 544.570 3009.340 ;
        RECT 207.070 2963.395 544.570 2996.800 ;
        RECT 207.070 2928.420 364.570 2963.395 ;
        RECT 67.075 2839.340 364.570 2928.420 ;
        RECT 67.075 2754.500 184.570 2839.340 ;
        RECT 188.470 2754.500 203.170 2839.340 ;
        RECT 67.075 2734.240 203.170 2754.500 ;
        RECT 67.075 2681.280 106.150 2734.240 ;
        RECT 113.730 2695.340 203.170 2734.240 ;
        RECT 113.730 2681.280 184.570 2695.340 ;
        RECT 67.075 2614.420 184.570 2681.280 ;
        RECT 188.470 2614.420 203.170 2695.340 ;
        RECT 207.070 2769.600 364.570 2839.340 ;
        RECT 207.070 2681.280 268.070 2769.600 ;
        RECT 271.970 2750.565 364.570 2769.600 ;
        RECT 368.470 2750.565 383.170 2963.395 ;
        RECT 387.070 2958.340 544.570 2963.395 ;
        RECT 548.470 2958.340 563.170 3009.340 ;
        RECT 567.070 2994.080 612.150 3009.340 ;
        RECT 616.050 2994.080 631.470 3072.960 ;
        RECT 635.370 2994.080 904.570 3073.360 ;
        RECT 567.070 2973.600 904.570 2994.080 ;
        RECT 567.070 2958.340 613.990 2973.600 ;
        RECT 387.070 2956.000 613.990 2958.340 ;
        RECT 617.890 2959.600 633.310 2973.600 ;
        RECT 637.210 2963.395 904.570 2973.600 ;
        RECT 637.210 2960.000 724.570 2963.395 ;
        RECT 617.890 2956.000 634.230 2959.600 ;
        RECT 387.070 2947.840 634.230 2956.000 ;
        RECT 638.130 2947.840 653.550 2960.000 ;
        RECT 657.450 2947.840 724.570 2960.000 ;
        RECT 387.070 2932.800 724.570 2947.840 ;
        RECT 387.070 2844.480 465.870 2932.800 ;
        RECT 469.770 2844.480 485.190 2932.800 ;
        RECT 489.090 2853.920 636.070 2932.800 ;
        RECT 639.970 2853.920 655.390 2932.800 ;
        RECT 659.290 2917.500 724.570 2932.800 ;
        RECT 728.470 2917.500 743.170 2963.395 ;
        RECT 747.070 2932.800 904.570 2963.395 ;
        RECT 747.070 2917.500 786.030 2932.800 ;
        RECT 659.290 2858.340 786.030 2917.500 ;
        RECT 489.090 2844.480 634.230 2853.920 ;
        RECT 639.970 2853.520 653.550 2853.920 ;
        RECT 659.290 2853.520 743.170 2858.340 ;
        RECT 387.070 2841.760 634.230 2844.480 ;
        RECT 638.130 2841.760 653.550 2853.520 ;
        RECT 657.450 2849.235 743.170 2853.520 ;
        RECT 657.450 2841.760 724.570 2849.235 ;
        RECT 387.070 2837.715 724.570 2841.760 ;
        RECT 387.070 2754.500 544.570 2837.715 ;
        RECT 548.470 2754.500 563.170 2837.715 ;
        RECT 567.070 2799.260 724.570 2837.715 ;
        RECT 728.470 2799.260 743.170 2849.235 ;
        RECT 747.070 2853.120 786.030 2858.340 ;
        RECT 789.930 2859.360 805.350 2932.800 ;
        RECT 789.930 2853.120 793.390 2859.360 ;
        RECT 747.070 2844.480 793.390 2853.120 ;
        RECT 800.970 2853.120 805.350 2859.360 ;
        RECT 809.250 2853.120 904.570 2932.800 ;
        RECT 800.970 2844.480 904.570 2853.120 ;
        RECT 747.070 2799.260 904.570 2844.480 ;
        RECT 567.070 2769.600 904.570 2799.260 ;
        RECT 567.070 2754.500 612.150 2769.600 ;
        RECT 387.070 2750.565 612.150 2754.500 ;
        RECT 271.970 2695.340 612.150 2750.565 ;
        RECT 271.970 2681.280 544.570 2695.340 ;
        RECT 207.070 2649.395 544.570 2681.280 ;
        RECT 207.070 2614.420 364.570 2649.395 ;
        RECT 67.075 2525.340 364.570 2614.420 ;
        RECT 67.075 2440.500 184.570 2525.340 ;
        RECT 188.470 2440.500 203.170 2525.340 ;
        RECT 67.075 2421.440 203.170 2440.500 ;
        RECT 67.075 2365.760 106.150 2421.440 ;
        RECT 113.730 2381.340 203.170 2421.440 ;
        RECT 113.730 2365.760 184.570 2381.340 ;
        RECT 67.075 2300.420 184.570 2365.760 ;
        RECT 188.470 2300.420 203.170 2381.340 ;
        RECT 207.070 2454.080 364.570 2525.340 ;
        RECT 207.070 2365.760 268.070 2454.080 ;
        RECT 271.970 2436.565 364.570 2454.080 ;
        RECT 368.470 2436.565 383.170 2649.395 ;
        RECT 387.070 2644.340 544.570 2649.395 ;
        RECT 548.470 2644.340 563.170 2695.340 ;
        RECT 567.070 2681.280 612.150 2695.340 ;
        RECT 616.050 2681.280 631.470 2769.600 ;
        RECT 635.370 2681.280 904.570 2769.600 ;
        RECT 567.070 2660.800 904.570 2681.280 ;
        RECT 567.070 2644.340 613.990 2660.800 ;
        RECT 387.070 2635.040 613.990 2644.340 ;
        RECT 617.890 2635.040 633.310 2660.800 ;
        RECT 637.210 2649.395 904.570 2660.800 ;
        RECT 637.210 2635.040 724.570 2649.395 ;
        RECT 387.070 2625.440 724.570 2635.040 ;
        RECT 387.070 2534.400 465.870 2625.440 ;
        RECT 469.770 2534.400 485.190 2625.440 ;
        RECT 489.090 2534.400 636.070 2625.440 ;
        RECT 639.970 2534.400 655.390 2625.440 ;
        RECT 659.290 2609.500 724.570 2625.440 ;
        RECT 728.470 2609.500 743.170 2649.395 ;
        RECT 747.070 2625.440 904.570 2649.395 ;
        RECT 747.070 2609.500 786.030 2625.440 ;
        RECT 659.290 2550.340 786.030 2609.500 ;
        RECT 659.290 2541.235 743.170 2550.340 ;
        RECT 659.290 2534.400 724.570 2541.235 ;
        RECT 387.070 2523.715 724.570 2534.400 ;
        RECT 387.070 2440.500 544.570 2523.715 ;
        RECT 548.470 2440.500 563.170 2523.715 ;
        RECT 567.070 2485.260 724.570 2523.715 ;
        RECT 728.470 2485.260 743.170 2541.235 ;
        RECT 747.070 2534.400 786.030 2550.340 ;
        RECT 789.930 2534.400 805.350 2625.440 ;
        RECT 809.250 2534.400 904.570 2625.440 ;
        RECT 747.070 2485.260 904.570 2534.400 ;
        RECT 567.070 2456.800 904.570 2485.260 ;
        RECT 567.070 2440.500 612.150 2456.800 ;
        RECT 387.070 2436.565 612.150 2440.500 ;
        RECT 271.970 2381.340 612.150 2436.565 ;
        RECT 271.970 2365.760 544.570 2381.340 ;
        RECT 207.070 2335.395 544.570 2365.760 ;
        RECT 207.070 2300.420 364.570 2335.395 ;
        RECT 67.075 2211.340 364.570 2300.420 ;
        RECT 67.075 2126.500 184.570 2211.340 ;
        RECT 188.470 2126.500 203.170 2211.340 ;
        RECT 67.075 2105.920 203.170 2126.500 ;
        RECT 67.075 2052.960 106.150 2105.920 ;
        RECT 113.730 2067.340 203.170 2105.920 ;
        RECT 113.730 2052.960 184.570 2067.340 ;
        RECT 67.075 1986.420 184.570 2052.960 ;
        RECT 188.470 1986.420 203.170 2067.340 ;
        RECT 207.070 2138.560 364.570 2211.340 ;
        RECT 207.070 2055.680 268.070 2138.560 ;
        RECT 271.970 2122.565 364.570 2138.560 ;
        RECT 368.470 2122.565 383.170 2335.395 ;
        RECT 387.070 2330.340 544.570 2335.395 ;
        RECT 548.470 2330.340 563.170 2381.340 ;
        RECT 567.070 2365.760 612.150 2381.340 ;
        RECT 616.050 2365.760 631.470 2456.800 ;
        RECT 635.370 2365.760 904.570 2456.800 ;
        RECT 567.070 2345.280 904.570 2365.760 ;
        RECT 567.070 2330.340 613.990 2345.280 ;
        RECT 387.070 2322.240 613.990 2330.340 ;
        RECT 617.890 2322.240 633.310 2345.280 ;
        RECT 637.210 2335.395 904.570 2345.280 ;
        RECT 637.210 2322.240 724.570 2335.395 ;
        RECT 387.070 2309.920 724.570 2322.240 ;
        RECT 387.070 2221.600 465.870 2309.920 ;
        RECT 469.770 2221.600 485.190 2309.920 ;
        RECT 489.090 2221.600 636.070 2309.920 ;
        RECT 639.970 2221.600 655.390 2309.920 ;
        RECT 659.290 2295.500 724.570 2309.920 ;
        RECT 728.470 2295.500 743.170 2335.395 ;
        RECT 747.070 2309.920 904.570 2335.395 ;
        RECT 747.070 2295.500 786.030 2309.920 ;
        RECT 659.290 2236.340 786.030 2295.500 ;
        RECT 659.290 2227.235 743.170 2236.340 ;
        RECT 659.290 2221.600 724.570 2227.235 ;
        RECT 387.070 2210.030 724.570 2221.600 ;
        RECT 387.070 2209.715 563.170 2210.030 ;
        RECT 387.070 2126.500 544.570 2209.715 ;
        RECT 548.470 2126.500 563.170 2209.715 ;
        RECT 567.070 2171.260 724.570 2210.030 ;
        RECT 728.470 2171.260 743.170 2227.235 ;
        RECT 747.070 2221.600 786.030 2236.340 ;
        RECT 789.930 2221.600 805.350 2309.920 ;
        RECT 809.250 2221.600 904.570 2309.920 ;
        RECT 747.070 2171.260 904.570 2221.600 ;
        RECT 567.070 2141.280 904.570 2171.260 ;
        RECT 567.070 2126.500 612.150 2141.280 ;
        RECT 387.070 2122.565 612.150 2126.500 ;
        RECT 271.970 2067.340 612.150 2122.565 ;
        RECT 271.970 2055.680 544.570 2067.340 ;
        RECT 207.070 2021.395 544.570 2055.680 ;
        RECT 207.070 1986.420 364.570 2021.395 ;
        RECT 67.075 1983.520 364.570 1986.420 ;
        RECT 67.075 1922.400 301.190 1983.520 ;
        RECT 305.090 1922.400 364.570 1983.520 ;
        RECT 67.075 1897.340 364.570 1922.400 ;
        RECT 67.075 1812.500 184.570 1897.340 ;
        RECT 188.470 1812.500 203.170 1897.340 ;
        RECT 67.075 1793.120 203.170 1812.500 ;
        RECT 67.075 1737.440 106.150 1793.120 ;
        RECT 113.730 1753.340 203.170 1793.120 ;
        RECT 113.730 1737.440 184.570 1753.340 ;
        RECT 67.075 1672.420 184.570 1737.440 ;
        RECT 188.470 1672.420 203.170 1753.340 ;
        RECT 207.070 1828.480 364.570 1897.340 ;
        RECT 207.070 1740.160 268.070 1828.480 ;
        RECT 271.970 1808.565 364.570 1828.480 ;
        RECT 368.470 1808.565 383.170 2021.395 ;
        RECT 387.070 2016.340 544.570 2021.395 ;
        RECT 548.470 2016.340 563.170 2067.340 ;
        RECT 567.070 2052.960 612.150 2067.340 ;
        RECT 616.050 2052.960 631.470 2141.280 ;
        RECT 635.370 2052.960 904.570 2141.280 ;
        RECT 567.070 2032.480 904.570 2052.960 ;
        RECT 567.070 2016.340 613.990 2032.480 ;
        RECT 387.070 2006.720 613.990 2016.340 ;
        RECT 617.890 2006.720 633.310 2032.480 ;
        RECT 637.210 2021.395 904.570 2032.480 ;
        RECT 637.210 2006.720 724.570 2021.395 ;
        RECT 387.070 1997.120 724.570 2006.720 ;
        RECT 387.070 1906.080 465.870 1997.120 ;
        RECT 469.770 1906.080 485.190 1997.120 ;
        RECT 489.090 1906.080 636.070 1997.120 ;
        RECT 639.970 1906.080 655.390 1997.120 ;
        RECT 659.290 1981.500 724.570 1997.120 ;
        RECT 728.470 1981.500 743.170 2021.395 ;
        RECT 747.070 1997.120 904.570 2021.395 ;
        RECT 747.070 1981.500 786.030 1997.120 ;
        RECT 659.290 1922.340 786.030 1981.500 ;
        RECT 659.290 1913.235 743.170 1922.340 ;
        RECT 659.290 1906.080 724.570 1913.235 ;
        RECT 387.070 1895.715 724.570 1906.080 ;
        RECT 387.070 1812.500 544.570 1895.715 ;
        RECT 548.470 1812.500 563.170 1895.715 ;
        RECT 567.070 1857.260 724.570 1895.715 ;
        RECT 728.470 1857.260 743.170 1913.235 ;
        RECT 747.070 1906.080 786.030 1922.340 ;
        RECT 789.930 1906.080 805.350 1997.120 ;
        RECT 809.250 1906.080 904.570 1997.120 ;
        RECT 747.070 1857.260 904.570 1906.080 ;
        RECT 567.070 1828.480 904.570 1857.260 ;
        RECT 567.070 1812.500 612.150 1828.480 ;
        RECT 387.070 1808.565 612.150 1812.500 ;
        RECT 271.970 1753.340 612.150 1808.565 ;
        RECT 271.970 1740.160 544.570 1753.340 ;
        RECT 207.070 1707.395 544.570 1740.160 ;
        RECT 207.070 1672.420 364.570 1707.395 ;
        RECT 67.075 1583.340 364.570 1672.420 ;
        RECT 67.075 1498.500 184.570 1583.340 ;
        RECT 188.470 1498.500 203.170 1583.340 ;
        RECT 67.075 1477.600 203.170 1498.500 ;
        RECT 67.075 1424.640 106.150 1477.600 ;
        RECT 113.730 1439.340 203.170 1477.600 ;
        RECT 113.730 1424.640 184.570 1439.340 ;
        RECT 67.075 1358.420 184.570 1424.640 ;
        RECT 188.470 1358.420 203.170 1439.340 ;
        RECT 207.070 1512.960 364.570 1583.340 ;
        RECT 207.070 1424.640 268.070 1512.960 ;
        RECT 271.970 1494.565 364.570 1512.960 ;
        RECT 368.470 1494.565 383.170 1707.395 ;
        RECT 387.070 1702.340 544.570 1707.395 ;
        RECT 548.470 1702.340 563.170 1753.340 ;
        RECT 567.070 1737.440 612.150 1753.340 ;
        RECT 616.050 1737.440 631.470 1828.480 ;
        RECT 635.370 1737.440 904.570 1828.480 ;
        RECT 567.070 1716.960 904.570 1737.440 ;
        RECT 567.070 1702.340 613.990 1716.960 ;
        RECT 387.070 1693.920 613.990 1702.340 ;
        RECT 617.890 1693.920 633.310 1716.960 ;
        RECT 637.210 1707.395 904.570 1716.960 ;
        RECT 637.210 1693.920 724.570 1707.395 ;
        RECT 387.070 1684.320 724.570 1693.920 ;
        RECT 387.070 1681.600 606.630 1684.320 ;
        RECT 387.070 1593.280 465.870 1681.600 ;
        RECT 469.770 1593.280 485.190 1681.600 ;
        RECT 489.090 1672.160 606.630 1681.600 ;
        RECT 610.530 1672.160 625.950 1684.320 ;
        RECT 629.850 1672.960 724.570 1684.320 ;
        RECT 629.850 1672.160 636.070 1672.960 ;
        RECT 489.090 1593.280 636.070 1672.160 ;
        RECT 639.970 1593.280 655.390 1672.960 ;
        RECT 659.290 1667.500 724.570 1672.960 ;
        RECT 728.470 1667.500 743.170 1707.395 ;
        RECT 747.070 1681.600 904.570 1707.395 ;
        RECT 747.070 1672.960 793.390 1681.600 ;
        RECT 747.070 1667.500 786.030 1672.960 ;
        RECT 659.290 1608.340 786.030 1667.500 ;
        RECT 659.290 1599.235 743.170 1608.340 ;
        RECT 659.290 1593.280 724.570 1599.235 ;
        RECT 387.070 1581.715 724.570 1593.280 ;
        RECT 387.070 1498.500 544.570 1581.715 ;
        RECT 548.470 1498.500 563.170 1581.715 ;
        RECT 567.070 1543.260 724.570 1581.715 ;
        RECT 728.470 1543.260 743.170 1599.235 ;
        RECT 747.070 1593.280 786.030 1608.340 ;
        RECT 789.930 1666.720 793.390 1672.960 ;
        RECT 800.970 1672.960 904.570 1681.600 ;
        RECT 800.970 1666.720 805.350 1672.960 ;
        RECT 789.930 1593.280 805.350 1666.720 ;
        RECT 809.250 1593.280 904.570 1672.960 ;
        RECT 747.070 1543.260 904.570 1593.280 ;
        RECT 567.070 1512.960 904.570 1543.260 ;
        RECT 567.070 1498.500 612.150 1512.960 ;
        RECT 387.070 1494.565 612.150 1498.500 ;
        RECT 271.970 1439.340 612.150 1494.565 ;
        RECT 271.970 1424.640 544.570 1439.340 ;
        RECT 207.070 1393.395 544.570 1424.640 ;
        RECT 207.070 1358.420 364.570 1393.395 ;
        RECT 67.075 1269.340 364.570 1358.420 ;
        RECT 67.075 1184.500 184.570 1269.340 ;
        RECT 188.470 1184.500 203.170 1269.340 ;
        RECT 67.075 1164.800 203.170 1184.500 ;
        RECT 67.075 1109.120 106.150 1164.800 ;
        RECT 113.730 1125.340 203.170 1164.800 ;
        RECT 113.730 1109.120 184.570 1125.340 ;
        RECT 67.075 1044.420 184.570 1109.120 ;
        RECT 188.470 1044.420 203.170 1125.340 ;
        RECT 207.070 1197.440 364.570 1269.340 ;
        RECT 207.070 1109.120 268.070 1197.440 ;
        RECT 271.970 1180.565 364.570 1197.440 ;
        RECT 368.470 1180.565 383.170 1393.395 ;
        RECT 387.070 1388.340 544.570 1393.395 ;
        RECT 548.470 1388.340 563.170 1439.340 ;
        RECT 567.070 1424.640 612.150 1439.340 ;
        RECT 616.050 1424.640 631.470 1512.960 ;
        RECT 635.370 1424.640 904.570 1512.960 ;
        RECT 567.070 1404.160 904.570 1424.640 ;
        RECT 567.070 1388.340 613.990 1404.160 ;
        RECT 387.070 1378.400 613.990 1388.340 ;
        RECT 617.890 1378.400 633.310 1404.160 ;
        RECT 637.210 1393.395 904.570 1404.160 ;
        RECT 637.210 1378.400 724.570 1393.395 ;
        RECT 387.070 1368.800 724.570 1378.400 ;
        RECT 387.070 1280.480 465.870 1368.800 ;
        RECT 469.770 1280.480 485.190 1368.800 ;
        RECT 489.090 1289.920 636.070 1368.800 ;
        RECT 639.970 1289.920 655.390 1368.800 ;
        RECT 659.290 1353.500 724.570 1368.800 ;
        RECT 728.470 1353.500 743.170 1393.395 ;
        RECT 747.070 1368.800 904.570 1393.395 ;
        RECT 747.070 1353.500 786.030 1368.800 ;
        RECT 659.290 1294.340 786.030 1353.500 ;
        RECT 489.090 1280.480 634.230 1289.920 ;
        RECT 639.970 1289.520 653.550 1289.920 ;
        RECT 659.290 1289.520 743.170 1294.340 ;
        RECT 387.070 1277.760 634.230 1280.480 ;
        RECT 638.130 1277.760 653.550 1289.520 ;
        RECT 657.450 1285.235 743.170 1289.520 ;
        RECT 657.450 1277.760 724.570 1285.235 ;
        RECT 387.070 1267.715 724.570 1277.760 ;
        RECT 387.070 1184.500 544.570 1267.715 ;
        RECT 548.470 1184.500 563.170 1267.715 ;
        RECT 567.070 1229.260 724.570 1267.715 ;
        RECT 728.470 1229.260 743.170 1285.235 ;
        RECT 747.070 1289.120 786.030 1294.340 ;
        RECT 789.930 1295.360 805.350 1368.800 ;
        RECT 789.930 1289.120 793.390 1295.360 ;
        RECT 747.070 1280.480 793.390 1289.120 ;
        RECT 800.970 1289.120 805.350 1295.360 ;
        RECT 809.250 1289.120 904.570 1368.800 ;
        RECT 800.970 1280.480 904.570 1289.120 ;
        RECT 747.070 1229.260 904.570 1280.480 ;
        RECT 567.070 1200.160 904.570 1229.260 ;
        RECT 567.070 1184.500 612.150 1200.160 ;
        RECT 387.070 1180.565 612.150 1184.500 ;
        RECT 271.970 1125.340 612.150 1180.565 ;
        RECT 271.970 1109.120 544.570 1125.340 ;
        RECT 207.070 1079.395 544.570 1109.120 ;
        RECT 207.070 1044.420 364.570 1079.395 ;
        RECT 67.075 1042.400 364.570 1044.420 ;
        RECT 67.075 981.280 301.190 1042.400 ;
        RECT 305.090 981.280 364.570 1042.400 ;
        RECT 67.075 955.340 364.570 981.280 ;
        RECT 67.075 870.500 184.570 955.340 ;
        RECT 188.470 870.500 203.170 955.340 ;
        RECT 67.075 852.000 203.170 870.500 ;
        RECT 67.075 796.320 106.150 852.000 ;
        RECT 113.730 811.340 203.170 852.000 ;
        RECT 113.730 796.320 184.570 811.340 ;
        RECT 67.075 730.420 184.570 796.320 ;
        RECT 188.470 730.420 203.170 811.340 ;
        RECT 207.070 881.920 364.570 955.340 ;
        RECT 207.070 799.040 268.070 881.920 ;
        RECT 271.970 866.565 364.570 881.920 ;
        RECT 368.470 866.565 383.170 1079.395 ;
        RECT 387.070 1074.340 544.570 1079.395 ;
        RECT 548.470 1074.340 563.170 1125.340 ;
        RECT 567.070 1109.120 612.150 1125.340 ;
        RECT 616.050 1109.120 631.470 1200.160 ;
        RECT 635.370 1109.120 904.570 1200.160 ;
        RECT 567.070 1091.360 904.570 1109.120 ;
        RECT 567.070 1079.200 611.230 1091.360 ;
        RECT 615.130 1079.600 630.550 1091.360 ;
        RECT 634.450 1079.600 904.570 1091.360 ;
        RECT 617.890 1079.200 630.550 1079.600 ;
        RECT 637.210 1079.395 904.570 1079.600 ;
        RECT 567.070 1074.340 613.990 1079.200 ;
        RECT 387.070 1065.600 613.990 1074.340 ;
        RECT 617.890 1065.600 633.310 1079.200 ;
        RECT 637.210 1065.600 724.570 1079.395 ;
        RECT 387.070 1056.000 724.570 1065.600 ;
        RECT 387.070 964.960 465.870 1056.000 ;
        RECT 469.770 964.960 485.190 1056.000 ;
        RECT 489.090 964.960 636.070 1056.000 ;
        RECT 639.970 964.960 655.390 1056.000 ;
        RECT 659.290 1039.500 724.570 1056.000 ;
        RECT 728.470 1039.500 743.170 1079.395 ;
        RECT 747.070 1056.000 904.570 1079.395 ;
        RECT 747.070 1039.500 786.030 1056.000 ;
        RECT 659.290 980.340 786.030 1039.500 ;
        RECT 659.290 971.235 743.170 980.340 ;
        RECT 659.290 964.960 724.570 971.235 ;
        RECT 387.070 953.715 724.570 964.960 ;
        RECT 387.070 870.500 544.570 953.715 ;
        RECT 548.470 870.500 563.170 953.715 ;
        RECT 567.070 915.260 724.570 953.715 ;
        RECT 728.470 915.260 743.170 971.235 ;
        RECT 747.070 964.960 786.030 980.340 ;
        RECT 789.930 964.960 805.350 1056.000 ;
        RECT 809.250 964.960 904.570 1056.000 ;
        RECT 747.070 915.260 904.570 964.960 ;
        RECT 567.070 887.360 904.570 915.260 ;
        RECT 567.070 875.200 611.230 887.360 ;
        RECT 615.130 875.600 630.550 887.360 ;
        RECT 634.450 875.600 904.570 887.360 ;
        RECT 616.050 875.200 630.550 875.600 ;
        RECT 567.070 870.500 612.150 875.200 ;
        RECT 387.070 866.565 612.150 870.500 ;
        RECT 271.970 811.340 612.150 866.565 ;
        RECT 271.970 799.040 544.570 811.340 ;
        RECT 207.070 765.395 544.570 799.040 ;
        RECT 207.070 730.420 364.570 765.395 ;
        RECT 67.075 641.340 364.570 730.420 ;
        RECT 67.075 589.500 184.570 641.340 ;
        RECT 188.470 589.500 203.170 641.340 ;
        RECT 67.075 536.480 203.170 589.500 ;
        RECT 67.075 516.160 106.150 536.480 ;
        RECT 113.730 530.340 203.170 536.480 ;
        RECT 113.730 516.160 184.570 530.340 ;
        RECT 67.075 416.420 184.570 516.160 ;
        RECT 188.470 416.420 203.170 530.340 ;
        RECT 207.070 604.480 364.570 641.340 ;
        RECT 207.070 516.160 268.070 604.480 ;
        RECT 271.970 552.565 364.570 604.480 ;
        RECT 368.470 552.565 383.170 765.395 ;
        RECT 387.070 760.340 544.570 765.395 ;
        RECT 548.470 760.340 563.170 811.340 ;
        RECT 567.070 796.320 612.150 811.340 ;
        RECT 616.050 796.320 631.470 875.200 ;
        RECT 635.370 796.320 904.570 875.600 ;
        RECT 567.070 775.840 904.570 796.320 ;
        RECT 567.070 760.340 613.990 775.840 ;
        RECT 387.070 750.080 613.990 760.340 ;
        RECT 617.890 750.080 633.310 775.840 ;
        RECT 637.210 765.395 904.570 775.840 ;
        RECT 637.210 750.080 724.570 765.395 ;
        RECT 387.070 740.480 724.570 750.080 ;
        RECT 387.070 652.160 465.870 740.480 ;
        RECT 469.770 652.160 485.190 740.480 ;
        RECT 489.090 652.160 636.070 740.480 ;
        RECT 639.970 652.160 655.390 740.480 ;
        RECT 659.290 725.500 724.570 740.480 ;
        RECT 728.470 725.500 743.170 765.395 ;
        RECT 747.070 740.480 904.570 765.395 ;
        RECT 747.070 725.500 786.030 740.480 ;
        RECT 659.290 666.340 786.030 725.500 ;
        RECT 659.290 657.235 743.170 666.340 ;
        RECT 659.290 652.160 724.570 657.235 ;
        RECT 387.070 639.715 724.570 652.160 ;
        RECT 387.070 589.500 544.570 639.715 ;
        RECT 548.470 589.500 563.170 639.715 ;
        RECT 567.070 604.480 724.570 639.715 ;
        RECT 567.070 589.500 612.150 604.480 ;
        RECT 387.070 552.565 612.150 589.500 ;
        RECT 271.970 530.340 612.150 552.565 ;
        RECT 271.970 516.160 544.570 530.340 ;
        RECT 207.070 451.395 544.570 516.160 ;
        RECT 207.070 416.420 364.570 451.395 ;
        RECT 67.075 327.340 364.570 416.420 ;
        RECT 67.075 14.640 184.570 327.340 ;
        RECT 188.470 14.640 203.170 327.340 ;
        RECT 207.070 242.720 364.570 327.340 ;
        RECT 207.070 181.600 331.550 242.720 ;
        RECT 335.450 181.600 364.570 242.720 ;
        RECT 207.070 14.640 364.570 181.600 ;
        RECT 368.470 14.640 383.170 451.395 ;
        RECT 387.070 446.340 544.570 451.395 ;
        RECT 548.470 446.340 563.170 530.340 ;
        RECT 567.070 516.160 612.150 530.340 ;
        RECT 616.050 516.160 631.470 604.480 ;
        RECT 635.370 601.260 724.570 604.480 ;
        RECT 728.470 601.260 743.170 657.235 ;
        RECT 747.070 652.160 786.030 666.340 ;
        RECT 789.930 652.160 805.350 740.480 ;
        RECT 809.250 652.160 904.570 740.480 ;
        RECT 747.070 601.260 904.570 652.160 ;
        RECT 635.370 516.160 904.570 601.260 ;
        RECT 567.070 463.040 904.570 516.160 ;
        RECT 567.070 446.340 613.990 463.040 ;
        RECT 387.070 437.280 613.990 446.340 ;
        RECT 617.890 437.280 633.310 463.040 ;
        RECT 637.210 451.395 904.570 463.040 ;
        RECT 637.210 437.280 724.570 451.395 ;
        RECT 387.070 427.680 724.570 437.280 ;
        RECT 387.070 414.080 636.070 427.680 ;
        RECT 387.070 325.760 465.870 414.080 ;
        RECT 469.770 325.760 485.190 414.080 ;
        RECT 489.090 336.640 636.070 414.080 ;
        RECT 639.970 336.640 655.390 427.680 ;
        RECT 659.290 411.500 724.570 427.680 ;
        RECT 728.470 411.500 743.170 451.395 ;
        RECT 747.070 427.680 904.570 451.395 ;
        RECT 747.070 411.500 786.030 427.680 ;
        RECT 659.290 352.340 786.030 411.500 ;
        RECT 659.290 343.235 743.170 352.340 ;
        RECT 659.290 336.640 724.570 343.235 ;
        RECT 489.090 325.760 724.570 336.640 ;
        RECT 387.070 325.715 724.570 325.760 ;
        RECT 387.070 277.580 544.570 325.715 ;
        RECT 548.470 277.580 563.170 325.715 ;
        RECT 567.070 277.580 724.570 325.715 ;
        RECT 387.070 253.600 724.570 277.580 ;
        RECT 387.070 165.280 465.870 253.600 ;
        RECT 469.770 165.280 485.190 253.600 ;
        RECT 489.090 180.340 636.070 253.600 ;
        RECT 489.090 165.280 544.570 180.340 ;
        RECT 387.070 14.640 544.570 165.280 ;
        RECT 548.470 14.640 563.170 180.340 ;
        RECT 567.070 165.280 636.070 180.340 ;
        RECT 639.970 165.280 655.390 253.600 ;
        RECT 659.290 239.500 724.570 253.600 ;
        RECT 728.470 239.500 743.170 343.235 ;
        RECT 747.070 336.640 786.030 352.340 ;
        RECT 789.930 336.640 805.350 427.680 ;
        RECT 809.250 336.640 904.570 427.680 ;
        RECT 747.070 253.600 904.570 336.640 ;
        RECT 747.070 239.500 786.030 253.600 ;
        RECT 659.290 180.340 786.030 239.500 ;
        RECT 659.290 165.280 724.570 180.340 ;
        RECT 567.070 14.640 724.570 165.280 ;
        RECT 728.470 63.500 743.170 180.340 ;
        RECT 747.070 165.280 786.030 180.340 ;
        RECT 789.930 165.280 805.350 253.600 ;
        RECT 809.250 165.280 904.570 253.600 ;
        RECT 747.070 63.500 904.570 165.280 ;
        RECT 728.470 14.640 904.570 63.500 ;
        RECT 908.470 14.640 923.170 3488.760 ;
        RECT 927.070 3378.880 1084.570 3488.760 ;
        RECT 927.070 3366.720 941.510 3378.880 ;
        RECT 945.410 3378.565 1084.570 3378.880 ;
        RECT 1088.470 3378.565 1103.170 3488.760 ;
        RECT 1107.070 3378.565 1264.570 3488.760 ;
        RECT 945.410 3366.720 1264.570 3378.565 ;
        RECT 927.070 3362.560 1264.570 3366.720 ;
        RECT 927.070 3350.400 941.510 3362.560 ;
        RECT 945.410 3350.400 1264.570 3362.560 ;
        RECT 927.070 3346.240 1264.570 3350.400 ;
        RECT 927.070 3334.080 941.510 3346.240 ;
        RECT 945.410 3334.080 1264.570 3346.240 ;
        RECT 927.070 3277.395 1264.570 3334.080 ;
        RECT 927.070 3253.760 1084.570 3277.395 ;
        RECT 927.070 3165.440 965.430 3253.760 ;
        RECT 969.330 3237.500 1084.570 3253.760 ;
        RECT 1088.470 3237.500 1103.170 3277.395 ;
        RECT 969.330 3178.340 1103.170 3237.500 ;
        RECT 969.330 3165.440 1084.570 3178.340 ;
        RECT 927.070 3068.800 1084.570 3165.440 ;
        RECT 927.070 3056.640 941.510 3068.800 ;
        RECT 945.410 3064.565 1084.570 3068.800 ;
        RECT 1088.470 3064.565 1103.170 3178.340 ;
        RECT 1107.070 3253.760 1264.570 3277.395 ;
        RECT 1107.070 3240.160 1115.390 3253.760 ;
        RECT 1107.070 3173.600 1107.110 3240.160 ;
        RECT 1111.010 3236.160 1115.390 3240.160 ;
        RECT 1119.290 3240.160 1264.570 3253.760 ;
        RECT 1119.290 3236.160 1126.430 3240.160 ;
        RECT 1111.010 3232.000 1126.430 3236.160 ;
        RECT 1111.010 3219.840 1115.390 3232.000 ;
        RECT 1119.290 3219.840 1126.430 3232.000 ;
        RECT 1111.010 3215.680 1126.430 3219.840 ;
        RECT 1111.010 3203.520 1115.390 3215.680 ;
        RECT 1119.290 3203.520 1126.430 3215.680 ;
        RECT 1111.010 3199.360 1126.430 3203.520 ;
        RECT 1111.010 3187.200 1115.390 3199.360 ;
        RECT 1119.290 3187.200 1126.430 3199.360 ;
        RECT 1111.010 3183.040 1126.430 3187.200 ;
        RECT 1111.010 3173.600 1115.390 3183.040 ;
        RECT 1107.070 3165.440 1115.390 3173.600 ;
        RECT 1119.290 3173.600 1126.430 3183.040 ;
        RECT 1130.330 3173.600 1264.570 3240.160 ;
        RECT 1119.290 3165.440 1264.570 3173.600 ;
        RECT 1107.070 3064.565 1264.570 3165.440 ;
        RECT 945.410 3056.640 1264.570 3064.565 ;
        RECT 927.070 3052.480 1264.570 3056.640 ;
        RECT 927.070 3040.320 941.510 3052.480 ;
        RECT 945.410 3040.320 1264.570 3052.480 ;
        RECT 927.070 3036.160 1264.570 3040.320 ;
        RECT 927.070 3024.000 941.510 3036.160 ;
        RECT 945.410 3024.000 1264.570 3036.160 ;
        RECT 927.070 3019.840 1264.570 3024.000 ;
        RECT 927.070 3007.680 941.510 3019.840 ;
        RECT 945.410 3007.680 1264.570 3019.840 ;
        RECT 927.070 2970.880 1264.570 3007.680 ;
        RECT 927.070 2953.280 943.350 2970.880 ;
        RECT 947.250 2963.395 1264.570 2970.880 ;
        RECT 947.250 2953.280 1084.570 2963.395 ;
        RECT 927.070 2932.800 1084.570 2953.280 ;
        RECT 927.070 2844.480 965.430 2932.800 ;
        RECT 969.330 2917.500 1084.570 2932.800 ;
        RECT 1088.470 2917.500 1103.170 2963.395 ;
        RECT 969.330 2858.340 1103.170 2917.500 ;
        RECT 969.330 2844.480 1084.570 2858.340 ;
        RECT 927.070 2750.565 1084.570 2844.480 ;
        RECT 1088.470 2750.565 1103.170 2858.340 ;
        RECT 1107.070 2932.800 1264.570 2963.395 ;
        RECT 1107.070 2844.480 1115.390 2932.800 ;
        RECT 1119.290 2844.480 1264.570 2932.800 ;
        RECT 1107.070 2750.565 1264.570 2844.480 ;
        RECT 927.070 2742.400 1264.570 2750.565 ;
        RECT 927.070 2730.240 941.510 2742.400 ;
        RECT 945.410 2730.240 1264.570 2742.400 ;
        RECT 927.070 2726.080 1264.570 2730.240 ;
        RECT 927.070 2713.920 941.510 2726.080 ;
        RECT 945.410 2713.920 1264.570 2726.080 ;
        RECT 927.070 2709.760 1264.570 2713.920 ;
        RECT 927.070 2697.600 941.510 2709.760 ;
        RECT 945.410 2697.600 1264.570 2709.760 ;
        RECT 927.070 2660.800 1264.570 2697.600 ;
        RECT 927.070 2637.760 943.350 2660.800 ;
        RECT 947.250 2649.395 1264.570 2660.800 ;
        RECT 947.250 2637.760 1084.570 2649.395 ;
        RECT 927.070 2622.720 1084.570 2637.760 ;
        RECT 927.070 2534.400 965.430 2622.720 ;
        RECT 969.330 2609.500 1084.570 2622.720 ;
        RECT 1088.470 2609.500 1103.170 2649.395 ;
        RECT 969.330 2550.340 1103.170 2609.500 ;
        RECT 969.330 2534.400 1084.570 2550.340 ;
        RECT 927.070 2436.565 1084.570 2534.400 ;
        RECT 1088.470 2436.565 1103.170 2550.340 ;
        RECT 1107.070 2622.720 1264.570 2649.395 ;
        RECT 1107.070 2534.400 1115.390 2622.720 ;
        RECT 1119.290 2534.400 1264.570 2622.720 ;
        RECT 1107.070 2436.565 1264.570 2534.400 ;
        RECT 927.070 2432.320 1264.570 2436.565 ;
        RECT 927.070 2420.160 941.510 2432.320 ;
        RECT 945.410 2420.160 1264.570 2432.320 ;
        RECT 927.070 2416.000 1264.570 2420.160 ;
        RECT 927.070 2403.840 941.510 2416.000 ;
        RECT 945.410 2403.840 1264.570 2416.000 ;
        RECT 927.070 2399.680 1264.570 2403.840 ;
        RECT 927.070 2387.520 941.510 2399.680 ;
        RECT 945.410 2387.520 1264.570 2399.680 ;
        RECT 927.070 2345.280 1264.570 2387.520 ;
        RECT 927.070 2322.240 943.350 2345.280 ;
        RECT 947.250 2335.395 1264.570 2345.280 ;
        RECT 947.250 2322.240 1084.570 2335.395 ;
        RECT 927.070 2307.200 1084.570 2322.240 ;
        RECT 927.070 2224.320 965.430 2307.200 ;
        RECT 969.330 2295.500 1084.570 2307.200 ;
        RECT 1088.470 2295.500 1103.170 2335.395 ;
        RECT 969.330 2236.340 1103.170 2295.500 ;
        RECT 969.330 2224.320 1084.570 2236.340 ;
        RECT 927.070 2122.565 1084.570 2224.320 ;
        RECT 1088.470 2122.565 1103.170 2236.340 ;
        RECT 1107.070 2307.200 1264.570 2335.395 ;
        RECT 1107.070 2224.320 1115.390 2307.200 ;
        RECT 1119.290 2224.320 1264.570 2307.200 ;
        RECT 1107.070 2122.565 1264.570 2224.320 ;
        RECT 927.070 2122.240 1264.570 2122.565 ;
        RECT 927.070 2110.080 941.510 2122.240 ;
        RECT 945.410 2110.080 1264.570 2122.240 ;
        RECT 927.070 2105.920 1264.570 2110.080 ;
        RECT 927.070 2093.760 941.510 2105.920 ;
        RECT 945.410 2093.760 1264.570 2105.920 ;
        RECT 927.070 2089.600 1264.570 2093.760 ;
        RECT 927.070 2077.440 941.510 2089.600 ;
        RECT 945.410 2077.440 1264.570 2089.600 ;
        RECT 927.070 2029.760 1264.570 2077.440 ;
        RECT 927.070 2006.720 943.350 2029.760 ;
        RECT 947.250 2021.395 1264.570 2029.760 ;
        RECT 947.250 2006.720 1084.570 2021.395 ;
        RECT 927.070 1997.120 1084.570 2006.720 ;
        RECT 927.070 1908.800 965.430 1997.120 ;
        RECT 969.330 1981.500 1084.570 1997.120 ;
        RECT 1088.470 1981.500 1103.170 2021.395 ;
        RECT 969.330 1922.340 1103.170 1981.500 ;
        RECT 969.330 1908.800 1084.570 1922.340 ;
        RECT 927.070 1812.160 1084.570 1908.800 ;
        RECT 927.070 1800.000 941.510 1812.160 ;
        RECT 945.410 1808.565 1084.570 1812.160 ;
        RECT 1088.470 1808.565 1103.170 1922.340 ;
        RECT 1107.070 1997.120 1264.570 2021.395 ;
        RECT 1107.070 1983.520 1115.390 1997.120 ;
        RECT 1107.070 1916.960 1107.110 1983.520 ;
        RECT 1111.010 1916.960 1115.390 1983.520 ;
        RECT 1107.070 1908.800 1115.390 1916.960 ;
        RECT 1119.290 1983.520 1264.570 1997.120 ;
        RECT 1119.290 1916.960 1126.430 1983.520 ;
        RECT 1130.330 1916.960 1264.570 1983.520 ;
        RECT 1119.290 1908.800 1264.570 1916.960 ;
        RECT 1107.070 1808.565 1264.570 1908.800 ;
        RECT 945.410 1800.000 1264.570 1808.565 ;
        RECT 927.070 1795.840 1264.570 1800.000 ;
        RECT 927.070 1783.680 941.510 1795.840 ;
        RECT 945.410 1783.680 1264.570 1795.840 ;
        RECT 927.070 1779.520 1264.570 1783.680 ;
        RECT 927.070 1767.360 941.510 1779.520 ;
        RECT 945.410 1767.360 1264.570 1779.520 ;
        RECT 927.070 1763.200 1264.570 1767.360 ;
        RECT 927.070 1751.040 941.510 1763.200 ;
        RECT 945.410 1751.040 1264.570 1763.200 ;
        RECT 927.070 1714.240 1264.570 1751.040 ;
        RECT 927.070 1696.640 943.350 1714.240 ;
        RECT 947.250 1707.395 1264.570 1714.240 ;
        RECT 947.250 1696.640 1084.570 1707.395 ;
        RECT 927.070 1681.600 1084.570 1696.640 ;
        RECT 927.070 1593.280 965.430 1681.600 ;
        RECT 969.330 1667.500 1084.570 1681.600 ;
        RECT 1088.470 1667.500 1103.170 1707.395 ;
        RECT 969.330 1608.340 1103.170 1667.500 ;
        RECT 969.330 1593.280 1084.570 1608.340 ;
        RECT 927.070 1494.565 1084.570 1593.280 ;
        RECT 1088.470 1494.565 1103.170 1608.340 ;
        RECT 1107.070 1681.600 1264.570 1707.395 ;
        RECT 1107.070 1593.280 1115.390 1681.600 ;
        RECT 1119.290 1593.280 1264.570 1681.600 ;
        RECT 1107.070 1494.565 1264.570 1593.280 ;
        RECT 927.070 1485.760 1264.570 1494.565 ;
        RECT 927.070 1473.600 941.510 1485.760 ;
        RECT 945.410 1473.600 1264.570 1485.760 ;
        RECT 927.070 1469.440 1264.570 1473.600 ;
        RECT 927.070 1457.280 941.510 1469.440 ;
        RECT 945.410 1457.280 1264.570 1469.440 ;
        RECT 927.070 1453.120 1264.570 1457.280 ;
        RECT 927.070 1440.960 941.510 1453.120 ;
        RECT 945.410 1440.960 1264.570 1453.120 ;
        RECT 927.070 1404.160 1264.570 1440.960 ;
        RECT 927.070 1381.120 943.350 1404.160 ;
        RECT 947.250 1393.395 1264.570 1404.160 ;
        RECT 947.250 1381.120 1084.570 1393.395 ;
        RECT 927.070 1366.080 1084.570 1381.120 ;
        RECT 927.070 1288.640 965.430 1366.080 ;
        RECT 969.330 1353.500 1084.570 1366.080 ;
        RECT 1088.470 1353.500 1103.170 1393.395 ;
        RECT 969.330 1294.340 1103.170 1353.500 ;
        RECT 969.330 1289.920 1084.570 1294.340 ;
        RECT 969.330 1288.640 1017.870 1289.920 ;
        RECT 927.070 1277.760 1017.870 1288.640 ;
        RECT 1021.770 1277.760 1084.570 1289.920 ;
        RECT 927.070 1181.120 1084.570 1277.760 ;
        RECT 927.070 1130.880 941.510 1181.120 ;
        RECT 945.410 1180.565 1084.570 1181.120 ;
        RECT 1088.470 1180.565 1103.170 1294.340 ;
        RECT 1107.070 1366.080 1264.570 1393.395 ;
        RECT 1107.070 1295.360 1115.390 1366.080 ;
        RECT 1107.070 1283.200 1109.870 1295.360 ;
        RECT 1113.770 1289.120 1115.390 1295.360 ;
        RECT 1119.290 1289.120 1264.570 1366.080 ;
        RECT 1113.770 1283.200 1264.570 1289.120 ;
        RECT 1107.070 1180.565 1264.570 1283.200 ;
        RECT 945.410 1130.880 1264.570 1180.565 ;
        RECT 927.070 1088.640 1264.570 1130.880 ;
        RECT 927.070 1065.600 943.350 1088.640 ;
        RECT 947.250 1079.395 1264.570 1088.640 ;
        RECT 947.250 1065.600 1084.570 1079.395 ;
        RECT 927.070 1056.000 1084.570 1065.600 ;
        RECT 927.070 967.680 965.430 1056.000 ;
        RECT 969.330 1039.500 1084.570 1056.000 ;
        RECT 1088.470 1039.500 1103.170 1079.395 ;
        RECT 969.330 980.340 1103.170 1039.500 ;
        RECT 969.330 967.680 1084.570 980.340 ;
        RECT 927.070 871.040 1084.570 967.680 ;
        RECT 927.070 809.920 941.510 871.040 ;
        RECT 945.410 866.565 1084.570 871.040 ;
        RECT 1088.470 866.565 1103.170 980.340 ;
        RECT 1107.070 1056.000 1264.570 1079.395 ;
        RECT 1107.070 1042.400 1115.390 1056.000 ;
        RECT 1107.070 975.840 1107.110 1042.400 ;
        RECT 1111.010 975.840 1115.390 1042.400 ;
        RECT 1107.070 967.680 1115.390 975.840 ;
        RECT 1119.290 1042.400 1264.570 1056.000 ;
        RECT 1119.290 975.840 1126.430 1042.400 ;
        RECT 1130.330 975.840 1264.570 1042.400 ;
        RECT 1119.290 967.680 1264.570 975.840 ;
        RECT 1107.070 866.565 1264.570 967.680 ;
        RECT 945.410 809.920 1264.570 866.565 ;
        RECT 927.070 773.120 1264.570 809.920 ;
        RECT 927.070 750.080 943.350 773.120 ;
        RECT 947.250 765.395 1264.570 773.120 ;
        RECT 947.250 750.080 1084.570 765.395 ;
        RECT 927.070 740.480 1084.570 750.080 ;
        RECT 927.070 652.160 965.430 740.480 ;
        RECT 969.330 725.500 1084.570 740.480 ;
        RECT 1088.470 725.500 1103.170 765.395 ;
        RECT 969.330 666.340 1103.170 725.500 ;
        RECT 969.330 652.160 1084.570 666.340 ;
        RECT 927.070 577.280 1084.570 652.160 ;
        RECT 927.070 565.120 941.510 577.280 ;
        RECT 945.410 565.120 1084.570 577.280 ;
        RECT 927.070 560.960 1084.570 565.120 ;
        RECT 927.070 548.800 941.510 560.960 ;
        RECT 945.410 552.565 1084.570 560.960 ;
        RECT 1088.470 552.565 1103.170 666.340 ;
        RECT 1107.070 740.480 1264.570 765.395 ;
        RECT 1107.070 652.160 1115.390 740.480 ;
        RECT 1119.290 652.160 1264.570 740.480 ;
        RECT 1107.070 552.565 1264.570 652.160 ;
        RECT 945.410 548.800 1264.570 552.565 ;
        RECT 927.070 544.640 1264.570 548.800 ;
        RECT 927.070 532.480 941.510 544.640 ;
        RECT 945.410 532.480 1264.570 544.640 ;
        RECT 927.070 463.040 1264.570 532.480 ;
        RECT 927.070 440.000 943.350 463.040 ;
        RECT 947.250 451.395 1264.570 463.040 ;
        RECT 947.250 440.000 1084.570 451.395 ;
        RECT 927.070 424.960 1084.570 440.000 ;
        RECT 927.070 336.640 965.430 424.960 ;
        RECT 969.330 411.500 1084.570 424.960 ;
        RECT 1088.470 411.500 1103.170 451.395 ;
        RECT 969.330 352.340 1103.170 411.500 ;
        RECT 969.330 336.640 1084.570 352.340 ;
        RECT 927.070 256.320 1084.570 336.640 ;
        RECT 927.070 244.960 1017.870 256.320 ;
        RECT 927.070 168.000 965.430 244.960 ;
        RECT 969.330 244.160 1017.870 244.960 ;
        RECT 1021.770 244.160 1084.570 256.320 ;
        RECT 969.330 239.500 1084.570 244.160 ;
        RECT 1088.470 239.500 1103.170 352.340 ;
        RECT 969.330 180.340 1103.170 239.500 ;
        RECT 969.330 168.000 1084.570 180.340 ;
        RECT 927.070 14.640 1084.570 168.000 ;
        RECT 1088.470 14.640 1103.170 180.340 ;
        RECT 1107.070 424.960 1264.570 451.395 ;
        RECT 1107.070 336.640 1115.390 424.960 ;
        RECT 1119.290 336.640 1264.570 424.960 ;
        RECT 1107.070 250.880 1264.570 336.640 ;
        RECT 1107.070 242.720 1115.390 250.880 ;
        RECT 1107.070 176.160 1107.110 242.720 ;
        RECT 1111.010 238.720 1115.390 242.720 ;
        RECT 1119.290 242.720 1264.570 250.880 ;
        RECT 1119.290 238.720 1126.430 242.720 ;
        RECT 1111.010 234.560 1126.430 238.720 ;
        RECT 1111.010 216.960 1115.390 234.560 ;
        RECT 1119.290 216.960 1126.430 234.560 ;
        RECT 1111.010 207.360 1126.430 216.960 ;
        RECT 1111.010 189.760 1115.390 207.360 ;
        RECT 1119.290 189.760 1126.430 207.360 ;
        RECT 1111.010 180.160 1126.430 189.760 ;
        RECT 1111.010 176.160 1115.390 180.160 ;
        RECT 1107.070 168.000 1115.390 176.160 ;
        RECT 1119.290 176.160 1126.430 180.160 ;
        RECT 1130.330 176.160 1264.570 242.720 ;
        RECT 1119.290 168.000 1264.570 176.160 ;
        RECT 1107.070 14.640 1264.570 168.000 ;
        RECT 1268.470 14.640 1283.170 3488.760 ;
        RECT 1287.070 3378.565 1444.570 3488.760 ;
        RECT 1448.470 3378.565 1463.170 3488.760 ;
        RECT 1287.070 3277.395 1463.170 3378.565 ;
        RECT 1287.070 3251.040 1444.570 3277.395 ;
        RECT 1287.070 3162.720 1435.550 3251.040 ;
        RECT 1439.450 3162.720 1444.570 3251.040 ;
        RECT 1287.070 3064.565 1444.570 3162.720 ;
        RECT 1448.470 3235.885 1463.170 3277.395 ;
        RECT 1467.070 3441.440 1624.570 3488.760 ;
        RECT 1467.070 3388.480 1570.790 3441.440 ;
        RECT 1574.690 3388.880 1590.110 3441.440 ;
        RECT 1594.010 3388.880 1624.570 3441.440 ;
        RECT 1576.530 3388.480 1590.110 3388.880 ;
        RECT 1467.070 3319.040 1572.630 3388.480 ;
        RECT 1576.530 3319.040 1591.950 3388.480 ;
        RECT 1467.070 3263.360 1570.790 3319.040 ;
        RECT 1576.530 3318.640 1590.110 3319.040 ;
        RECT 1595.850 3318.640 1624.570 3388.880 ;
        RECT 1574.690 3263.360 1590.110 3318.640 ;
        RECT 1594.010 3263.360 1624.570 3318.640 ;
        RECT 1467.070 3235.885 1624.570 3263.360 ;
        RECT 1448.470 3146.275 1624.570 3235.885 ;
        RECT 1448.470 3064.565 1463.170 3146.275 ;
        RECT 1287.070 2963.395 1463.170 3064.565 ;
        RECT 1287.070 2930.080 1444.570 2963.395 ;
        RECT 1287.070 2847.200 1435.550 2930.080 ;
        RECT 1439.450 2847.200 1444.570 2930.080 ;
        RECT 1287.070 2750.565 1444.570 2847.200 ;
        RECT 1448.470 2953.165 1463.170 2963.395 ;
        RECT 1467.070 3128.640 1624.570 3146.275 ;
        RECT 1467.070 3072.960 1570.790 3128.640 ;
        RECT 1574.690 3073.360 1590.110 3128.640 ;
        RECT 1594.010 3073.360 1624.570 3128.640 ;
        RECT 1576.530 3072.960 1590.110 3073.360 ;
        RECT 1467.070 3003.520 1572.630 3072.960 ;
        RECT 1576.530 3003.520 1591.950 3072.960 ;
        RECT 1467.070 2964.160 1570.790 3003.520 ;
        RECT 1576.530 3003.120 1590.110 3003.520 ;
        RECT 1595.850 3003.120 1624.570 3073.360 ;
        RECT 1574.690 2964.560 1590.110 3003.120 ;
        RECT 1594.010 2964.560 1624.570 3003.120 ;
        RECT 1577.450 2964.160 1590.110 2964.560 ;
        RECT 1467.070 2953.165 1573.550 2964.160 ;
        RECT 1448.470 2950.560 1573.550 2953.165 ;
        RECT 1577.450 2950.560 1592.870 2964.160 ;
        RECT 1596.770 2950.560 1624.570 2964.560 ;
        RECT 1448.470 2837.715 1624.570 2950.560 ;
        RECT 1448.470 2750.565 1463.170 2837.715 ;
        RECT 1287.070 2649.395 1463.170 2750.565 ;
        RECT 1287.070 2625.440 1444.570 2649.395 ;
        RECT 1287.070 2537.120 1435.550 2625.440 ;
        RECT 1439.450 2537.120 1444.570 2625.440 ;
        RECT 1287.070 2436.565 1444.570 2537.120 ;
        RECT 1448.470 2639.165 1463.170 2649.395 ;
        RECT 1467.070 2815.840 1624.570 2837.715 ;
        RECT 1467.070 2760.160 1570.790 2815.840 ;
        RECT 1574.690 2760.560 1590.110 2815.840 ;
        RECT 1594.010 2760.560 1624.570 2815.840 ;
        RECT 1576.530 2760.160 1590.110 2760.560 ;
        RECT 1467.070 2690.720 1572.630 2760.160 ;
        RECT 1576.530 2690.720 1591.950 2760.160 ;
        RECT 1467.070 2651.360 1570.790 2690.720 ;
        RECT 1576.530 2690.320 1590.110 2690.720 ;
        RECT 1595.850 2690.320 1624.570 2760.560 ;
        RECT 1574.690 2651.760 1590.110 2690.320 ;
        RECT 1594.010 2651.760 1624.570 2690.320 ;
        RECT 1577.450 2651.360 1590.110 2651.760 ;
        RECT 1467.070 2639.165 1573.550 2651.360 ;
        RECT 1448.470 2635.040 1573.550 2639.165 ;
        RECT 1577.450 2635.040 1592.870 2651.360 ;
        RECT 1596.770 2635.040 1624.570 2651.760 ;
        RECT 1448.470 2523.715 1624.570 2635.040 ;
        RECT 1448.470 2436.565 1463.170 2523.715 ;
        RECT 1287.070 2335.395 1463.170 2436.565 ;
        RECT 1287.070 2309.920 1444.570 2335.395 ;
        RECT 1287.070 2221.600 1435.550 2309.920 ;
        RECT 1439.450 2221.600 1444.570 2309.920 ;
        RECT 1287.070 2122.565 1444.570 2221.600 ;
        RECT 1448.470 2325.165 1463.170 2335.395 ;
        RECT 1467.070 2500.320 1624.570 2523.715 ;
        RECT 1467.070 2447.360 1533.990 2500.320 ;
        RECT 1537.890 2447.360 1553.310 2500.320 ;
        RECT 1557.210 2456.800 1624.570 2500.320 ;
        RECT 1557.210 2447.360 1572.630 2456.800 ;
        RECT 1467.070 2375.200 1572.630 2447.360 ;
        RECT 1576.530 2375.200 1591.950 2456.800 ;
        RECT 1467.070 2335.840 1570.790 2375.200 ;
        RECT 1576.530 2374.800 1590.110 2375.200 ;
        RECT 1595.850 2374.800 1624.570 2456.800 ;
        RECT 1574.690 2336.240 1590.110 2374.800 ;
        RECT 1594.010 2336.240 1624.570 2374.800 ;
        RECT 1577.450 2335.840 1590.110 2336.240 ;
        RECT 1467.070 2325.165 1573.550 2335.840 ;
        RECT 1448.470 2322.240 1573.550 2325.165 ;
        RECT 1577.450 2322.240 1592.870 2335.840 ;
        RECT 1596.770 2322.240 1624.570 2336.240 ;
        RECT 1448.470 2210.030 1624.570 2322.240 ;
        RECT 1448.470 2122.565 1463.170 2210.030 ;
        RECT 1287.070 2021.395 1463.170 2122.565 ;
        RECT 1287.070 1994.400 1444.570 2021.395 ;
        RECT 1287.070 1906.080 1435.550 1994.400 ;
        RECT 1439.450 1906.080 1444.570 1994.400 ;
        RECT 1287.070 1808.565 1444.570 1906.080 ;
        RECT 1448.470 2011.165 1463.170 2021.395 ;
        RECT 1467.070 2187.520 1624.570 2210.030 ;
        RECT 1467.070 2131.840 1570.790 2187.520 ;
        RECT 1574.690 2132.240 1590.110 2187.520 ;
        RECT 1594.010 2132.240 1624.570 2187.520 ;
        RECT 1576.530 2131.840 1590.110 2132.240 ;
        RECT 1467.070 2062.400 1572.630 2131.840 ;
        RECT 1576.530 2062.400 1591.950 2131.840 ;
        RECT 1467.070 2023.040 1570.790 2062.400 ;
        RECT 1576.530 2062.000 1590.110 2062.400 ;
        RECT 1595.850 2062.000 1624.570 2132.240 ;
        RECT 1574.690 2023.440 1590.110 2062.000 ;
        RECT 1594.010 2023.440 1624.570 2062.000 ;
        RECT 1577.450 2023.040 1590.110 2023.440 ;
        RECT 1467.070 2011.165 1573.550 2023.040 ;
        RECT 1448.470 2006.720 1573.550 2011.165 ;
        RECT 1577.450 2006.720 1592.870 2023.040 ;
        RECT 1596.770 2006.720 1624.570 2023.440 ;
        RECT 1448.470 1895.715 1624.570 2006.720 ;
        RECT 1448.470 1808.565 1463.170 1895.715 ;
        RECT 1287.070 1707.395 1463.170 1808.565 ;
        RECT 1287.070 1678.880 1444.570 1707.395 ;
        RECT 1287.070 1596.000 1435.550 1678.880 ;
        RECT 1439.450 1596.000 1444.570 1678.880 ;
        RECT 1287.070 1494.565 1444.570 1596.000 ;
        RECT 1448.470 1697.165 1463.170 1707.395 ;
        RECT 1467.070 1872.000 1624.570 1895.715 ;
        RECT 1467.070 1819.040 1570.790 1872.000 ;
        RECT 1574.690 1819.440 1590.110 1872.000 ;
        RECT 1594.010 1819.440 1624.570 1872.000 ;
        RECT 1576.530 1819.040 1590.110 1819.440 ;
        RECT 1467.070 1746.880 1572.630 1819.040 ;
        RECT 1576.530 1746.880 1591.950 1819.040 ;
        RECT 1467.070 1707.520 1570.790 1746.880 ;
        RECT 1576.530 1746.480 1590.110 1746.880 ;
        RECT 1595.850 1746.480 1624.570 1819.440 ;
        RECT 1574.690 1707.920 1590.110 1746.480 ;
        RECT 1594.010 1707.920 1624.570 1746.480 ;
        RECT 1577.450 1707.520 1590.110 1707.920 ;
        RECT 1467.070 1697.165 1573.550 1707.520 ;
        RECT 1448.470 1693.920 1573.550 1697.165 ;
        RECT 1577.450 1693.920 1592.870 1707.520 ;
        RECT 1596.770 1693.920 1624.570 1707.920 ;
        RECT 1448.470 1581.715 1624.570 1693.920 ;
        RECT 1448.470 1494.565 1463.170 1581.715 ;
        RECT 1287.070 1393.395 1463.170 1494.565 ;
        RECT 1287.070 1368.800 1444.570 1393.395 ;
        RECT 1287.070 1280.480 1435.550 1368.800 ;
        RECT 1439.450 1280.480 1444.570 1368.800 ;
        RECT 1287.070 1180.565 1444.570 1280.480 ;
        RECT 1448.470 1383.165 1463.170 1393.395 ;
        RECT 1467.070 1559.200 1624.570 1581.715 ;
        RECT 1467.070 1503.520 1570.790 1559.200 ;
        RECT 1574.690 1503.920 1590.110 1559.200 ;
        RECT 1594.010 1503.920 1624.570 1559.200 ;
        RECT 1576.530 1503.520 1590.110 1503.920 ;
        RECT 1467.070 1434.080 1572.630 1503.520 ;
        RECT 1576.530 1434.080 1591.950 1503.520 ;
        RECT 1467.070 1394.720 1570.790 1434.080 ;
        RECT 1576.530 1433.680 1590.110 1434.080 ;
        RECT 1595.850 1433.680 1624.570 1503.920 ;
        RECT 1574.690 1395.120 1590.110 1433.680 ;
        RECT 1594.010 1395.120 1624.570 1433.680 ;
        RECT 1577.450 1394.720 1590.110 1395.120 ;
        RECT 1467.070 1383.165 1573.550 1394.720 ;
        RECT 1448.470 1378.400 1573.550 1383.165 ;
        RECT 1577.450 1378.400 1592.870 1394.720 ;
        RECT 1596.770 1378.400 1624.570 1395.120 ;
        RECT 1448.470 1267.715 1624.570 1378.400 ;
        RECT 1448.470 1180.565 1463.170 1267.715 ;
        RECT 1287.070 1079.395 1463.170 1180.565 ;
        RECT 1287.070 1053.280 1444.570 1079.395 ;
        RECT 1287.070 964.960 1435.550 1053.280 ;
        RECT 1439.450 964.960 1444.570 1053.280 ;
        RECT 1287.070 866.565 1444.570 964.960 ;
        RECT 1448.470 1069.165 1463.170 1079.395 ;
        RECT 1467.070 1243.680 1624.570 1267.715 ;
        RECT 1467.070 1190.720 1570.790 1243.680 ;
        RECT 1574.690 1191.120 1590.110 1243.680 ;
        RECT 1594.010 1191.120 1624.570 1243.680 ;
        RECT 1576.530 1190.720 1590.110 1191.120 ;
        RECT 1467.070 1118.560 1572.630 1190.720 ;
        RECT 1576.530 1118.560 1591.950 1190.720 ;
        RECT 1467.070 1079.200 1570.790 1118.560 ;
        RECT 1576.530 1118.160 1590.110 1118.560 ;
        RECT 1595.850 1118.160 1624.570 1191.120 ;
        RECT 1574.690 1079.600 1590.110 1118.160 ;
        RECT 1594.010 1079.600 1624.570 1118.160 ;
        RECT 1577.450 1079.200 1590.110 1079.600 ;
        RECT 1467.070 1069.165 1573.550 1079.200 ;
        RECT 1448.470 1065.600 1573.550 1069.165 ;
        RECT 1577.450 1065.600 1592.870 1079.200 ;
        RECT 1596.770 1065.600 1624.570 1079.600 ;
        RECT 1448.470 953.715 1624.570 1065.600 ;
        RECT 1448.470 866.565 1463.170 953.715 ;
        RECT 1287.070 765.395 1463.170 866.565 ;
        RECT 1287.070 737.760 1444.570 765.395 ;
        RECT 1287.070 654.880 1435.550 737.760 ;
        RECT 1439.450 654.880 1444.570 737.760 ;
        RECT 1287.070 552.565 1444.570 654.880 ;
        RECT 1448.470 755.165 1463.170 765.395 ;
        RECT 1467.070 930.880 1624.570 953.715 ;
        RECT 1467.070 875.200 1570.790 930.880 ;
        RECT 1574.690 875.600 1590.110 930.880 ;
        RECT 1594.010 875.600 1624.570 930.880 ;
        RECT 1576.530 875.200 1590.110 875.600 ;
        RECT 1467.070 805.760 1572.630 875.200 ;
        RECT 1576.530 805.760 1591.950 875.200 ;
        RECT 1467.070 766.400 1570.790 805.760 ;
        RECT 1576.530 805.360 1590.110 805.760 ;
        RECT 1595.850 805.360 1624.570 875.600 ;
        RECT 1574.690 766.800 1590.110 805.360 ;
        RECT 1594.010 766.800 1624.570 805.360 ;
        RECT 1577.450 766.400 1590.110 766.800 ;
        RECT 1467.070 755.165 1573.550 766.400 ;
        RECT 1448.470 750.080 1573.550 755.165 ;
        RECT 1577.450 750.080 1592.870 766.400 ;
        RECT 1596.770 750.080 1624.570 766.800 ;
        RECT 1448.470 639.715 1624.570 750.080 ;
        RECT 1448.470 552.565 1463.170 639.715 ;
        RECT 1287.070 451.395 1463.170 552.565 ;
        RECT 1287.070 427.680 1444.570 451.395 ;
        RECT 1287.070 339.360 1435.550 427.680 ;
        RECT 1439.450 339.360 1444.570 427.680 ;
        RECT 1287.070 253.600 1444.570 339.360 ;
        RECT 1287.070 165.280 1435.550 253.600 ;
        RECT 1439.450 165.280 1444.570 253.600 ;
        RECT 1287.070 14.640 1444.570 165.280 ;
        RECT 1448.470 441.165 1463.170 451.395 ;
        RECT 1467.070 615.360 1624.570 639.715 ;
        RECT 1467.070 595.040 1570.790 615.360 ;
        RECT 1574.690 595.440 1590.110 615.360 ;
        RECT 1594.010 595.440 1624.570 615.360 ;
        RECT 1576.530 595.040 1590.110 595.440 ;
        RECT 1467.070 525.600 1572.630 595.040 ;
        RECT 1576.530 525.600 1591.950 595.040 ;
        RECT 1467.070 453.600 1570.790 525.600 ;
        RECT 1576.530 525.200 1590.110 525.600 ;
        RECT 1595.850 525.200 1624.570 595.440 ;
        RECT 1574.690 454.000 1590.110 525.200 ;
        RECT 1594.010 454.000 1624.570 525.200 ;
        RECT 1577.450 453.600 1590.110 454.000 ;
        RECT 1467.070 441.165 1573.550 453.600 ;
        RECT 1448.470 437.280 1573.550 441.165 ;
        RECT 1577.450 437.280 1592.870 453.600 ;
        RECT 1596.770 437.280 1624.570 454.000 ;
        RECT 1448.470 325.715 1624.570 437.280 ;
        RECT 1448.470 14.640 1463.170 325.715 ;
        RECT 1467.070 14.640 1624.570 325.715 ;
        RECT 1628.470 3378.565 1643.170 3488.760 ;
        RECT 1647.070 3382.500 1804.570 3488.760 ;
        RECT 1808.470 3382.500 1823.170 3488.760 ;
        RECT 1827.070 3397.920 1984.570 3488.760 ;
        RECT 1827.070 3382.500 1891.870 3397.920 ;
        RECT 1647.070 3378.565 1891.870 3382.500 ;
        RECT 1628.470 3323.340 1891.870 3378.565 ;
        RECT 1628.470 3277.395 1804.570 3323.340 ;
        RECT 1628.470 3064.565 1643.170 3277.395 ;
        RECT 1647.070 3253.760 1804.570 3277.395 ;
        RECT 1647.070 3162.720 1746.510 3253.760 ;
        RECT 1750.410 3162.720 1765.830 3253.760 ;
        RECT 1769.730 3235.885 1804.570 3253.760 ;
        RECT 1808.470 3235.885 1823.170 3323.340 ;
        RECT 1827.070 3319.040 1891.870 3323.340 ;
        RECT 1895.770 3319.040 1911.190 3397.920 ;
        RECT 1915.090 3378.565 1984.570 3397.920 ;
        RECT 1988.470 3382.500 2164.570 3488.760 ;
        RECT 2168.470 3382.500 2183.170 3488.760 ;
        RECT 1988.470 3378.565 2183.170 3382.500 ;
        RECT 1915.090 3323.340 2183.170 3378.565 ;
        RECT 1827.070 3306.880 1890.950 3319.040 ;
        RECT 1895.770 3318.640 1910.270 3319.040 ;
        RECT 1915.090 3318.640 2164.570 3323.340 ;
        RECT 1894.850 3306.880 1910.270 3318.640 ;
        RECT 1914.170 3306.880 2164.570 3318.640 ;
        RECT 1827.070 3277.395 2164.570 3306.880 ;
        RECT 1827.070 3253.760 1984.570 3277.395 ;
        RECT 1827.070 3235.885 1916.710 3253.760 ;
        RECT 1769.730 3162.720 1916.710 3235.885 ;
        RECT 1920.610 3162.720 1936.030 3253.760 ;
        RECT 1939.930 3162.720 1984.570 3253.760 ;
        RECT 1647.070 3146.275 1984.570 3162.720 ;
        RECT 1647.070 3068.500 1804.570 3146.275 ;
        RECT 1808.470 3068.500 1823.170 3146.275 ;
        RECT 1827.070 3085.120 1984.570 3146.275 ;
        RECT 1827.070 3072.960 1890.950 3085.120 ;
        RECT 1894.850 3073.360 1910.270 3085.120 ;
        RECT 1914.170 3073.360 1984.570 3085.120 ;
        RECT 1895.770 3072.960 1910.270 3073.360 ;
        RECT 1827.070 3068.500 1891.870 3072.960 ;
        RECT 1647.070 3064.565 1891.870 3068.500 ;
        RECT 1628.470 3009.340 1891.870 3064.565 ;
        RECT 1628.470 2963.395 1804.570 3009.340 ;
        RECT 1628.470 2750.565 1643.170 2963.395 ;
        RECT 1647.070 2953.165 1804.570 2963.395 ;
        RECT 1808.470 2953.165 1823.170 3009.340 ;
        RECT 1827.070 2994.080 1891.870 3009.340 ;
        RECT 1895.770 2994.080 1911.190 3072.960 ;
        RECT 1915.090 3064.565 1984.570 3073.360 ;
        RECT 1988.470 3237.500 2003.170 3277.395 ;
        RECT 2007.070 3253.760 2164.570 3277.395 ;
        RECT 2007.070 3237.500 2066.670 3253.760 ;
        RECT 1988.470 3178.340 2066.670 3237.500 ;
        RECT 1988.470 3113.260 2003.170 3178.340 ;
        RECT 2007.070 3162.720 2066.670 3178.340 ;
        RECT 2070.570 3162.720 2085.990 3253.760 ;
        RECT 2089.890 3250.580 2164.570 3253.760 ;
        RECT 2168.470 3250.580 2183.170 3323.340 ;
        RECT 2089.890 3162.720 2183.170 3250.580 ;
        RECT 2007.070 3146.275 2183.170 3162.720 ;
        RECT 2007.070 3113.260 2164.570 3146.275 ;
        RECT 1988.470 3068.500 2164.570 3113.260 ;
        RECT 2168.470 3068.500 2183.170 3146.275 ;
        RECT 1988.470 3064.565 2183.170 3068.500 ;
        RECT 1915.090 3009.340 2183.170 3064.565 ;
        RECT 1915.090 2994.080 2164.570 3009.340 ;
        RECT 1827.070 2973.600 2164.570 2994.080 ;
        RECT 1827.070 2953.165 1893.710 2973.600 ;
        RECT 1647.070 2950.560 1893.710 2953.165 ;
        RECT 1897.610 2950.560 1913.030 2973.600 ;
        RECT 1916.930 2963.395 2164.570 2973.600 ;
        RECT 1916.930 2950.560 1984.570 2963.395 ;
        RECT 1647.070 2932.800 1984.570 2950.560 ;
        RECT 1647.070 2844.480 1746.510 2932.800 ;
        RECT 1750.410 2844.480 1765.830 2932.800 ;
        RECT 1769.730 2853.920 1916.710 2932.800 ;
        RECT 1920.610 2853.920 1936.030 2932.800 ;
        RECT 1769.730 2844.480 1913.950 2853.920 ;
        RECT 1920.610 2853.520 1933.270 2853.920 ;
        RECT 1939.930 2853.520 1984.570 2932.800 ;
        RECT 1647.070 2841.760 1913.950 2844.480 ;
        RECT 1917.850 2841.760 1933.270 2853.520 ;
        RECT 1937.170 2841.760 1984.570 2853.520 ;
        RECT 1647.070 2837.715 1984.570 2841.760 ;
        RECT 1647.070 2754.500 1804.570 2837.715 ;
        RECT 1808.470 2754.500 1823.170 2837.715 ;
        RECT 1827.070 2769.600 1984.570 2837.715 ;
        RECT 1827.070 2754.500 1891.870 2769.600 ;
        RECT 1647.070 2750.565 1891.870 2754.500 ;
        RECT 1628.470 2695.340 1891.870 2750.565 ;
        RECT 1628.470 2649.395 1804.570 2695.340 ;
        RECT 1628.470 2436.565 1643.170 2649.395 ;
        RECT 1647.070 2639.165 1804.570 2649.395 ;
        RECT 1808.470 2639.165 1823.170 2695.340 ;
        RECT 1827.070 2690.720 1891.870 2695.340 ;
        RECT 1895.770 2690.720 1911.190 2769.600 ;
        RECT 1915.090 2750.565 1984.570 2769.600 ;
        RECT 1988.470 2917.500 2003.170 2963.395 ;
        RECT 2007.070 2958.340 2164.570 2963.395 ;
        RECT 2168.470 2958.340 2183.170 3009.340 ;
        RECT 2007.070 2932.800 2183.170 2958.340 ;
        RECT 2007.070 2917.500 2066.670 2932.800 ;
        RECT 1988.470 2853.120 2066.670 2917.500 ;
        RECT 2070.570 2859.360 2085.990 2932.800 ;
        RECT 2070.570 2853.120 2074.030 2859.360 ;
        RECT 1988.470 2849.235 2074.030 2853.120 ;
        RECT 1988.470 2799.260 2003.170 2849.235 ;
        RECT 2007.070 2844.480 2074.030 2849.235 ;
        RECT 2081.610 2853.120 2085.990 2859.360 ;
        RECT 2089.890 2853.120 2183.170 2932.800 ;
        RECT 2081.610 2844.480 2183.170 2853.120 ;
        RECT 2007.070 2837.715 2183.170 2844.480 ;
        RECT 2007.070 2799.260 2164.570 2837.715 ;
        RECT 1988.470 2754.500 2164.570 2799.260 ;
        RECT 2168.470 2754.500 2183.170 2837.715 ;
        RECT 1988.470 2750.565 2183.170 2754.500 ;
        RECT 1915.090 2695.340 2183.170 2750.565 ;
        RECT 1827.070 2678.560 1890.950 2690.720 ;
        RECT 1895.770 2690.320 1910.270 2690.720 ;
        RECT 1915.090 2690.320 2164.570 2695.340 ;
        RECT 1894.850 2678.560 1910.270 2690.320 ;
        RECT 1914.170 2678.560 2164.570 2690.320 ;
        RECT 1827.070 2660.800 2164.570 2678.560 ;
        RECT 1827.070 2639.165 1893.710 2660.800 ;
        RECT 1647.070 2635.040 1893.710 2639.165 ;
        RECT 1897.610 2635.040 1913.030 2660.800 ;
        RECT 1916.930 2649.395 2164.570 2660.800 ;
        RECT 1916.930 2635.040 1984.570 2649.395 ;
        RECT 1647.070 2625.440 1984.570 2635.040 ;
        RECT 1647.070 2534.400 1746.510 2625.440 ;
        RECT 1750.410 2534.400 1765.830 2625.440 ;
        RECT 1769.730 2534.400 1916.710 2625.440 ;
        RECT 1920.610 2534.400 1936.030 2625.440 ;
        RECT 1939.930 2534.400 1984.570 2625.440 ;
        RECT 1647.070 2523.715 1984.570 2534.400 ;
        RECT 1647.070 2440.500 1804.570 2523.715 ;
        RECT 1808.470 2440.500 1823.170 2523.715 ;
        RECT 1827.070 2456.800 1984.570 2523.715 ;
        RECT 1827.070 2440.500 1891.870 2456.800 ;
        RECT 1647.070 2436.565 1891.870 2440.500 ;
        RECT 1628.470 2381.340 1891.870 2436.565 ;
        RECT 1628.470 2335.395 1804.570 2381.340 ;
        RECT 1628.470 2122.565 1643.170 2335.395 ;
        RECT 1647.070 2325.165 1804.570 2335.395 ;
        RECT 1808.470 2325.165 1823.170 2381.340 ;
        RECT 1827.070 2365.760 1891.870 2381.340 ;
        RECT 1895.770 2365.760 1911.190 2456.800 ;
        RECT 1915.090 2436.565 1984.570 2456.800 ;
        RECT 1988.470 2609.500 2003.170 2649.395 ;
        RECT 2007.070 2644.340 2164.570 2649.395 ;
        RECT 2168.470 2644.340 2183.170 2695.340 ;
        RECT 2007.070 2625.440 2183.170 2644.340 ;
        RECT 2007.070 2609.500 2066.670 2625.440 ;
        RECT 1988.470 2541.235 2066.670 2609.500 ;
        RECT 1988.470 2485.260 2003.170 2541.235 ;
        RECT 2007.070 2534.400 2066.670 2541.235 ;
        RECT 2070.570 2534.400 2085.990 2625.440 ;
        RECT 2089.890 2534.400 2183.170 2625.440 ;
        RECT 2007.070 2523.715 2183.170 2534.400 ;
        RECT 2007.070 2485.260 2164.570 2523.715 ;
        RECT 1988.470 2440.500 2164.570 2485.260 ;
        RECT 2168.470 2440.500 2183.170 2523.715 ;
        RECT 1988.470 2436.565 2183.170 2440.500 ;
        RECT 1915.090 2381.340 2183.170 2436.565 ;
        RECT 1915.090 2365.760 2164.570 2381.340 ;
        RECT 1827.070 2345.280 2164.570 2365.760 ;
        RECT 1827.070 2325.165 1893.710 2345.280 ;
        RECT 1647.070 2322.240 1893.710 2325.165 ;
        RECT 1897.610 2322.240 1913.030 2345.280 ;
        RECT 1916.930 2335.395 2164.570 2345.280 ;
        RECT 1916.930 2322.240 1984.570 2335.395 ;
        RECT 1647.070 2309.920 1984.570 2322.240 ;
        RECT 1647.070 2221.600 1746.510 2309.920 ;
        RECT 1750.410 2221.600 1765.830 2309.920 ;
        RECT 1769.730 2221.600 1916.710 2309.920 ;
        RECT 1920.610 2221.600 1936.030 2309.920 ;
        RECT 1939.930 2221.600 1984.570 2309.920 ;
        RECT 1647.070 2210.030 1984.570 2221.600 ;
        RECT 1647.070 2209.715 1823.170 2210.030 ;
        RECT 1647.070 2126.500 1804.570 2209.715 ;
        RECT 1808.470 2126.500 1823.170 2209.715 ;
        RECT 1827.070 2141.280 1984.570 2210.030 ;
        RECT 1827.070 2126.500 1891.870 2141.280 ;
        RECT 1647.070 2122.565 1891.870 2126.500 ;
        RECT 1628.470 2067.340 1891.870 2122.565 ;
        RECT 1628.470 2021.395 1804.570 2067.340 ;
        RECT 1628.470 1808.565 1643.170 2021.395 ;
        RECT 1647.070 2011.165 1804.570 2021.395 ;
        RECT 1808.470 2011.165 1823.170 2067.340 ;
        RECT 1827.070 2052.960 1891.870 2067.340 ;
        RECT 1895.770 2052.960 1911.190 2141.280 ;
        RECT 1915.090 2122.565 1984.570 2141.280 ;
        RECT 1988.470 2295.500 2003.170 2335.395 ;
        RECT 2007.070 2330.340 2164.570 2335.395 ;
        RECT 2168.470 2330.340 2183.170 2381.340 ;
        RECT 2007.070 2309.920 2183.170 2330.340 ;
        RECT 2007.070 2295.500 2066.670 2309.920 ;
        RECT 1988.470 2227.235 2066.670 2295.500 ;
        RECT 1988.470 2171.260 2003.170 2227.235 ;
        RECT 2007.070 2221.600 2066.670 2227.235 ;
        RECT 2070.570 2221.600 2085.990 2309.920 ;
        RECT 2089.890 2221.600 2183.170 2309.920 ;
        RECT 2007.070 2209.715 2183.170 2221.600 ;
        RECT 2007.070 2171.260 2164.570 2209.715 ;
        RECT 1988.470 2126.500 2164.570 2171.260 ;
        RECT 2168.470 2126.500 2183.170 2209.715 ;
        RECT 1988.470 2122.565 2183.170 2126.500 ;
        RECT 1915.090 2067.340 2183.170 2122.565 ;
        RECT 1915.090 2052.960 2164.570 2067.340 ;
        RECT 1827.070 2032.480 2164.570 2052.960 ;
        RECT 1827.070 2011.165 1893.710 2032.480 ;
        RECT 1647.070 2006.720 1893.710 2011.165 ;
        RECT 1897.610 2006.720 1913.030 2032.480 ;
        RECT 1916.930 2021.395 2164.570 2032.480 ;
        RECT 1916.930 2006.720 1984.570 2021.395 ;
        RECT 1647.070 1997.120 1984.570 2006.720 ;
        RECT 1647.070 1906.080 1746.510 1997.120 ;
        RECT 1750.410 1906.080 1765.830 1997.120 ;
        RECT 1769.730 1906.080 1916.710 1997.120 ;
        RECT 1920.610 1906.080 1936.030 1997.120 ;
        RECT 1939.930 1906.080 1984.570 1997.120 ;
        RECT 1647.070 1895.715 1984.570 1906.080 ;
        RECT 1647.070 1812.500 1804.570 1895.715 ;
        RECT 1808.470 1812.500 1823.170 1895.715 ;
        RECT 1827.070 1828.480 1984.570 1895.715 ;
        RECT 1827.070 1812.500 1891.870 1828.480 ;
        RECT 1647.070 1808.565 1891.870 1812.500 ;
        RECT 1628.470 1753.340 1891.870 1808.565 ;
        RECT 1628.470 1707.395 1804.570 1753.340 ;
        RECT 1628.470 1494.565 1643.170 1707.395 ;
        RECT 1647.070 1697.165 1804.570 1707.395 ;
        RECT 1808.470 1697.165 1823.170 1753.340 ;
        RECT 1827.070 1737.440 1891.870 1753.340 ;
        RECT 1895.770 1737.440 1911.190 1828.480 ;
        RECT 1915.090 1808.565 1984.570 1828.480 ;
        RECT 1988.470 1981.500 2003.170 2021.395 ;
        RECT 2007.070 2016.340 2164.570 2021.395 ;
        RECT 2168.470 2016.340 2183.170 2067.340 ;
        RECT 2007.070 1997.120 2183.170 2016.340 ;
        RECT 2007.070 1981.500 2066.670 1997.120 ;
        RECT 1988.470 1913.235 2066.670 1981.500 ;
        RECT 1988.470 1857.260 2003.170 1913.235 ;
        RECT 2007.070 1906.080 2066.670 1913.235 ;
        RECT 2070.570 1906.080 2085.990 1997.120 ;
        RECT 2089.890 1906.080 2183.170 1997.120 ;
        RECT 2007.070 1895.715 2183.170 1906.080 ;
        RECT 2007.070 1857.260 2164.570 1895.715 ;
        RECT 1988.470 1812.500 2164.570 1857.260 ;
        RECT 2168.470 1812.500 2183.170 1895.715 ;
        RECT 1988.470 1808.565 2183.170 1812.500 ;
        RECT 1915.090 1753.340 2183.170 1808.565 ;
        RECT 1915.090 1737.440 2164.570 1753.340 ;
        RECT 1827.070 1716.960 2164.570 1737.440 ;
        RECT 1827.070 1697.165 1893.710 1716.960 ;
        RECT 1647.070 1693.920 1893.710 1697.165 ;
        RECT 1897.610 1693.920 1913.030 1716.960 ;
        RECT 1916.930 1707.395 2164.570 1716.960 ;
        RECT 1916.930 1693.920 1984.570 1707.395 ;
        RECT 1647.070 1684.320 1984.570 1693.920 ;
        RECT 1647.070 1681.600 1886.350 1684.320 ;
        RECT 1647.070 1593.280 1746.510 1681.600 ;
        RECT 1750.410 1593.280 1765.830 1681.600 ;
        RECT 1769.730 1672.160 1886.350 1681.600 ;
        RECT 1890.250 1672.160 1905.670 1684.320 ;
        RECT 1909.570 1672.960 1984.570 1684.320 ;
        RECT 1909.570 1672.160 1916.710 1672.960 ;
        RECT 1769.730 1593.280 1916.710 1672.160 ;
        RECT 1920.610 1593.280 1936.030 1672.960 ;
        RECT 1939.930 1593.280 1984.570 1672.960 ;
        RECT 1647.070 1581.715 1984.570 1593.280 ;
        RECT 1647.070 1498.500 1804.570 1581.715 ;
        RECT 1808.470 1498.500 1823.170 1581.715 ;
        RECT 1827.070 1512.960 1984.570 1581.715 ;
        RECT 1827.070 1498.500 1891.870 1512.960 ;
        RECT 1647.070 1494.565 1891.870 1498.500 ;
        RECT 1628.470 1439.340 1891.870 1494.565 ;
        RECT 1628.470 1393.395 1804.570 1439.340 ;
        RECT 1628.470 1180.565 1643.170 1393.395 ;
        RECT 1647.070 1383.165 1804.570 1393.395 ;
        RECT 1808.470 1383.165 1823.170 1439.340 ;
        RECT 1827.070 1424.640 1891.870 1439.340 ;
        RECT 1895.770 1424.640 1911.190 1512.960 ;
        RECT 1915.090 1494.565 1984.570 1512.960 ;
        RECT 1988.470 1667.500 2003.170 1707.395 ;
        RECT 2007.070 1702.340 2164.570 1707.395 ;
        RECT 2168.470 1702.340 2183.170 1753.340 ;
        RECT 2007.070 1681.600 2183.170 1702.340 ;
        RECT 2007.070 1672.960 2074.030 1681.600 ;
        RECT 2007.070 1667.500 2066.670 1672.960 ;
        RECT 1988.470 1599.235 2066.670 1667.500 ;
        RECT 1988.470 1543.260 2003.170 1599.235 ;
        RECT 2007.070 1593.280 2066.670 1599.235 ;
        RECT 2070.570 1666.720 2074.030 1672.960 ;
        RECT 2081.610 1672.960 2183.170 1681.600 ;
        RECT 2081.610 1666.720 2085.990 1672.960 ;
        RECT 2070.570 1593.280 2085.990 1666.720 ;
        RECT 2089.890 1593.280 2183.170 1672.960 ;
        RECT 2007.070 1581.715 2183.170 1593.280 ;
        RECT 2007.070 1543.260 2164.570 1581.715 ;
        RECT 1988.470 1498.500 2164.570 1543.260 ;
        RECT 2168.470 1498.500 2183.170 1581.715 ;
        RECT 1988.470 1494.565 2183.170 1498.500 ;
        RECT 1915.090 1439.340 2183.170 1494.565 ;
        RECT 1915.090 1424.640 2164.570 1439.340 ;
        RECT 1827.070 1404.160 2164.570 1424.640 ;
        RECT 1827.070 1383.165 1893.710 1404.160 ;
        RECT 1647.070 1378.400 1893.710 1383.165 ;
        RECT 1897.610 1378.400 1913.030 1404.160 ;
        RECT 1916.930 1393.395 2164.570 1404.160 ;
        RECT 1916.930 1378.400 1984.570 1393.395 ;
        RECT 1647.070 1368.800 1984.570 1378.400 ;
        RECT 1647.070 1280.480 1746.510 1368.800 ;
        RECT 1750.410 1280.480 1765.830 1368.800 ;
        RECT 1769.730 1280.480 1916.710 1368.800 ;
        RECT 1920.610 1280.480 1936.030 1368.800 ;
        RECT 1939.930 1280.480 1984.570 1368.800 ;
        RECT 1647.070 1267.715 1984.570 1280.480 ;
        RECT 1647.070 1184.500 1804.570 1267.715 ;
        RECT 1808.470 1184.500 1823.170 1267.715 ;
        RECT 1827.070 1200.160 1984.570 1267.715 ;
        RECT 1827.070 1184.500 1891.870 1200.160 ;
        RECT 1647.070 1180.565 1891.870 1184.500 ;
        RECT 1628.470 1125.340 1891.870 1180.565 ;
        RECT 1628.470 1079.395 1804.570 1125.340 ;
        RECT 1628.470 866.565 1643.170 1079.395 ;
        RECT 1647.070 1069.165 1804.570 1079.395 ;
        RECT 1808.470 1069.165 1823.170 1125.340 ;
        RECT 1827.070 1109.120 1891.870 1125.340 ;
        RECT 1895.770 1109.120 1911.190 1200.160 ;
        RECT 1915.090 1180.565 1984.570 1200.160 ;
        RECT 1988.470 1353.500 2003.170 1393.395 ;
        RECT 2007.070 1388.340 2164.570 1393.395 ;
        RECT 2168.470 1388.340 2183.170 1439.340 ;
        RECT 2007.070 1368.800 2183.170 1388.340 ;
        RECT 2007.070 1353.500 2066.670 1368.800 ;
        RECT 1988.470 1285.235 2066.670 1353.500 ;
        RECT 1988.470 1229.260 2003.170 1285.235 ;
        RECT 2007.070 1280.480 2066.670 1285.235 ;
        RECT 2070.570 1280.480 2085.990 1368.800 ;
        RECT 2089.890 1280.480 2183.170 1368.800 ;
        RECT 2007.070 1267.715 2183.170 1280.480 ;
        RECT 2007.070 1229.260 2164.570 1267.715 ;
        RECT 1988.470 1184.500 2164.570 1229.260 ;
        RECT 2168.470 1184.500 2183.170 1267.715 ;
        RECT 1988.470 1180.565 2183.170 1184.500 ;
        RECT 1915.090 1125.340 2183.170 1180.565 ;
        RECT 1915.090 1109.120 2164.570 1125.340 ;
        RECT 1827.070 1091.360 2164.570 1109.120 ;
        RECT 1827.070 1079.200 1890.950 1091.360 ;
        RECT 1894.850 1079.600 1910.270 1091.360 ;
        RECT 1914.170 1079.600 2164.570 1091.360 ;
        RECT 1897.610 1079.200 1910.270 1079.600 ;
        RECT 1916.930 1079.395 2164.570 1079.600 ;
        RECT 1827.070 1069.165 1893.710 1079.200 ;
        RECT 1647.070 1065.600 1893.710 1069.165 ;
        RECT 1897.610 1065.600 1913.030 1079.200 ;
        RECT 1916.930 1065.600 1984.570 1079.395 ;
        RECT 1647.070 1056.000 1984.570 1065.600 ;
        RECT 1647.070 964.960 1746.510 1056.000 ;
        RECT 1750.410 964.960 1765.830 1056.000 ;
        RECT 1769.730 964.960 1916.710 1056.000 ;
        RECT 1920.610 964.960 1936.030 1056.000 ;
        RECT 1939.930 964.960 1984.570 1056.000 ;
        RECT 1647.070 953.715 1984.570 964.960 ;
        RECT 1647.070 870.500 1804.570 953.715 ;
        RECT 1808.470 870.500 1823.170 953.715 ;
        RECT 1827.070 887.360 1984.570 953.715 ;
        RECT 1827.070 875.200 1890.950 887.360 ;
        RECT 1894.850 875.600 1910.270 887.360 ;
        RECT 1914.170 875.600 1984.570 887.360 ;
        RECT 1895.770 875.200 1910.270 875.600 ;
        RECT 1827.070 870.500 1891.870 875.200 ;
        RECT 1647.070 866.565 1891.870 870.500 ;
        RECT 1628.470 811.340 1891.870 866.565 ;
        RECT 1628.470 765.395 1804.570 811.340 ;
        RECT 1628.470 552.565 1643.170 765.395 ;
        RECT 1647.070 755.165 1804.570 765.395 ;
        RECT 1808.470 755.165 1823.170 811.340 ;
        RECT 1827.070 796.320 1891.870 811.340 ;
        RECT 1895.770 796.320 1911.190 875.200 ;
        RECT 1915.090 866.565 1984.570 875.600 ;
        RECT 1988.470 1039.500 2003.170 1079.395 ;
        RECT 2007.070 1074.340 2164.570 1079.395 ;
        RECT 2168.470 1074.340 2183.170 1125.340 ;
        RECT 2007.070 1056.000 2183.170 1074.340 ;
        RECT 2007.070 1039.500 2066.670 1056.000 ;
        RECT 1988.470 971.235 2066.670 1039.500 ;
        RECT 1988.470 915.260 2003.170 971.235 ;
        RECT 2007.070 964.960 2066.670 971.235 ;
        RECT 2070.570 964.960 2085.990 1056.000 ;
        RECT 2089.890 964.960 2183.170 1056.000 ;
        RECT 2007.070 953.715 2183.170 964.960 ;
        RECT 2007.070 915.260 2164.570 953.715 ;
        RECT 1988.470 870.500 2164.570 915.260 ;
        RECT 2168.470 870.500 2183.170 953.715 ;
        RECT 1988.470 866.565 2183.170 870.500 ;
        RECT 1915.090 811.340 2183.170 866.565 ;
        RECT 1915.090 796.320 2164.570 811.340 ;
        RECT 1827.070 775.840 2164.570 796.320 ;
        RECT 1827.070 755.165 1893.710 775.840 ;
        RECT 1647.070 750.080 1893.710 755.165 ;
        RECT 1897.610 750.080 1913.030 775.840 ;
        RECT 1916.930 765.395 2164.570 775.840 ;
        RECT 1916.930 750.080 1984.570 765.395 ;
        RECT 1647.070 740.480 1984.570 750.080 ;
        RECT 1647.070 652.160 1746.510 740.480 ;
        RECT 1750.410 652.160 1765.830 740.480 ;
        RECT 1769.730 652.160 1916.710 740.480 ;
        RECT 1920.610 652.160 1936.030 740.480 ;
        RECT 1939.930 652.160 1984.570 740.480 ;
        RECT 1647.070 639.715 1984.570 652.160 ;
        RECT 1647.070 589.500 1804.570 639.715 ;
        RECT 1808.470 589.500 1823.170 639.715 ;
        RECT 1827.070 604.480 1984.570 639.715 ;
        RECT 1827.070 589.500 1891.870 604.480 ;
        RECT 1647.070 552.565 1891.870 589.500 ;
        RECT 1628.470 530.340 1891.870 552.565 ;
        RECT 1628.470 451.395 1804.570 530.340 ;
        RECT 1628.470 14.640 1643.170 451.395 ;
        RECT 1647.070 441.165 1804.570 451.395 ;
        RECT 1808.470 441.165 1823.170 530.340 ;
        RECT 1827.070 516.160 1891.870 530.340 ;
        RECT 1895.770 516.160 1911.190 604.480 ;
        RECT 1915.090 552.565 1984.570 604.480 ;
        RECT 1988.470 725.500 2003.170 765.395 ;
        RECT 2007.070 760.340 2164.570 765.395 ;
        RECT 2168.470 760.340 2183.170 811.340 ;
        RECT 2007.070 740.480 2183.170 760.340 ;
        RECT 2007.070 725.500 2066.670 740.480 ;
        RECT 1988.470 657.235 2066.670 725.500 ;
        RECT 1988.470 601.260 2003.170 657.235 ;
        RECT 2007.070 652.160 2066.670 657.235 ;
        RECT 2070.570 652.160 2085.990 740.480 ;
        RECT 2089.890 652.160 2183.170 740.480 ;
        RECT 2007.070 639.715 2183.170 652.160 ;
        RECT 2007.070 601.260 2164.570 639.715 ;
        RECT 1988.470 589.500 2164.570 601.260 ;
        RECT 2168.470 589.500 2183.170 639.715 ;
        RECT 1988.470 552.565 2183.170 589.500 ;
        RECT 1915.090 530.340 2183.170 552.565 ;
        RECT 1915.090 516.160 2164.570 530.340 ;
        RECT 1827.070 463.040 2164.570 516.160 ;
        RECT 1827.070 441.165 1893.710 463.040 ;
        RECT 1647.070 437.280 1893.710 441.165 ;
        RECT 1897.610 437.280 1913.030 463.040 ;
        RECT 1916.930 451.395 2164.570 463.040 ;
        RECT 1916.930 437.280 1984.570 451.395 ;
        RECT 1647.070 427.680 1984.570 437.280 ;
        RECT 1647.070 336.640 1746.510 427.680 ;
        RECT 1750.410 336.640 1765.830 427.680 ;
        RECT 1769.730 336.640 1916.710 427.680 ;
        RECT 1920.610 336.640 1936.030 427.680 ;
        RECT 1939.930 336.640 1984.570 427.680 ;
        RECT 1647.070 325.715 1984.570 336.640 ;
        RECT 1647.070 253.600 1804.570 325.715 ;
        RECT 1647.070 165.280 1746.510 253.600 ;
        RECT 1750.410 165.280 1765.830 253.600 ;
        RECT 1769.730 165.280 1804.570 253.600 ;
        RECT 1647.070 14.640 1804.570 165.280 ;
        RECT 1808.470 14.640 1823.170 325.715 ;
        RECT 1827.070 253.600 1984.570 325.715 ;
        RECT 1827.070 165.280 1916.710 253.600 ;
        RECT 1920.610 165.280 1936.030 253.600 ;
        RECT 1939.930 165.280 1984.570 253.600 ;
        RECT 1827.070 14.640 1984.570 165.280 ;
        RECT 1988.470 411.500 2003.170 451.395 ;
        RECT 2007.070 446.340 2164.570 451.395 ;
        RECT 2168.470 446.340 2183.170 530.340 ;
        RECT 2007.070 427.680 2183.170 446.340 ;
        RECT 2007.070 411.500 2066.670 427.680 ;
        RECT 1988.470 343.235 2066.670 411.500 ;
        RECT 1988.470 239.500 2003.170 343.235 ;
        RECT 2007.070 336.640 2066.670 343.235 ;
        RECT 2070.570 336.640 2085.990 427.680 ;
        RECT 2089.890 336.640 2183.170 427.680 ;
        RECT 2007.070 325.715 2183.170 336.640 ;
        RECT 2007.070 277.580 2164.570 325.715 ;
        RECT 2168.470 277.580 2183.170 325.715 ;
        RECT 2007.070 253.600 2183.170 277.580 ;
        RECT 2007.070 239.500 2066.670 253.600 ;
        RECT 1988.470 180.340 2066.670 239.500 ;
        RECT 1988.470 14.640 2003.170 180.340 ;
        RECT 2007.070 165.280 2066.670 180.340 ;
        RECT 2070.570 165.280 2085.990 253.600 ;
        RECT 2089.890 180.340 2183.170 253.600 ;
        RECT 2089.890 165.280 2164.570 180.340 ;
        RECT 2007.070 14.640 2164.570 165.280 ;
        RECT 2168.470 14.640 2183.170 180.340 ;
        RECT 2187.070 3427.260 2344.570 3488.760 ;
        RECT 2348.470 3427.260 2363.170 3488.760 ;
        RECT 2367.070 3427.260 2524.570 3488.760 ;
        RECT 2187.070 3397.920 2524.570 3427.260 ;
        RECT 2187.070 3319.040 2212.030 3397.920 ;
        RECT 2215.930 3319.040 2231.350 3397.920 ;
        RECT 2187.070 3306.880 2211.110 3319.040 ;
        RECT 2215.930 3318.640 2230.430 3319.040 ;
        RECT 2235.250 3318.640 2524.570 3397.920 ;
        RECT 2215.010 3306.880 2230.430 3318.640 ;
        RECT 2234.330 3306.880 2524.570 3318.640 ;
        RECT 2187.070 3277.395 2524.570 3306.880 ;
        RECT 2187.070 3253.760 2344.570 3277.395 ;
        RECT 2187.070 3162.720 2235.950 3253.760 ;
        RECT 2239.850 3162.720 2255.270 3253.760 ;
        RECT 2259.170 3237.500 2344.570 3253.760 ;
        RECT 2348.470 3237.500 2363.170 3277.395 ;
        RECT 2367.070 3253.760 2524.570 3277.395 ;
        RECT 2367.070 3237.500 2385.910 3253.760 ;
        RECT 2259.170 3178.340 2385.910 3237.500 ;
        RECT 2259.170 3162.720 2344.570 3178.340 ;
        RECT 2187.070 3113.260 2344.570 3162.720 ;
        RECT 2348.470 3113.260 2363.170 3178.340 ;
        RECT 2367.070 3162.720 2385.910 3178.340 ;
        RECT 2389.810 3162.720 2405.230 3253.760 ;
        RECT 2409.130 3162.720 2524.570 3253.760 ;
        RECT 2367.070 3113.260 2524.570 3162.720 ;
        RECT 2187.070 3085.120 2524.570 3113.260 ;
        RECT 2187.070 3072.960 2211.110 3085.120 ;
        RECT 2215.010 3073.360 2230.430 3085.120 ;
        RECT 2234.330 3073.360 2524.570 3085.120 ;
        RECT 2215.930 3072.960 2230.430 3073.360 ;
        RECT 2187.070 2994.080 2212.030 3072.960 ;
        RECT 2215.930 2994.080 2231.350 3072.960 ;
        RECT 2235.250 2994.080 2524.570 3073.360 ;
        RECT 2187.070 2973.600 2524.570 2994.080 ;
        RECT 2187.070 2950.560 2213.870 2973.600 ;
        RECT 2217.770 2950.560 2233.190 2973.600 ;
        RECT 2237.090 2963.395 2524.570 2973.600 ;
        RECT 2237.090 2950.560 2344.570 2963.395 ;
        RECT 2187.070 2932.800 2344.570 2950.560 ;
        RECT 2187.070 2844.480 2235.950 2932.800 ;
        RECT 2239.850 2844.480 2255.270 2932.800 ;
        RECT 2259.170 2917.500 2344.570 2932.800 ;
        RECT 2348.470 2917.500 2363.170 2963.395 ;
        RECT 2367.070 2932.800 2524.570 2963.395 ;
        RECT 2367.070 2917.500 2385.910 2932.800 ;
        RECT 2259.170 2858.340 2385.910 2917.500 ;
        RECT 2259.170 2844.480 2344.570 2858.340 ;
        RECT 2187.070 2799.260 2344.570 2844.480 ;
        RECT 2348.470 2799.260 2363.170 2858.340 ;
        RECT 2367.070 2844.480 2385.910 2858.340 ;
        RECT 2389.810 2844.480 2405.230 2932.800 ;
        RECT 2409.130 2844.480 2524.570 2932.800 ;
        RECT 2367.070 2799.260 2524.570 2844.480 ;
        RECT 2187.070 2769.600 2524.570 2799.260 ;
        RECT 2187.070 2681.280 2212.030 2769.600 ;
        RECT 2215.930 2681.280 2231.350 2769.600 ;
        RECT 2235.250 2681.280 2524.570 2769.600 ;
        RECT 2187.070 2660.800 2524.570 2681.280 ;
        RECT 2187.070 2635.040 2213.870 2660.800 ;
        RECT 2217.770 2635.040 2233.190 2660.800 ;
        RECT 2237.090 2649.395 2524.570 2660.800 ;
        RECT 2237.090 2635.040 2344.570 2649.395 ;
        RECT 2187.070 2625.440 2344.570 2635.040 ;
        RECT 2187.070 2534.400 2235.950 2625.440 ;
        RECT 2239.850 2534.400 2255.270 2625.440 ;
        RECT 2259.170 2609.500 2344.570 2625.440 ;
        RECT 2348.470 2609.500 2363.170 2649.395 ;
        RECT 2367.070 2625.440 2524.570 2649.395 ;
        RECT 2367.070 2609.500 2385.910 2625.440 ;
        RECT 2259.170 2550.340 2385.910 2609.500 ;
        RECT 2259.170 2534.400 2344.570 2550.340 ;
        RECT 2187.070 2485.260 2344.570 2534.400 ;
        RECT 2348.470 2485.260 2363.170 2550.340 ;
        RECT 2367.070 2534.400 2385.910 2550.340 ;
        RECT 2389.810 2534.400 2405.230 2625.440 ;
        RECT 2409.130 2534.400 2524.570 2625.440 ;
        RECT 2367.070 2485.260 2524.570 2534.400 ;
        RECT 2187.070 2456.800 2524.570 2485.260 ;
        RECT 2187.070 2365.760 2212.030 2456.800 ;
        RECT 2215.930 2365.760 2231.350 2456.800 ;
        RECT 2235.250 2365.760 2524.570 2456.800 ;
        RECT 2187.070 2345.280 2524.570 2365.760 ;
        RECT 2187.070 2322.240 2213.870 2345.280 ;
        RECT 2217.770 2322.240 2233.190 2345.280 ;
        RECT 2237.090 2335.395 2524.570 2345.280 ;
        RECT 2237.090 2322.240 2344.570 2335.395 ;
        RECT 2187.070 2309.920 2344.570 2322.240 ;
        RECT 2187.070 2221.600 2235.950 2309.920 ;
        RECT 2239.850 2221.600 2255.270 2309.920 ;
        RECT 2259.170 2295.500 2344.570 2309.920 ;
        RECT 2348.470 2295.500 2363.170 2335.395 ;
        RECT 2367.070 2309.920 2524.570 2335.395 ;
        RECT 2367.070 2295.500 2385.910 2309.920 ;
        RECT 2259.170 2236.340 2385.910 2295.500 ;
        RECT 2259.170 2221.600 2344.570 2236.340 ;
        RECT 2187.070 2171.260 2344.570 2221.600 ;
        RECT 2348.470 2171.260 2363.170 2236.340 ;
        RECT 2367.070 2221.600 2385.910 2236.340 ;
        RECT 2389.810 2221.600 2405.230 2309.920 ;
        RECT 2409.130 2221.600 2524.570 2309.920 ;
        RECT 2367.070 2171.260 2524.570 2221.600 ;
        RECT 2187.070 2141.280 2524.570 2171.260 ;
        RECT 2187.070 2052.960 2212.030 2141.280 ;
        RECT 2215.930 2052.960 2231.350 2141.280 ;
        RECT 2235.250 2052.960 2524.570 2141.280 ;
        RECT 2187.070 2032.480 2524.570 2052.960 ;
        RECT 2187.070 2006.720 2213.870 2032.480 ;
        RECT 2217.770 2006.720 2233.190 2032.480 ;
        RECT 2237.090 2021.395 2524.570 2032.480 ;
        RECT 2237.090 2006.720 2344.570 2021.395 ;
        RECT 2187.070 1997.120 2344.570 2006.720 ;
        RECT 2187.070 1906.080 2235.950 1997.120 ;
        RECT 2239.850 1906.080 2255.270 1997.120 ;
        RECT 2259.170 1981.500 2344.570 1997.120 ;
        RECT 2348.470 1981.500 2363.170 2021.395 ;
        RECT 2367.070 1997.120 2524.570 2021.395 ;
        RECT 2367.070 1981.500 2385.910 1997.120 ;
        RECT 2259.170 1922.340 2385.910 1981.500 ;
        RECT 2259.170 1906.080 2344.570 1922.340 ;
        RECT 2187.070 1857.260 2344.570 1906.080 ;
        RECT 2348.470 1857.260 2363.170 1922.340 ;
        RECT 2367.070 1906.080 2385.910 1922.340 ;
        RECT 2389.810 1906.080 2405.230 1997.120 ;
        RECT 2409.130 1906.080 2524.570 1997.120 ;
        RECT 2367.070 1857.260 2524.570 1906.080 ;
        RECT 2187.070 1828.480 2524.570 1857.260 ;
        RECT 2187.070 1737.440 2212.030 1828.480 ;
        RECT 2215.930 1737.440 2231.350 1828.480 ;
        RECT 2235.250 1737.440 2524.570 1828.480 ;
        RECT 2187.070 1716.960 2524.570 1737.440 ;
        RECT 2187.070 1693.920 2213.870 1716.960 ;
        RECT 2217.770 1693.920 2233.190 1716.960 ;
        RECT 2237.090 1707.395 2524.570 1716.960 ;
        RECT 2237.090 1693.920 2344.570 1707.395 ;
        RECT 2187.070 1684.320 2344.570 1693.920 ;
        RECT 2187.070 1672.160 2206.510 1684.320 ;
        RECT 2210.410 1672.160 2225.830 1684.320 ;
        RECT 2229.730 1672.960 2344.570 1684.320 ;
        RECT 2229.730 1672.160 2235.950 1672.960 ;
        RECT 2187.070 1593.280 2235.950 1672.160 ;
        RECT 2239.850 1593.280 2255.270 1672.960 ;
        RECT 2259.170 1667.500 2344.570 1672.960 ;
        RECT 2348.470 1667.500 2363.170 1707.395 ;
        RECT 2367.070 1681.600 2524.570 1707.395 ;
        RECT 2367.070 1672.960 2394.190 1681.600 ;
        RECT 2367.070 1667.500 2385.910 1672.960 ;
        RECT 2259.170 1608.340 2385.910 1667.500 ;
        RECT 2259.170 1593.280 2344.570 1608.340 ;
        RECT 2187.070 1543.260 2344.570 1593.280 ;
        RECT 2348.470 1543.260 2363.170 1608.340 ;
        RECT 2367.070 1593.280 2385.910 1608.340 ;
        RECT 2389.810 1666.720 2394.190 1672.960 ;
        RECT 2401.770 1672.960 2524.570 1681.600 ;
        RECT 2401.770 1666.720 2405.230 1672.960 ;
        RECT 2389.810 1593.280 2405.230 1666.720 ;
        RECT 2409.130 1593.280 2524.570 1672.960 ;
        RECT 2367.070 1543.260 2524.570 1593.280 ;
        RECT 2187.070 1512.960 2524.570 1543.260 ;
        RECT 2187.070 1424.640 2212.030 1512.960 ;
        RECT 2215.930 1424.640 2231.350 1512.960 ;
        RECT 2235.250 1424.640 2524.570 1512.960 ;
        RECT 2187.070 1404.160 2524.570 1424.640 ;
        RECT 2187.070 1378.400 2213.870 1404.160 ;
        RECT 2217.770 1378.400 2233.190 1404.160 ;
        RECT 2237.090 1393.395 2524.570 1404.160 ;
        RECT 2237.090 1378.400 2344.570 1393.395 ;
        RECT 2187.070 1368.800 2344.570 1378.400 ;
        RECT 2187.070 1280.480 2235.950 1368.800 ;
        RECT 2239.850 1280.480 2255.270 1368.800 ;
        RECT 2259.170 1353.500 2344.570 1368.800 ;
        RECT 2348.470 1353.500 2363.170 1393.395 ;
        RECT 2367.070 1368.800 2524.570 1393.395 ;
        RECT 2367.070 1353.500 2385.910 1368.800 ;
        RECT 2259.170 1294.340 2385.910 1353.500 ;
        RECT 2259.170 1280.480 2344.570 1294.340 ;
        RECT 2187.070 1229.260 2344.570 1280.480 ;
        RECT 2348.470 1229.260 2363.170 1294.340 ;
        RECT 2367.070 1280.480 2385.910 1294.340 ;
        RECT 2389.810 1280.480 2405.230 1368.800 ;
        RECT 2409.130 1280.480 2524.570 1368.800 ;
        RECT 2367.070 1229.260 2524.570 1280.480 ;
        RECT 2187.070 1200.160 2524.570 1229.260 ;
        RECT 2187.070 1109.120 2212.030 1200.160 ;
        RECT 2215.930 1109.120 2231.350 1200.160 ;
        RECT 2235.250 1109.120 2524.570 1200.160 ;
        RECT 2187.070 1088.640 2524.570 1109.120 ;
        RECT 2187.070 1065.600 2213.870 1088.640 ;
        RECT 2217.770 1065.600 2233.190 1088.640 ;
        RECT 2237.090 1079.395 2524.570 1088.640 ;
        RECT 2237.090 1065.600 2344.570 1079.395 ;
        RECT 2187.070 1056.000 2344.570 1065.600 ;
        RECT 2187.070 964.960 2235.950 1056.000 ;
        RECT 2239.850 964.960 2255.270 1056.000 ;
        RECT 2259.170 1039.500 2344.570 1056.000 ;
        RECT 2348.470 1039.500 2363.170 1079.395 ;
        RECT 2367.070 1056.000 2524.570 1079.395 ;
        RECT 2367.070 1039.500 2385.910 1056.000 ;
        RECT 2259.170 980.340 2385.910 1039.500 ;
        RECT 2259.170 964.960 2344.570 980.340 ;
        RECT 2187.070 915.260 2344.570 964.960 ;
        RECT 2348.470 915.260 2363.170 980.340 ;
        RECT 2367.070 964.960 2385.910 980.340 ;
        RECT 2389.810 964.960 2405.230 1056.000 ;
        RECT 2409.130 964.960 2524.570 1056.000 ;
        RECT 2367.070 915.260 2524.570 964.960 ;
        RECT 2187.070 887.360 2524.570 915.260 ;
        RECT 2187.070 875.200 2188.110 887.360 ;
        RECT 2192.010 875.200 2207.430 887.360 ;
        RECT 2211.330 876.000 2524.570 887.360 ;
        RECT 2211.330 875.200 2212.030 876.000 ;
        RECT 2187.070 796.320 2212.030 875.200 ;
        RECT 2215.930 796.320 2231.350 876.000 ;
        RECT 2235.250 796.320 2524.570 876.000 ;
        RECT 2187.070 775.840 2524.570 796.320 ;
        RECT 2187.070 750.080 2213.870 775.840 ;
        RECT 2217.770 750.080 2233.190 775.840 ;
        RECT 2237.090 765.395 2524.570 775.840 ;
        RECT 2237.090 750.080 2344.570 765.395 ;
        RECT 2187.070 740.480 2344.570 750.080 ;
        RECT 2187.070 652.160 2235.950 740.480 ;
        RECT 2239.850 652.160 2255.270 740.480 ;
        RECT 2259.170 725.500 2344.570 740.480 ;
        RECT 2348.470 725.500 2363.170 765.395 ;
        RECT 2367.070 740.480 2524.570 765.395 ;
        RECT 2367.070 725.500 2385.910 740.480 ;
        RECT 2259.170 666.340 2385.910 725.500 ;
        RECT 2259.170 652.160 2344.570 666.340 ;
        RECT 2187.070 604.480 2344.570 652.160 ;
        RECT 2187.070 516.160 2212.030 604.480 ;
        RECT 2215.930 516.160 2231.350 604.480 ;
        RECT 2235.250 601.260 2344.570 604.480 ;
        RECT 2348.470 601.260 2363.170 666.340 ;
        RECT 2367.070 652.160 2385.910 666.340 ;
        RECT 2389.810 652.160 2405.230 740.480 ;
        RECT 2409.130 652.160 2524.570 740.480 ;
        RECT 2367.070 601.260 2524.570 652.160 ;
        RECT 2235.250 516.160 2524.570 601.260 ;
        RECT 2187.070 463.040 2524.570 516.160 ;
        RECT 2187.070 437.280 2213.870 463.040 ;
        RECT 2217.770 437.280 2233.190 463.040 ;
        RECT 2237.090 451.395 2524.570 463.040 ;
        RECT 2237.090 437.280 2344.570 451.395 ;
        RECT 2187.070 427.680 2344.570 437.280 ;
        RECT 2187.070 336.640 2235.950 427.680 ;
        RECT 2239.850 336.640 2255.270 427.680 ;
        RECT 2259.170 411.500 2344.570 427.680 ;
        RECT 2348.470 411.500 2363.170 451.395 ;
        RECT 2367.070 427.680 2524.570 451.395 ;
        RECT 2367.070 411.500 2385.910 427.680 ;
        RECT 2259.170 352.340 2385.910 411.500 ;
        RECT 2259.170 336.640 2344.570 352.340 ;
        RECT 2187.070 253.600 2344.570 336.640 ;
        RECT 2187.070 165.280 2235.950 253.600 ;
        RECT 2239.850 165.280 2255.270 253.600 ;
        RECT 2259.170 239.500 2344.570 253.600 ;
        RECT 2348.470 239.500 2363.170 352.340 ;
        RECT 2367.070 336.640 2385.910 352.340 ;
        RECT 2389.810 336.640 2405.230 427.680 ;
        RECT 2409.130 336.640 2524.570 427.680 ;
        RECT 2367.070 253.600 2524.570 336.640 ;
        RECT 2367.070 239.500 2385.910 253.600 ;
        RECT 2259.170 180.340 2385.910 239.500 ;
        RECT 2259.170 165.280 2344.570 180.340 ;
        RECT 2187.070 63.500 2344.570 165.280 ;
        RECT 2348.470 63.500 2363.170 180.340 ;
        RECT 2187.070 14.640 2363.170 63.500 ;
        RECT 2367.070 165.280 2385.910 180.340 ;
        RECT 2389.810 165.280 2405.230 253.600 ;
        RECT 2409.130 165.280 2524.570 253.600 ;
        RECT 2367.070 14.640 2524.570 165.280 ;
        RECT 2528.470 14.640 2543.170 3488.760 ;
        RECT 2547.070 3378.565 2704.570 3488.760 ;
        RECT 2708.470 3378.565 2723.170 3488.760 ;
        RECT 2727.070 3378.565 2880.175 3488.760 ;
        RECT 2547.070 3373.440 2880.175 3378.565 ;
        RECT 2547.070 3319.040 2832.110 3373.440 ;
        RECT 2547.070 3277.395 2829.350 3319.040 ;
        RECT 2839.690 3318.640 2880.175 3373.440 ;
        RECT 2547.070 3064.565 2704.570 3277.395 ;
        RECT 2708.470 3064.565 2723.170 3277.395 ;
        RECT 2727.070 3263.360 2829.350 3277.395 ;
        RECT 2836.930 3263.360 2880.175 3318.640 ;
        RECT 2727.070 3064.565 2880.175 3263.360 ;
        RECT 2547.070 3057.920 2880.175 3064.565 ;
        RECT 2547.070 3003.520 2832.110 3057.920 ;
        RECT 2547.070 2963.395 2829.350 3003.520 ;
        RECT 2839.690 3003.120 2880.175 3057.920 ;
        RECT 2547.070 2750.565 2704.570 2963.395 ;
        RECT 2708.470 2750.565 2723.170 2963.395 ;
        RECT 2727.070 2950.560 2829.350 2963.395 ;
        RECT 2836.930 2950.560 2880.175 3003.120 ;
        RECT 2727.070 2750.565 2880.175 2950.560 ;
        RECT 2547.070 2745.120 2880.175 2750.565 ;
        RECT 2547.070 2690.720 2832.110 2745.120 ;
        RECT 2547.070 2649.395 2829.350 2690.720 ;
        RECT 2839.690 2690.320 2880.175 2745.120 ;
        RECT 2547.070 2436.565 2704.570 2649.395 ;
        RECT 2708.470 2611.840 2723.170 2649.395 ;
        RECT 2708.470 2545.280 2715.270 2611.840 ;
        RECT 2719.170 2545.280 2723.170 2611.840 ;
        RECT 2708.470 2436.565 2723.170 2545.280 ;
        RECT 2727.070 2635.040 2829.350 2649.395 ;
        RECT 2836.930 2635.040 2880.175 2690.320 ;
        RECT 2727.070 2436.565 2880.175 2635.040 ;
        RECT 2547.070 2429.600 2880.175 2436.565 ;
        RECT 2547.070 2375.200 2836.710 2429.600 ;
        RECT 2547.070 2335.395 2810.030 2375.200 ;
        RECT 2547.070 2122.565 2704.570 2335.395 ;
        RECT 2708.470 2122.565 2723.170 2335.395 ;
        RECT 2727.070 2322.240 2810.030 2335.395 ;
        RECT 2813.930 2322.240 2829.350 2375.200 ;
        RECT 2833.250 2368.480 2836.710 2375.200 ;
        RECT 2844.290 2368.480 2880.175 2429.600 ;
        RECT 2833.250 2322.240 2880.175 2368.480 ;
        RECT 2727.070 2122.565 2880.175 2322.240 ;
        RECT 2547.070 2116.800 2880.175 2122.565 ;
        RECT 2547.070 2062.400 2832.110 2116.800 ;
        RECT 2547.070 2021.395 2829.350 2062.400 ;
        RECT 2839.690 2062.000 2880.175 2116.800 ;
        RECT 2547.070 1808.565 2704.570 2021.395 ;
        RECT 2708.470 1808.565 2723.170 2021.395 ;
        RECT 2727.070 2006.720 2829.350 2021.395 ;
        RECT 2836.930 2006.720 2880.175 2062.000 ;
        RECT 2727.070 1808.565 2880.175 2006.720 ;
        RECT 2547.070 1804.000 2880.175 1808.565 ;
        RECT 2547.070 1746.880 2836.710 1804.000 ;
        RECT 2547.070 1707.395 2810.030 1746.880 ;
        RECT 2547.070 1494.565 2704.570 1707.395 ;
        RECT 2708.470 1670.720 2723.170 1707.395 ;
        RECT 2708.470 1604.160 2715.270 1670.720 ;
        RECT 2719.170 1604.160 2723.170 1670.720 ;
        RECT 2708.470 1494.565 2723.170 1604.160 ;
        RECT 2727.070 1693.920 2810.030 1707.395 ;
        RECT 2813.930 1693.920 2829.350 1746.880 ;
        RECT 2833.250 1737.440 2836.710 1746.880 ;
        RECT 2844.290 1737.440 2880.175 1804.000 ;
        RECT 2833.250 1693.920 2880.175 1737.440 ;
        RECT 2727.070 1494.565 2880.175 1693.920 ;
        RECT 2547.070 1488.480 2880.175 1494.565 ;
        RECT 2547.070 1434.080 2832.110 1488.480 ;
        RECT 2547.070 1393.395 2829.350 1434.080 ;
        RECT 2839.690 1433.680 2880.175 1488.480 ;
        RECT 2547.070 1180.565 2704.570 1393.395 ;
        RECT 2708.470 1180.565 2723.170 1393.395 ;
        RECT 2727.070 1378.400 2829.350 1393.395 ;
        RECT 2836.930 1378.400 2880.175 1433.680 ;
        RECT 2727.070 1180.565 2880.175 1378.400 ;
        RECT 2547.070 1175.680 2880.175 1180.565 ;
        RECT 2547.070 1118.560 2836.710 1175.680 ;
        RECT 2547.070 1079.395 2810.030 1118.560 ;
        RECT 2547.070 866.565 2704.570 1079.395 ;
        RECT 2708.470 866.565 2723.170 1079.395 ;
        RECT 2727.070 1065.600 2810.030 1079.395 ;
        RECT 2813.930 1065.600 2829.350 1118.560 ;
        RECT 2833.250 1111.840 2836.710 1118.560 ;
        RECT 2844.290 1111.840 2880.175 1175.680 ;
        RECT 2833.250 1065.600 2880.175 1111.840 ;
        RECT 2727.070 866.565 2880.175 1065.600 ;
        RECT 2547.070 860.160 2880.175 866.565 ;
        RECT 2547.070 805.760 2832.110 860.160 ;
        RECT 2547.070 765.395 2829.350 805.760 ;
        RECT 2839.690 805.360 2880.175 860.160 ;
        RECT 2547.070 552.565 2704.570 765.395 ;
        RECT 2708.470 552.565 2723.170 765.395 ;
        RECT 2727.070 750.080 2829.350 765.395 ;
        RECT 2836.930 750.080 2880.175 805.360 ;
        RECT 2727.070 552.565 2880.175 750.080 ;
        RECT 2547.070 547.360 2880.175 552.565 ;
        RECT 2547.070 525.600 2832.110 547.360 ;
        RECT 2547.070 451.395 2829.350 525.600 ;
        RECT 2839.690 525.200 2880.175 547.360 ;
        RECT 2547.070 14.640 2704.570 451.395 ;
        RECT 2708.470 414.080 2723.170 451.395 ;
        RECT 2708.470 347.520 2715.270 414.080 ;
        RECT 2719.170 347.520 2723.170 414.080 ;
        RECT 2708.470 14.640 2723.170 347.520 ;
        RECT 2727.070 437.280 2829.350 451.395 ;
        RECT 2836.930 437.280 2880.175 525.200 ;
        RECT 2727.070 14.640 2880.175 437.280 ;
  END
END user_project_wrapper
END LIBRARY

