magic
tech sky130A
magscale 1 2
timestamp 1710358026
<< obsli1 >>
rect 1104 2159 4876 8721
<< obsm1 >>
rect 1104 2128 5138 8752
<< metal2 >>
rect 2962 10200 3018 11000
<< obsm2 >>
rect 1421 10144 2906 10282
rect 3074 10144 5134 10282
rect 1421 1391 5134 10144
<< metal3 >>
rect 5200 9528 6000 9648
rect 0 8168 800 8288
rect 5200 6808 6000 6928
rect 5200 4088 6000 4208
rect 5200 1368 6000 1488
<< obsm3 >>
rect 800 9448 5120 9621
rect 800 8368 5200 9448
rect 880 8088 5200 8368
rect 800 7008 5200 8088
rect 800 6728 5120 7008
rect 800 4288 5200 6728
rect 800 4008 5120 4288
rect 800 1568 5200 4008
rect 800 1395 5120 1568
<< metal4 >>
rect 1415 2128 1735 8752
rect 1886 2128 2206 8752
rect 2358 2128 2678 8752
rect 2829 2128 3149 8752
rect 3301 2128 3621 8752
rect 3772 2128 4092 8752
rect 4244 2128 4564 8752
rect 4715 2128 5035 8752
<< labels >>
rlabel metal3 s 5200 6808 6000 6928 6 bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal output
rlabel metal3 s 5200 9528 6000 9648 6 bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 2 nsew signal input
rlabel metal3 s 5200 1368 6000 1488 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 5200 4088 6000 4208 6 ccff_tail
port 4 nsew signal output
rlabel metal2 s 2962 10200 3018 11000 6 gfpga_pad_GPIO_PAD
port 5 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 prog_clk
port 6 nsew signal input
rlabel metal4 s 1415 2128 1735 8752 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 2358 2128 2678 8752 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 3301 2128 3621 8752 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 4244 2128 4564 8752 6 vdd
port 7 nsew power bidirectional
rlabel metal4 s 1886 2128 2206 8752 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 2829 2128 3149 8752 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 3772 2128 4092 8752 6 vss
port 8 nsew ground bidirectional
rlabel metal4 s 4715 2128 5035 8752 6 vss
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 11000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 120000
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/grid_io_top_out/runs/24_03_13_13_26/results/signoff/grid_io_top_out.magic.gds
string GDS_START 47994
<< end >>

