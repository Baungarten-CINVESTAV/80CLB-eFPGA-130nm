magic
tech sky130A
magscale 1 2
timestamp 1708041581
<< viali >>
rect 13737 17289 13771 17323
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 3893 17153 3927 17187
rect 4261 17153 4295 17187
rect 5457 17153 5491 17187
rect 5641 17153 5675 17187
rect 6837 17153 6871 17187
rect 8033 17153 8067 17187
rect 9413 17153 9447 17187
rect 10977 17153 11011 17187
rect 12357 17153 12391 17187
rect 13093 17153 13127 17187
rect 13829 17153 13863 17187
rect 14197 17153 14231 17187
rect 1869 17017 1903 17051
rect 4077 17017 4111 17051
rect 1593 16949 1627 16983
rect 1961 16949 1995 16983
rect 2237 16949 2271 16983
rect 2697 16949 2731 16983
rect 4445 16949 4479 16983
rect 5273 16949 5307 16983
rect 5825 16949 5859 16983
rect 6653 16949 6687 16983
rect 8217 16949 8251 16983
rect 9597 16949 9631 16983
rect 10793 16949 10827 16983
rect 12173 16949 12207 16983
rect 13277 16949 13311 16983
rect 14381 16949 14415 16983
rect 5641 16745 5675 16779
rect 2973 16677 3007 16711
rect 11713 16677 11747 16711
rect 13369 16677 13403 16711
rect 3985 16609 4019 16643
rect 6377 16609 6411 16643
rect 7941 16609 7975 16643
rect 1777 16541 1811 16575
rect 1869 16541 1903 16575
rect 2789 16541 2823 16575
rect 3065 16541 3099 16575
rect 3525 16541 3559 16575
rect 3801 16541 3835 16575
rect 5457 16541 5491 16575
rect 6561 16541 6595 16575
rect 6745 16541 6779 16575
rect 7113 16541 7147 16575
rect 7205 16541 7239 16575
rect 7757 16541 7791 16575
rect 9413 16541 9447 16575
rect 9873 16541 9907 16575
rect 10793 16541 10827 16575
rect 11805 16541 11839 16575
rect 13093 16541 13127 16575
rect 13553 16541 13587 16575
rect 13737 16541 13771 16575
rect 14197 16541 14231 16575
rect 4721 16473 4755 16507
rect 4813 16473 4847 16507
rect 5365 16473 5399 16507
rect 9505 16473 9539 16507
rect 1685 16405 1719 16439
rect 2053 16405 2087 16439
rect 3249 16405 3283 16439
rect 4445 16405 4479 16439
rect 5917 16405 5951 16439
rect 6929 16405 6963 16439
rect 7297 16405 7331 16439
rect 10057 16405 10091 16439
rect 10701 16405 10735 16439
rect 13001 16405 13035 16439
rect 13829 16405 13863 16439
rect 14381 16405 14415 16439
rect 2605 16201 2639 16235
rect 3341 16201 3375 16235
rect 5549 16201 5583 16235
rect 7205 16201 7239 16235
rect 7481 16201 7515 16235
rect 9321 16201 9355 16235
rect 14197 16201 14231 16235
rect 4537 16133 4571 16167
rect 5089 16133 5123 16167
rect 8125 16133 8159 16167
rect 1777 16065 1811 16099
rect 2053 16065 2087 16099
rect 2421 16065 2455 16099
rect 2881 16065 2915 16099
rect 3065 16065 3099 16099
rect 3525 16065 3559 16099
rect 3801 16065 3835 16099
rect 5273 16065 5307 16099
rect 7297 16065 7331 16099
rect 9137 16065 9171 16099
rect 10149 16065 10183 16099
rect 10609 16065 10643 16099
rect 14105 16065 14139 16099
rect 3617 15997 3651 16031
rect 4445 15997 4479 16031
rect 6009 15997 6043 16031
rect 6193 15997 6227 16031
rect 6561 15997 6595 16031
rect 6745 15997 6779 16031
rect 8217 15997 8251 16031
rect 10793 15997 10827 16031
rect 1869 15929 1903 15963
rect 4261 15929 4295 15963
rect 7665 15929 7699 15963
rect 1685 15861 1719 15895
rect 2789 15861 2823 15895
rect 3157 15861 3191 15895
rect 5365 15861 5399 15895
rect 10333 15861 10367 15895
rect 11069 15861 11103 15895
rect 4077 15657 4111 15691
rect 4721 15657 4755 15691
rect 6193 15657 6227 15691
rect 7481 15657 7515 15691
rect 11161 15657 11195 15691
rect 14381 15657 14415 15691
rect 4261 15589 4295 15623
rect 6561 15589 6595 15623
rect 2237 15521 2271 15555
rect 2421 15521 2455 15555
rect 4905 15521 4939 15555
rect 5089 15521 5123 15555
rect 1409 15453 1443 15487
rect 1869 15453 1903 15487
rect 2145 15453 2179 15487
rect 3617 15453 3651 15487
rect 3893 15453 3927 15487
rect 4169 15453 4203 15487
rect 5917 15453 5951 15487
rect 6101 15453 6135 15487
rect 6377 15453 6411 15487
rect 7205 15453 7239 15487
rect 7389 15453 7423 15487
rect 9505 15453 9539 15487
rect 9873 15453 9907 15487
rect 9965 15453 9999 15487
rect 10425 15453 10459 15487
rect 10609 15453 10643 15487
rect 11069 15453 11103 15487
rect 11345 15453 11379 15487
rect 14197 15453 14231 15487
rect 2881 15385 2915 15419
rect 7757 15385 7791 15419
rect 8309 15385 8343 15419
rect 8401 15385 8435 15419
rect 8585 15385 8619 15419
rect 1593 15317 1627 15351
rect 1685 15317 1719 15351
rect 2053 15317 2087 15351
rect 2973 15317 3007 15351
rect 5365 15317 5399 15351
rect 6653 15317 6687 15351
rect 8953 15317 8987 15351
rect 9689 15317 9723 15351
rect 10057 15317 10091 15351
rect 4261 15113 4295 15147
rect 6101 15113 6135 15147
rect 8033 15113 8067 15147
rect 9505 15113 9539 15147
rect 3056 15045 3090 15079
rect 5374 15045 5408 15079
rect 6644 15045 6678 15079
rect 8392 15045 8426 15079
rect 1593 14977 1627 15011
rect 1685 14977 1719 15011
rect 5917 14977 5951 15011
rect 6009 14977 6043 15011
rect 7849 14977 7883 15011
rect 9597 14977 9631 15011
rect 9781 14977 9815 15011
rect 10333 14977 10367 15011
rect 11161 14977 11195 15011
rect 11253 14977 11287 15011
rect 12449 14977 12483 15011
rect 13001 14977 13035 15011
rect 13093 14977 13127 15011
rect 14197 14977 14231 15011
rect 1869 14909 1903 14943
rect 2421 14909 2455 14943
rect 2789 14909 2823 14943
rect 5641 14909 5675 14943
rect 6377 14909 6411 14943
rect 8125 14909 8159 14943
rect 10517 14909 10551 14943
rect 11529 14909 11563 14943
rect 11713 14909 11747 14943
rect 12357 14909 12391 14943
rect 12725 14909 12759 14943
rect 1501 14841 1535 14875
rect 10241 14841 10275 14875
rect 10701 14841 10735 14875
rect 2053 14773 2087 14807
rect 4169 14773 4203 14807
rect 5825 14773 5859 14807
rect 7757 14773 7791 14807
rect 12173 14773 12207 14807
rect 12909 14773 12943 14807
rect 13277 14773 13311 14807
rect 14381 14773 14415 14807
rect 2053 14569 2087 14603
rect 6653 14569 6687 14603
rect 8125 14569 8159 14603
rect 8493 14569 8527 14603
rect 10149 14569 10183 14603
rect 10517 14569 10551 14603
rect 10793 14569 10827 14603
rect 14197 14569 14231 14603
rect 2513 14501 2547 14535
rect 3433 14501 3467 14535
rect 4077 14501 4111 14535
rect 13185 14501 13219 14535
rect 13645 14501 13679 14535
rect 2421 14433 2455 14467
rect 4445 14433 4479 14467
rect 8033 14433 8067 14467
rect 11069 14433 11103 14467
rect 12725 14433 12759 14467
rect 1501 14365 1535 14399
rect 2237 14365 2271 14399
rect 2697 14365 2731 14399
rect 2973 14365 3007 14399
rect 3249 14365 3283 14399
rect 3893 14365 3927 14399
rect 4353 14365 4387 14399
rect 6561 14365 6595 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 10057 14365 10091 14399
rect 10333 14365 10367 14399
rect 10609 14365 10643 14399
rect 10701 14365 10735 14399
rect 12541 14365 12575 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 14105 14365 14139 14399
rect 4261 14297 4295 14331
rect 6316 14297 6350 14331
rect 7766 14297 7800 14331
rect 9413 14297 9447 14331
rect 11314 14297 11348 14331
rect 1593 14229 1627 14263
rect 2789 14229 2823 14263
rect 5089 14229 5123 14263
rect 5181 14229 5215 14263
rect 12449 14229 12483 14263
rect 3525 14025 3559 14059
rect 7113 14025 7147 14059
rect 7389 14025 7423 14059
rect 9505 14025 9539 14059
rect 12173 14025 12207 14059
rect 12265 14025 12299 14059
rect 13185 14025 13219 14059
rect 13921 14025 13955 14059
rect 4660 13957 4694 13991
rect 14105 13957 14139 13991
rect 1593 13889 1627 13923
rect 3157 13889 3191 13923
rect 4905 13889 4939 13923
rect 4997 13889 5031 13923
rect 5181 13889 5215 13923
rect 5733 13889 5767 13923
rect 6929 13889 6963 13923
rect 7205 13889 7239 13923
rect 7941 13889 7975 13923
rect 8493 13889 8527 13923
rect 9321 13889 9355 13923
rect 9781 13889 9815 13923
rect 10609 13889 10643 13923
rect 11345 13889 11379 13923
rect 11529 13889 11563 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 13737 13889 13771 13923
rect 1685 13821 1719 13855
rect 2329 13821 2363 13855
rect 2513 13821 2547 13855
rect 8125 13821 8159 13855
rect 8217 13821 8251 13855
rect 9965 13821 9999 13855
rect 10149 13821 10183 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 11713 13821 11747 13855
rect 12725 13821 12759 13855
rect 14381 13821 14415 13855
rect 8677 13753 8711 13787
rect 9597 13753 9631 13787
rect 1869 13685 1903 13719
rect 2605 13685 2639 13719
rect 5365 13685 5399 13719
rect 5825 13685 5859 13719
rect 7757 13685 7791 13719
rect 2881 13481 2915 13515
rect 4537 13481 4571 13515
rect 10793 13481 10827 13515
rect 11437 13481 11471 13515
rect 12265 13481 12299 13515
rect 12909 13481 12943 13515
rect 5641 13413 5675 13447
rect 12633 13413 12667 13447
rect 2789 13345 2823 13379
rect 3525 13345 3559 13379
rect 4721 13345 4755 13379
rect 5917 13345 5951 13379
rect 8217 13345 8251 13379
rect 9413 13345 9447 13379
rect 10057 13345 10091 13379
rect 12081 13345 12115 13379
rect 2522 13277 2556 13311
rect 3341 13277 3375 13311
rect 4905 13277 4939 13311
rect 5181 13277 5215 13311
rect 5457 13277 5491 13311
rect 5733 13277 5767 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 7757 13277 7791 13311
rect 10885 13277 10919 13311
rect 11161 13277 11195 13311
rect 12333 13271 12367 13305
rect 12449 13273 12483 13307
rect 12725 13277 12759 13311
rect 13737 13277 13771 13311
rect 14197 13277 14231 13311
rect 7113 13209 7147 13243
rect 9045 13209 9079 13243
rect 9137 13209 9171 13243
rect 1409 13141 1443 13175
rect 5365 13141 5399 13175
rect 6377 13141 6411 13175
rect 7205 13141 7239 13175
rect 8769 13141 8803 13175
rect 10609 13141 10643 13175
rect 11345 13141 11379 13175
rect 13921 13141 13955 13175
rect 14381 13141 14415 13175
rect 2697 12937 2731 12971
rect 6193 12937 6227 12971
rect 6837 12937 6871 12971
rect 8401 12937 8435 12971
rect 10885 12937 10919 12971
rect 4169 12869 4203 12903
rect 12173 12869 12207 12903
rect 1777 12801 1811 12835
rect 1869 12801 1903 12835
rect 2329 12801 2363 12835
rect 2605 12801 2639 12835
rect 3065 12801 3099 12835
rect 3249 12801 3283 12835
rect 4077 12801 4111 12835
rect 4353 12801 4387 12835
rect 4629 12801 4663 12835
rect 5549 12801 5583 12835
rect 6561 12801 6595 12835
rect 6929 12801 6963 12835
rect 7021 12801 7055 12835
rect 7288 12801 7322 12835
rect 8493 12801 8527 12835
rect 8760 12801 8794 12835
rect 11069 12801 11103 12835
rect 11161 12801 11195 12835
rect 12449 12825 12483 12859
rect 4813 12733 4847 12767
rect 5733 12733 5767 12767
rect 6469 12733 6503 12767
rect 10701 12733 10735 12767
rect 11529 12733 11563 12767
rect 11713 12733 11747 12767
rect 2513 12665 2547 12699
rect 2881 12665 2915 12699
rect 12265 12665 12299 12699
rect 1685 12597 1719 12631
rect 2053 12597 2087 12631
rect 3433 12597 3467 12631
rect 4537 12597 4571 12631
rect 5273 12597 5307 12631
rect 9873 12597 9907 12631
rect 10149 12597 10183 12631
rect 11253 12597 11287 12631
rect 2881 12393 2915 12427
rect 4445 12393 4479 12427
rect 4813 12393 4847 12427
rect 7113 12393 7147 12427
rect 11437 12393 11471 12427
rect 14381 12393 14415 12427
rect 11897 12325 11931 12359
rect 2973 12257 3007 12291
rect 3985 12257 4019 12291
rect 5641 12257 5675 12291
rect 7389 12257 7423 12291
rect 8033 12257 8067 12291
rect 11713 12257 11747 12291
rect 1409 12189 1443 12223
rect 2421 12189 2455 12223
rect 2689 12189 2723 12223
rect 3157 12189 3191 12223
rect 3801 12189 3835 12223
rect 4905 12189 4939 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 5733 12189 5767 12223
rect 7205 12189 7239 12223
rect 7941 12189 7975 12223
rect 8585 12189 8619 12223
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 10313 12189 10347 12223
rect 11529 12189 11563 12223
rect 14197 12189 14231 12223
rect 2513 12121 2547 12155
rect 6000 12121 6034 12155
rect 7849 12121 7883 12155
rect 9045 12121 9079 12155
rect 9137 12121 9171 12155
rect 9689 12121 9723 12155
rect 1593 12053 1627 12087
rect 3617 12053 3651 12087
rect 8677 12053 8711 12087
rect 9965 12053 9999 12087
rect 2421 11849 2455 11883
rect 4629 11849 4663 11883
rect 4905 11849 4939 11883
rect 7205 11849 7239 11883
rect 7481 11849 7515 11883
rect 10977 11849 11011 11883
rect 1409 11713 1443 11747
rect 1869 11713 1903 11747
rect 1961 11713 1995 11747
rect 2237 11713 2271 11747
rect 2513 11713 2547 11747
rect 3249 11713 3283 11747
rect 4721 11713 4755 11747
rect 5181 11713 5215 11747
rect 8125 11713 8159 11747
rect 8401 11713 8435 11747
rect 9965 11713 9999 11747
rect 13921 11713 13955 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 3433 11645 3467 11679
rect 3985 11645 4019 11679
rect 4169 11645 4203 11679
rect 6561 11645 6595 11679
rect 7941 11645 7975 11679
rect 10333 11645 10367 11679
rect 10517 11645 10551 11679
rect 11529 11645 11563 11679
rect 2145 11577 2179 11611
rect 4997 11577 5031 11611
rect 8217 11577 8251 11611
rect 10149 11577 10183 11611
rect 1501 11509 1535 11543
rect 1685 11509 1719 11543
rect 3157 11509 3191 11543
rect 3893 11509 3927 11543
rect 14381 11509 14415 11543
rect 3433 11305 3467 11339
rect 5273 11305 5307 11339
rect 6285 11305 6319 11339
rect 7389 11305 7423 11339
rect 3065 11237 3099 11271
rect 5365 11237 5399 11271
rect 7573 11237 7607 11271
rect 5825 11169 5859 11203
rect 9321 11169 9355 11203
rect 10057 11169 10091 11203
rect 11529 11169 11563 11203
rect 1593 11101 1627 11135
rect 2973 11101 3007 11135
rect 3525 11101 3559 11135
rect 5089 11101 5123 11135
rect 5549 11101 5583 11135
rect 5641 11101 5675 11135
rect 6837 11101 6871 11135
rect 7205 11101 7239 11135
rect 8217 11101 8251 11135
rect 8493 11101 8527 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10324 11101 10358 11135
rect 11713 11101 11747 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 1685 11033 1719 11067
rect 6745 10965 6779 10999
rect 7113 10965 7147 10999
rect 8309 10965 8343 10999
rect 11437 10965 11471 10999
rect 12173 10965 12207 10999
rect 11345 10761 11379 10795
rect 12173 10761 12207 10795
rect 1777 10625 1811 10659
rect 2053 10625 2087 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5273 10625 5307 10659
rect 5549 10625 5583 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 7849 10625 7883 10659
rect 9689 10625 9723 10659
rect 9965 10625 9999 10659
rect 10241 10625 10275 10659
rect 11161 10625 11195 10659
rect 11529 10625 11563 10659
rect 12449 10625 12483 10659
rect 14197 10625 14231 10659
rect 5733 10557 5767 10591
rect 7113 10557 7147 10591
rect 7297 10557 7331 10591
rect 9781 10557 9815 10591
rect 11713 10557 11747 10591
rect 1869 10489 1903 10523
rect 4905 10489 4939 10523
rect 5457 10489 5491 10523
rect 10057 10489 10091 10523
rect 12265 10489 12299 10523
rect 1685 10421 1719 10455
rect 5089 10421 5123 10455
rect 6009 10421 6043 10455
rect 7021 10421 7055 10455
rect 7757 10421 7791 10455
rect 9137 10421 9171 10455
rect 10333 10421 10367 10455
rect 14381 10421 14415 10455
rect 12081 10217 12115 10251
rect 3801 10149 3835 10183
rect 9045 10149 9079 10183
rect 11161 10149 11195 10183
rect 11621 10149 11655 10183
rect 10517 10081 10551 10115
rect 11253 10081 11287 10115
rect 11437 10081 11471 10115
rect 3166 10013 3200 10047
rect 3433 10013 3467 10047
rect 5181 10013 5215 10047
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 8585 10013 8619 10047
rect 10425 10013 10459 10047
rect 10701 10013 10735 10047
rect 12173 10013 12207 10047
rect 1777 9945 1811 9979
rect 4914 9945 4948 9979
rect 5273 9945 5307 9979
rect 7358 9945 7392 9979
rect 10158 9945 10192 9979
rect 13553 9945 13587 9979
rect 1501 9877 1535 9911
rect 2053 9877 2087 9911
rect 8493 9877 8527 9911
rect 8769 9877 8803 9911
rect 13829 9877 13863 9911
rect 4537 9673 4571 9707
rect 6193 9673 6227 9707
rect 10057 9673 10091 9707
rect 1777 9537 1811 9571
rect 2881 9537 2915 9571
rect 3065 9537 3099 9571
rect 3525 9537 3559 9571
rect 3617 9537 3651 9571
rect 5273 9537 5307 9571
rect 5549 9537 5583 9571
rect 5733 9537 5767 9571
rect 6377 9537 6411 9571
rect 7297 9537 7331 9571
rect 9137 9537 9171 9571
rect 9505 9537 9539 9571
rect 10793 9537 10827 9571
rect 11161 9537 11195 9571
rect 11253 9537 11287 9571
rect 11529 9537 11563 9571
rect 3893 9469 3927 9503
rect 5089 9469 5123 9503
rect 6561 9469 6595 9503
rect 10977 9469 11011 9503
rect 11713 9469 11747 9503
rect 12265 9469 12299 9503
rect 3433 9401 3467 9435
rect 8585 9401 8619 9435
rect 1685 9333 1719 9367
rect 2237 9333 2271 9367
rect 3157 9333 3191 9367
rect 3709 9333 3743 9367
rect 4721 9333 4755 9367
rect 7021 9333 7055 9367
rect 9229 9333 9263 9367
rect 10425 9333 10459 9367
rect 11897 9333 11931 9367
rect 3617 9129 3651 9163
rect 4721 9129 4755 9163
rect 7205 9129 7239 9163
rect 10333 9129 10367 9163
rect 10517 9129 10551 9163
rect 11805 9129 11839 9163
rect 13737 9129 13771 9163
rect 14381 9129 14415 9163
rect 9781 9061 9815 9095
rect 11069 9061 11103 9095
rect 12265 9061 12299 9095
rect 12541 9061 12575 9095
rect 4905 8993 4939 9027
rect 5181 8993 5215 9027
rect 7849 8993 7883 9027
rect 9229 8993 9263 9027
rect 11989 8993 12023 9027
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 2493 8925 2527 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 5641 8925 5675 8959
rect 8677 8925 8711 8959
rect 10149 8925 10183 8959
rect 10425 8925 10459 8959
rect 10701 8925 10735 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 12173 8925 12207 8959
rect 12449 8925 12483 8959
rect 12725 8925 12759 8959
rect 13921 8925 13955 8959
rect 14197 8925 14231 8959
rect 1409 8857 1443 8891
rect 4997 8857 5031 8891
rect 5908 8857 5942 8891
rect 8125 8857 8159 8891
rect 9321 8857 9355 8891
rect 3985 8789 4019 8823
rect 7021 8789 7055 8823
rect 9965 8789 9999 8823
rect 10793 8789 10827 8823
rect 1869 8585 1903 8619
rect 3709 8585 3743 8619
rect 4261 8585 4295 8619
rect 4537 8585 4571 8619
rect 7941 8585 7975 8619
rect 10701 8585 10735 8619
rect 11161 8585 11195 8619
rect 4813 8517 4847 8551
rect 9045 8517 9079 8551
rect 9137 8517 9171 8551
rect 9689 8517 9723 8551
rect 13093 8517 13127 8551
rect 13185 8517 13219 8551
rect 2982 8449 3016 8483
rect 3525 8449 3559 8483
rect 3801 8449 3835 8483
rect 4077 8449 4111 8483
rect 4353 8449 4387 8483
rect 6745 8449 6779 8483
rect 8861 8449 8895 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 11069 8449 11103 8483
rect 12653 8449 12687 8483
rect 12909 8449 12943 8483
rect 14105 8449 14139 8483
rect 3249 8381 3283 8415
rect 4721 8381 4755 8415
rect 4997 8381 5031 8415
rect 6101 8381 6135 8415
rect 6561 8381 6595 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 7481 8381 7515 8415
rect 8677 8381 8711 8415
rect 9781 8381 9815 8415
rect 9965 8381 9999 8415
rect 13369 8381 13403 8415
rect 3985 8313 4019 8347
rect 10977 8313 11011 8347
rect 11529 8313 11563 8347
rect 14381 8313 14415 8347
rect 5457 8245 5491 8279
rect 8217 8245 8251 8279
rect 10149 8245 10183 8279
rect 7205 8041 7239 8075
rect 7665 8041 7699 8075
rect 9045 8041 9079 8075
rect 10149 8041 10183 8075
rect 12817 8041 12851 8075
rect 14105 8041 14139 8075
rect 6285 7973 6319 8007
rect 10057 7973 10091 8007
rect 11345 7973 11379 8007
rect 12633 7973 12667 8007
rect 13737 7973 13771 8007
rect 4261 7905 4295 7939
rect 4629 7905 4663 7939
rect 6929 7905 6963 7939
rect 8769 7905 8803 7939
rect 9413 7905 9447 7939
rect 10609 7905 10643 7939
rect 10793 7905 10827 7939
rect 13369 7905 13403 7939
rect 1409 7837 1443 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 4445 7837 4479 7871
rect 4905 7837 4939 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9597 7837 9631 7871
rect 10333 7837 10367 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 13553 7837 13587 7871
rect 14289 7837 14323 7871
rect 1777 7769 1811 7803
rect 2053 7769 2087 7803
rect 5172 7769 5206 7803
rect 8125 7769 8159 7803
rect 11253 7769 11287 7803
rect 12081 7769 12115 7803
rect 12173 7769 12207 7803
rect 2513 7701 2547 7735
rect 3525 7701 3559 7735
rect 3801 7701 3835 7735
rect 6469 7701 6503 7735
rect 8033 7701 8067 7735
rect 11805 7701 11839 7735
rect 4261 7497 4295 7531
rect 5273 7497 5307 7531
rect 6193 7497 6227 7531
rect 7297 7497 7331 7531
rect 8585 7497 8619 7531
rect 9045 7497 9079 7531
rect 10885 7497 10919 7531
rect 12909 7429 12943 7463
rect 1777 7361 1811 7395
rect 2329 7361 2363 7395
rect 3157 7361 3191 7395
rect 3525 7361 3559 7395
rect 4445 7361 4479 7395
rect 4905 7361 4939 7395
rect 4997 7361 5031 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 7113 7361 7147 7395
rect 8125 7361 8159 7395
rect 8401 7361 8435 7395
rect 8861 7361 8895 7395
rect 9137 7361 9171 7395
rect 9588 7361 9622 7395
rect 10977 7361 11011 7395
rect 11069 7361 11103 7395
rect 11161 7361 11195 7395
rect 12449 7361 12483 7395
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 14197 7361 14231 7395
rect 2237 7293 2271 7327
rect 2605 7293 2639 7327
rect 3709 7293 3743 7327
rect 6377 7293 6411 7327
rect 6561 7293 6595 7327
rect 7389 7293 7423 7327
rect 7573 7293 7607 7327
rect 9321 7293 9355 7327
rect 12081 7293 12115 7327
rect 12265 7293 12299 7327
rect 2513 7225 2547 7259
rect 4813 7225 4847 7259
rect 8769 7225 8803 7259
rect 10701 7225 10735 7259
rect 1501 7157 1535 7191
rect 4169 7157 4203 7191
rect 5181 7157 5215 7191
rect 6929 7157 6963 7191
rect 7757 7157 7791 7191
rect 8309 7157 8343 7191
rect 11529 7157 11563 7191
rect 14381 7157 14415 7191
rect 1685 6953 1719 6987
rect 3525 6953 3559 6987
rect 5365 6953 5399 6987
rect 9873 6953 9907 6987
rect 7297 6885 7331 6919
rect 11989 6885 12023 6919
rect 1869 6817 1903 6851
rect 2605 6817 2639 6851
rect 3985 6817 4019 6851
rect 6745 6817 6779 6851
rect 6929 6817 6963 6851
rect 7113 6817 7147 6851
rect 8033 6817 8067 6851
rect 10609 6817 10643 6851
rect 12817 6817 12851 6851
rect 13185 6817 13219 6851
rect 1777 6749 1811 6783
rect 2053 6749 2087 6783
rect 2789 6749 2823 6783
rect 3341 6749 3375 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 7757 6749 7791 6783
rect 8217 6749 8251 6783
rect 10517 6749 10551 6783
rect 10876 6749 10910 6783
rect 13001 6749 13035 6783
rect 13093 6749 13127 6783
rect 14197 6749 14231 6783
rect 4252 6681 4286 6715
rect 5457 6681 5491 6715
rect 6009 6681 6043 6715
rect 6101 6681 6135 6715
rect 2513 6613 2547 6647
rect 3249 6613 3283 6647
rect 6561 6613 6595 6647
rect 7941 6613 7975 6647
rect 8677 6613 8711 6647
rect 12357 6613 12391 6647
rect 14381 6613 14415 6647
rect 2053 6409 2087 6443
rect 2421 6409 2455 6443
rect 3341 6409 3375 6443
rect 3893 6409 3927 6443
rect 4169 6409 4203 6443
rect 6193 6409 6227 6443
rect 6469 6409 6503 6443
rect 7297 6409 7331 6443
rect 7941 6409 7975 6443
rect 8861 6409 8895 6443
rect 10701 6409 10735 6443
rect 4905 6341 4939 6375
rect 5457 6341 5491 6375
rect 7757 6341 7791 6375
rect 1409 6273 1443 6307
rect 1777 6273 1811 6307
rect 2145 6273 2179 6307
rect 2237 6273 2271 6307
rect 2697 6273 2731 6307
rect 3525 6273 3559 6307
rect 3617 6273 3651 6307
rect 4077 6273 4111 6307
rect 6009 6273 6043 6307
rect 6377 6273 6411 6307
rect 6837 6273 6871 6307
rect 7573 6273 7607 6307
rect 7849 6273 7883 6307
rect 8125 6273 8159 6307
rect 9137 6273 9171 6307
rect 9505 6273 9539 6307
rect 9965 6273 9999 6307
rect 4813 6205 4847 6239
rect 5549 6205 5583 6239
rect 5733 6205 5767 6239
rect 6653 6205 6687 6239
rect 8217 6205 8251 6239
rect 8401 6205 8435 6239
rect 9045 6205 9079 6239
rect 10057 6205 10091 6239
rect 10241 6205 10275 6239
rect 2513 6137 2547 6171
rect 7389 6137 7423 6171
rect 9781 6137 9815 6171
rect 3801 6069 3835 6103
rect 9689 6069 9723 6103
rect 2053 5865 2087 5899
rect 6469 5865 6503 5899
rect 6745 5865 6779 5899
rect 10333 5865 10367 5899
rect 14289 5865 14323 5899
rect 3341 5797 3375 5831
rect 2513 5729 2547 5763
rect 5089 5729 5123 5763
rect 8953 5729 8987 5763
rect 2145 5661 2179 5695
rect 3525 5661 3559 5695
rect 3985 5661 4019 5695
rect 4169 5661 4203 5695
rect 4629 5661 4663 5695
rect 6837 5661 6871 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 14105 5661 14139 5695
rect 1777 5593 1811 5627
rect 2605 5593 2639 5627
rect 3157 5593 3191 5627
rect 5356 5593 5390 5627
rect 7941 5593 7975 5627
rect 9198 5593 9232 5627
rect 13553 5593 13587 5627
rect 13921 5593 13955 5627
rect 1501 5525 1535 5559
rect 4997 5525 5031 5559
rect 2237 5321 2271 5355
rect 3065 5321 3099 5355
rect 9321 5321 9355 5355
rect 2421 5253 2455 5287
rect 4353 5253 4387 5287
rect 5365 5253 5399 5287
rect 5549 5253 5583 5287
rect 5641 5253 5675 5287
rect 6929 5253 6963 5287
rect 7849 5253 7883 5287
rect 9781 5253 9815 5287
rect 9873 5253 9907 5287
rect 10701 5253 10735 5287
rect 1777 5185 1811 5219
rect 2053 5185 2087 5219
rect 2513 5185 2547 5219
rect 4445 5185 4479 5219
rect 7297 5185 7331 5219
rect 14197 5185 14231 5219
rect 4721 5117 4755 5151
rect 5825 5117 5859 5151
rect 6377 5117 6411 5151
rect 7021 5117 7055 5151
rect 10609 5117 10643 5151
rect 10885 5117 10919 5151
rect 7481 5049 7515 5083
rect 10333 5049 10367 5083
rect 1501 4981 1535 5015
rect 4629 4981 4663 5015
rect 14381 4981 14415 5015
rect 3065 4777 3099 4811
rect 3617 4777 3651 4811
rect 9045 4777 9079 4811
rect 9873 4777 9907 4811
rect 10517 4777 10551 4811
rect 11069 4777 11103 4811
rect 4169 4709 4203 4743
rect 8769 4709 8803 4743
rect 2881 4641 2915 4675
rect 9597 4641 9631 4675
rect 10609 4641 10643 4675
rect 2614 4573 2648 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 6009 4573 6043 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7389 4573 7423 4607
rect 9965 4573 9999 4607
rect 10057 4573 10091 4607
rect 10333 4573 10367 4607
rect 10885 4573 10919 4607
rect 14105 4573 14139 4607
rect 5764 4505 5798 4539
rect 7656 4505 7690 4539
rect 1501 4437 1535 4471
rect 4629 4437 4663 4471
rect 6101 4437 6135 4471
rect 6929 4437 6963 4471
rect 10241 4437 10275 4471
rect 14197 4437 14231 4471
rect 4629 4233 4663 4267
rect 5089 4233 5123 4267
rect 8125 4233 8159 4267
rect 9597 4233 9631 4267
rect 3433 4165 3467 4199
rect 5825 4165 5859 4199
rect 1777 4097 1811 4131
rect 2145 4097 2179 4131
rect 4537 4097 4571 4131
rect 4905 4097 4939 4131
rect 6377 4097 6411 4131
rect 6653 4097 6687 4131
rect 6920 4097 6954 4131
rect 8769 4097 8803 4131
rect 9781 4097 9815 4131
rect 14197 4097 14231 4131
rect 3249 4029 3283 4063
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 4445 4029 4479 4063
rect 5273 4029 5307 4063
rect 5917 4029 5951 4063
rect 9321 4029 9355 4063
rect 9505 4029 9539 4063
rect 10609 4029 10643 4063
rect 4077 3961 4111 3995
rect 9965 3961 9999 3995
rect 1501 3893 1535 3927
rect 2789 3893 2823 3927
rect 6469 3893 6503 3927
rect 8033 3893 8067 3927
rect 8861 3893 8895 3927
rect 14381 3893 14415 3927
rect 2145 3689 2179 3723
rect 6285 3689 6319 3723
rect 7205 3689 7239 3723
rect 7757 3689 7791 3723
rect 9781 3689 9815 3723
rect 12081 3689 12115 3723
rect 4905 3553 4939 3587
rect 6745 3553 6779 3587
rect 9597 3553 9631 3587
rect 1777 3485 1811 3519
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 4537 3485 4571 3519
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 7573 3485 7607 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 9413 3485 9447 3519
rect 9873 3485 9907 3519
rect 12173 3485 12207 3519
rect 14197 3485 14231 3519
rect 1409 3417 1443 3451
rect 2504 3417 2538 3451
rect 5172 3417 5206 3451
rect 3617 3349 3651 3383
rect 3985 3349 4019 3383
rect 7389 3349 7423 3383
rect 8309 3349 8343 3383
rect 8953 3349 8987 3383
rect 14381 3349 14415 3383
rect 1685 3145 1719 3179
rect 2145 3145 2179 3179
rect 5365 3145 5399 3179
rect 8677 3145 8711 3179
rect 14289 3145 14323 3179
rect 2513 3077 2547 3111
rect 4230 3077 4264 3111
rect 6009 3077 6043 3111
rect 1777 3009 1811 3043
rect 1869 3009 1903 3043
rect 2329 3009 2363 3043
rect 2605 3009 2639 3043
rect 3709 3009 3743 3043
rect 3985 3009 4019 3043
rect 5457 3009 5491 3043
rect 6561 3009 6595 3043
rect 8401 3009 8435 3043
rect 9965 3009 9999 3043
rect 10885 3009 10919 3043
rect 11345 3009 11379 3043
rect 11529 3009 11563 3043
rect 11796 3009 11830 3043
rect 14473 3009 14507 3043
rect 1961 2941 1995 2975
rect 6101 2941 6135 2975
rect 9137 2941 9171 2975
rect 9321 2941 9355 2975
rect 10793 2941 10827 2975
rect 6745 2873 6779 2907
rect 8585 2873 8619 2907
rect 9873 2873 9907 2907
rect 11253 2873 11287 2907
rect 3893 2805 3927 2839
rect 12909 2805 12943 2839
rect 2421 2601 2455 2635
rect 4629 2601 4663 2635
rect 5273 2601 5307 2635
rect 6009 2601 6043 2635
rect 7573 2601 7607 2635
rect 9137 2601 9171 2635
rect 10149 2601 10183 2635
rect 11529 2601 11563 2635
rect 12541 2601 12575 2635
rect 13737 2601 13771 2635
rect 14105 2601 14139 2635
rect 4445 2533 4479 2567
rect 2237 2397 2271 2431
rect 3801 2397 3835 2431
rect 4261 2397 4295 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6561 2397 6595 2431
rect 7389 2397 7423 2431
rect 8953 2397 8987 2431
rect 9965 2397 9999 2431
rect 11713 2397 11747 2431
rect 12725 2397 12759 2431
rect 13921 2397 13955 2431
rect 14289 2397 14323 2431
rect 3985 2261 4019 2295
rect 6377 2261 6411 2295
<< metal1 >>
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 1026 17280 1032 17332
rect 1084 17280 1090 17332
rect 1118 17280 1124 17332
rect 1176 17320 1182 17332
rect 1176 17292 2176 17320
rect 1176 17280 1182 17292
rect 1044 17252 1072 17280
rect 1044 17224 1716 17252
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1688 17193 1716 17224
rect 2148 17193 2176 17292
rect 2406 17280 2412 17332
rect 2464 17280 2470 17332
rect 3786 17280 3792 17332
rect 3844 17280 3850 17332
rect 5166 17280 5172 17332
rect 5224 17280 5230 17332
rect 6546 17280 6552 17332
rect 6604 17280 6610 17332
rect 8202 17280 8208 17332
rect 8260 17280 8266 17332
rect 9306 17280 9312 17332
rect 9364 17280 9370 17332
rect 10686 17280 10692 17332
rect 10744 17280 10750 17332
rect 12066 17280 12072 17332
rect 12124 17280 12130 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 14458 17320 14464 17332
rect 13771 17292 14464 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 2424 17252 2452 17280
rect 2424 17224 2544 17252
rect 2516 17193 2544 17224
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 3804 17184 3832 17280
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3804 17156 3893 17184
rect 2501 17147 2559 17153
rect 3881 17153 3893 17156
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 2424 17116 2452 17147
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 4212 17156 4261 17184
rect 4212 17144 4218 17156
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 5184 17184 5212 17280
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 5184 17156 5457 17184
rect 4249 17147 4307 17153
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 6564 17184 6592 17280
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6564 17156 6837 17184
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 8220 17184 8248 17280
rect 8067 17156 8248 17184
rect 9324 17184 9352 17280
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9324 17156 9413 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 9401 17153 9413 17156
rect 9447 17153 9459 17187
rect 10704 17184 10732 17280
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10704 17156 10977 17184
rect 9401 17147 9459 17153
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 12084 17184 12112 17280
rect 14568 17252 14596 17280
rect 13096 17224 14596 17252
rect 13096 17193 13124 17224
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 12084 17156 12357 17184
rect 10965 17147 11023 17153
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 13817 17187 13875 17193
rect 13817 17153 13829 17187
rect 13863 17184 13875 17187
rect 13998 17184 14004 17196
rect 13863 17156 14004 17184
rect 13863 17153 13875 17156
rect 13817 17147 13875 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14090 17144 14096 17196
rect 14148 17184 14154 17196
rect 14185 17187 14243 17193
rect 14185 17184 14197 17187
rect 14148 17156 14197 17184
rect 14148 17144 14154 17156
rect 14185 17153 14197 17156
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 2774 17116 2780 17128
rect 2424 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 11146 17116 11152 17128
rect 3988 17088 11152 17116
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 3694 17048 3700 17060
rect 1903 17020 3700 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 1578 16940 1584 16992
rect 1636 16940 1642 16992
rect 1946 16940 1952 16992
rect 2004 16940 2010 16992
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 2188 16952 2237 16980
rect 2188 16940 2194 16952
rect 2225 16949 2237 16952
rect 2271 16949 2283 16983
rect 2225 16943 2283 16949
rect 2685 16983 2743 16989
rect 2685 16949 2697 16983
rect 2731 16980 2743 16983
rect 3988 16980 4016 17088
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 4065 17051 4123 17057
rect 4065 17017 4077 17051
rect 4111 17048 4123 17051
rect 4111 17020 5764 17048
rect 4111 17017 4123 17020
rect 4065 17011 4123 17017
rect 5736 16992 5764 17020
rect 7208 17020 9628 17048
rect 7208 16992 7236 17020
rect 2731 16952 4016 16980
rect 2731 16949 2743 16952
rect 2685 16943 2743 16949
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 4304 16952 4445 16980
rect 4304 16940 4310 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 5261 16983 5319 16989
rect 5261 16980 5273 16983
rect 4948 16952 5273 16980
rect 4948 16940 4954 16952
rect 5261 16949 5273 16952
rect 5307 16949 5319 16983
rect 5261 16943 5319 16949
rect 5718 16940 5724 16992
rect 5776 16940 5782 16992
rect 5810 16940 5816 16992
rect 5868 16940 5874 16992
rect 6638 16940 6644 16992
rect 6696 16940 6702 16992
rect 7190 16940 7196 16992
rect 7248 16940 7254 16992
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 9030 16980 9036 16992
rect 8251 16952 9036 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9600 16989 9628 17020
rect 9585 16983 9643 16989
rect 9585 16949 9597 16983
rect 9631 16980 9643 16983
rect 9858 16980 9864 16992
rect 9631 16952 9864 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10778 16940 10784 16992
rect 10836 16940 10842 16992
rect 12158 16940 12164 16992
rect 12216 16940 12222 16992
rect 13262 16940 13268 16992
rect 13320 16940 13326 16992
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 1636 16748 5580 16776
rect 1636 16736 1642 16748
rect 2961 16711 3019 16717
rect 2961 16677 2973 16711
rect 3007 16677 3019 16711
rect 5552 16708 5580 16748
rect 5626 16736 5632 16788
rect 5684 16736 5690 16788
rect 7944 16748 9674 16776
rect 5552 16680 7880 16708
rect 2961 16671 3019 16677
rect 1946 16640 1952 16652
rect 1780 16612 1952 16640
rect 1780 16581 1808 16612
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2976 16640 3004 16671
rect 3973 16643 4031 16649
rect 3973 16640 3985 16643
rect 2976 16612 3985 16640
rect 3973 16609 3985 16612
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 5810 16600 5816 16652
rect 5868 16640 5874 16652
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 5868 16612 6377 16640
rect 5868 16600 5874 16612
rect 6365 16609 6377 16612
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 6564 16612 6960 16640
rect 6564 16584 6592 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16541 1915 16575
rect 1857 16535 1915 16541
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1872 16504 1900 16535
rect 2774 16532 2780 16584
rect 2832 16532 2838 16584
rect 3050 16532 3056 16584
rect 3108 16532 3114 16584
rect 3513 16575 3571 16581
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3559 16544 3801 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5491 16544 5856 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 992 16476 1900 16504
rect 2746 16476 4568 16504
rect 992 16464 998 16476
rect 1670 16396 1676 16448
rect 1728 16396 1734 16448
rect 2041 16439 2099 16445
rect 2041 16405 2053 16439
rect 2087 16436 2099 16439
rect 2746 16436 2774 16476
rect 2087 16408 2774 16436
rect 3237 16439 3295 16445
rect 2087 16405 2099 16408
rect 2041 16399 2099 16405
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3510 16436 3516 16448
rect 3283 16408 3516 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4433 16439 4491 16445
rect 4433 16436 4445 16439
rect 3936 16408 4445 16436
rect 3936 16396 3942 16408
rect 4433 16405 4445 16408
rect 4479 16405 4491 16439
rect 4540 16436 4568 16476
rect 4706 16464 4712 16516
rect 4764 16464 4770 16516
rect 4798 16464 4804 16516
rect 4856 16464 4862 16516
rect 5350 16464 5356 16516
rect 5408 16464 5414 16516
rect 5828 16448 5856 16544
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 6932 16572 6960 16612
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6779 16544 6868 16572
rect 6932 16544 7113 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 6840 16448 6868 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7190 16532 7196 16584
rect 7248 16532 7254 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7524 16544 7757 16572
rect 7524 16532 7530 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7852 16572 7880 16680
rect 7944 16649 7972 16748
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 9646 16640 9674 16748
rect 12158 16736 12164 16788
rect 12216 16736 12222 16788
rect 13262 16736 13268 16788
rect 13320 16736 13326 16788
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 9784 16680 11713 16708
rect 9784 16640 9812 16680
rect 11701 16677 11713 16680
rect 11747 16677 11759 16711
rect 11701 16671 11759 16677
rect 12176 16640 12204 16736
rect 9646 16612 9812 16640
rect 11808 16612 12204 16640
rect 13280 16640 13308 16736
rect 13354 16668 13360 16720
rect 13412 16668 13418 16720
rect 13280 16612 13768 16640
rect 7929 16603 7987 16609
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 7852 16544 9413 16572
rect 7745 16535 7803 16541
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 10594 16572 10600 16584
rect 9968 16544 10600 16572
rect 9493 16507 9551 16513
rect 9493 16473 9505 16507
rect 9539 16504 9551 16507
rect 9968 16504 9996 16544
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10778 16532 10784 16584
rect 10836 16532 10842 16584
rect 11808 16581 11836 16612
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16572 13139 16575
rect 13354 16572 13360 16584
rect 13127 16544 13360 16572
rect 13127 16541 13139 16544
rect 13081 16535 13139 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 13740 16581 13768 16612
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13504 16544 13553 16572
rect 13504 16532 13510 16544
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14185 16575 14243 16581
rect 14185 16572 14197 16575
rect 13964 16544 14197 16572
rect 13964 16532 13970 16544
rect 14185 16541 14197 16544
rect 14231 16541 14243 16575
rect 14185 16535 14243 16541
rect 14090 16504 14096 16516
rect 9539 16476 9996 16504
rect 10060 16476 14096 16504
rect 9539 16473 9551 16476
rect 9493 16467 9551 16473
rect 5258 16436 5264 16448
rect 4540 16408 5264 16436
rect 4433 16399 4491 16405
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5810 16396 5816 16448
rect 5868 16396 5874 16448
rect 5902 16396 5908 16448
rect 5960 16396 5966 16448
rect 6822 16396 6828 16448
rect 6880 16396 6886 16448
rect 6914 16396 6920 16448
rect 6972 16396 6978 16448
rect 7282 16396 7288 16448
rect 7340 16396 7346 16448
rect 10060 16445 10088 16476
rect 14090 16464 14096 16476
rect 14148 16464 14154 16516
rect 10045 16439 10103 16445
rect 10045 16405 10057 16439
rect 10091 16405 10103 16439
rect 10045 16399 10103 16405
rect 10686 16396 10692 16448
rect 10744 16396 10750 16448
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12584 16408 13001 16436
rect 12584 16396 12590 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 13814 16396 13820 16448
rect 13872 16396 13878 16448
rect 14366 16396 14372 16448
rect 14424 16396 14430 16448
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16232 2651 16235
rect 2774 16232 2780 16244
rect 2639 16204 2780 16232
rect 2639 16201 2651 16204
rect 2593 16195 2651 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 3329 16235 3387 16241
rect 3329 16232 3341 16235
rect 3108 16204 3341 16232
rect 3108 16192 3114 16204
rect 3329 16201 3341 16204
rect 3375 16201 3387 16235
rect 3329 16195 3387 16201
rect 3510 16192 3516 16244
rect 3568 16192 3574 16244
rect 5537 16235 5595 16241
rect 5537 16201 5549 16235
rect 5583 16232 5595 16235
rect 5902 16232 5908 16244
rect 5583 16204 5908 16232
rect 5583 16201 5595 16204
rect 5537 16195 5595 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6914 16192 6920 16244
rect 6972 16192 6978 16244
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7282 16232 7288 16244
rect 7239 16204 7288 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 7466 16192 7472 16244
rect 7524 16192 7530 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 13906 16232 13912 16244
rect 9355 16204 13912 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 14056 16204 14197 16232
rect 14056 16192 14062 16204
rect 14185 16201 14197 16204
rect 14231 16201 14243 16235
rect 14185 16195 14243 16201
rect 1026 16124 1032 16176
rect 1084 16164 1090 16176
rect 3528 16164 3556 16192
rect 1084 16136 2084 16164
rect 3528 16136 3832 16164
rect 1084 16124 1090 16136
rect 2056 16105 2084 16136
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2041 16099 2099 16105
rect 1811 16068 1900 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1872 15969 1900 16068
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 2455 16068 2881 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2869 16065 2881 16068
rect 2915 16096 2927 16099
rect 3053 16099 3111 16105
rect 3053 16096 3065 16099
rect 2915 16068 3065 16096
rect 2915 16065 2927 16068
rect 2869 16059 2927 16065
rect 3053 16065 3065 16068
rect 3099 16096 3111 16099
rect 3510 16096 3516 16108
rect 3099 16068 3516 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 3804 16105 3832 16136
rect 4246 16124 4252 16176
rect 4304 16164 4310 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 4304 16136 4537 16164
rect 4304 16124 4310 16136
rect 4525 16133 4537 16136
rect 4571 16133 4583 16167
rect 4525 16127 4583 16133
rect 5077 16167 5135 16173
rect 5077 16133 5089 16167
rect 5123 16164 5135 16167
rect 5350 16164 5356 16176
rect 5123 16136 5356 16164
rect 5123 16133 5135 16136
rect 5077 16127 5135 16133
rect 5350 16124 5356 16136
rect 5408 16164 5414 16176
rect 5408 16136 6868 16164
rect 5408 16124 5414 16136
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16065 3847 16099
rect 3789 16059 3847 16065
rect 5258 16056 5264 16108
rect 5316 16056 5322 16108
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 16028 3663 16031
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 3651 16000 3740 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15929 1915 15963
rect 1857 15923 1915 15929
rect 1670 15852 1676 15904
rect 1728 15852 1734 15904
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 2777 15895 2835 15901
rect 2777 15892 2789 15895
rect 2464 15864 2789 15892
rect 2464 15852 2470 15864
rect 2777 15861 2789 15864
rect 2823 15861 2835 15895
rect 2777 15855 2835 15861
rect 3142 15852 3148 15904
rect 3200 15852 3206 15904
rect 3712 15892 3740 16000
rect 3896 16000 4445 16028
rect 3896 15972 3924 16000
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 5994 15988 6000 16040
rect 6052 15988 6058 16040
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 16028 6239 16031
rect 6549 16031 6607 16037
rect 6549 16028 6561 16031
rect 6227 16000 6561 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 3878 15920 3884 15972
rect 3936 15920 3942 15972
rect 4249 15963 4307 15969
rect 4249 15929 4261 15963
rect 4295 15960 4307 15963
rect 4724 15960 4752 15988
rect 4295 15932 4752 15960
rect 4295 15929 4307 15932
rect 4249 15923 4307 15929
rect 6472 15904 6500 16000
rect 6549 15997 6561 16000
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6730 15988 6736 16040
rect 6788 15988 6794 16040
rect 6840 16028 6868 16136
rect 6932 16096 6960 16192
rect 7300 16164 7328 16192
rect 8113 16167 8171 16173
rect 7300 16136 7604 16164
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6932 16068 7297 16096
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7576 16028 7604 16136
rect 8113 16133 8125 16167
rect 8159 16164 8171 16167
rect 8478 16164 8484 16176
rect 8159 16136 8484 16164
rect 8159 16133 8171 16136
rect 8113 16127 8171 16133
rect 8478 16124 8484 16136
rect 8536 16124 8542 16176
rect 9030 16124 9036 16176
rect 9088 16124 9094 16176
rect 10686 16124 10692 16176
rect 10744 16124 10750 16176
rect 9048 16096 9076 16124
rect 9125 16099 9183 16105
rect 9125 16096 9137 16099
rect 9048 16068 9137 16096
rect 9125 16065 9137 16068
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 10134 16056 10140 16108
rect 10192 16056 10198 16108
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16096 10655 16099
rect 10704 16096 10732 16124
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 10643 16068 10732 16096
rect 12406 16068 14105 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 6840 16000 7420 16028
rect 7576 16000 8217 16028
rect 4522 15892 4528 15904
rect 3712 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5353 15895 5411 15901
rect 5353 15861 5365 15895
rect 5399 15892 5411 15895
rect 5534 15892 5540 15904
rect 5399 15864 5540 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6454 15852 6460 15904
rect 6512 15852 6518 15904
rect 7392 15892 7420 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 10778 15988 10784 16040
rect 10836 15988 10842 16040
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 7524 15932 7665 15960
rect 7524 15920 7530 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 12406 15960 12434 16068
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 7653 15923 7711 15929
rect 7760 15932 12434 15960
rect 7760 15892 7788 15932
rect 7392 15864 7788 15892
rect 10318 15852 10324 15904
rect 10376 15852 10382 15904
rect 11054 15852 11060 15904
rect 11112 15852 11118 15904
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 1670 15648 1676 15700
rect 1728 15648 1734 15700
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4154 15688 4160 15700
rect 4111 15660 4160 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4706 15648 4712 15700
rect 4764 15648 4770 15700
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 5902 15648 5908 15700
rect 5960 15648 5966 15700
rect 6181 15691 6239 15697
rect 6181 15657 6193 15691
rect 6227 15688 6239 15691
rect 6454 15688 6460 15700
rect 6227 15660 6460 15688
rect 6227 15657 6239 15660
rect 6181 15651 6239 15657
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 7469 15691 7527 15697
rect 7469 15688 7481 15691
rect 6788 15660 7481 15688
rect 6788 15648 6794 15660
rect 7469 15657 7481 15660
rect 7515 15657 7527 15691
rect 7469 15651 7527 15657
rect 10318 15648 10324 15700
rect 10376 15648 10382 15700
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 11149 15691 11207 15697
rect 11149 15688 11161 15691
rect 10836 15660 11161 15688
rect 10836 15648 10842 15660
rect 11149 15657 11161 15660
rect 11195 15657 11207 15691
rect 11149 15651 11207 15657
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 14415 15660 14872 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 1688 15552 1716 15648
rect 2225 15555 2283 15561
rect 2225 15552 2237 15555
rect 1688 15524 2237 15552
rect 2225 15521 2237 15524
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 1854 15444 1860 15496
rect 1912 15444 1918 15496
rect 2130 15444 2136 15496
rect 2188 15444 2194 15496
rect 2240 15484 2268 15515
rect 2406 15512 2412 15564
rect 2464 15512 2470 15564
rect 3160 15552 3188 15648
rect 4249 15623 4307 15629
rect 4249 15589 4261 15623
rect 4295 15620 4307 15623
rect 4816 15620 4844 15648
rect 4295 15592 4844 15620
rect 4295 15589 4307 15592
rect 4249 15583 4307 15589
rect 4893 15555 4951 15561
rect 4893 15552 4905 15555
rect 3160 15524 4905 15552
rect 4893 15521 4905 15524
rect 4939 15521 4951 15555
rect 4893 15515 4951 15521
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15552 5135 15555
rect 5920 15552 5948 15648
rect 6549 15623 6607 15629
rect 6549 15589 6561 15623
rect 6595 15620 6607 15623
rect 6595 15592 10272 15620
rect 6595 15589 6607 15592
rect 6549 15583 6607 15589
rect 5123 15524 5948 15552
rect 6104 15524 10180 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 3418 15484 3424 15496
rect 2240 15456 3424 15484
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3602 15444 3608 15496
rect 3660 15444 3666 15496
rect 3881 15487 3939 15493
rect 3881 15453 3893 15487
rect 3927 15484 3939 15487
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3927 15456 4169 15484
rect 3927 15453 3939 15456
rect 3881 15447 3939 15453
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15416 2927 15419
rect 2915 15388 3556 15416
rect 2915 15385 2927 15388
rect 2869 15379 2927 15385
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 1670 15308 1676 15360
rect 1728 15308 1734 15360
rect 2038 15308 2044 15360
rect 2096 15308 2102 15360
rect 2961 15351 3019 15357
rect 2961 15317 2973 15351
rect 3007 15348 3019 15351
rect 3050 15348 3056 15360
rect 3007 15320 3056 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3528 15348 3556 15388
rect 4172 15360 4200 15447
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 6104 15493 6132 15524
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 5718 15376 5724 15428
rect 5776 15416 5782 15428
rect 6104 15416 6132 15447
rect 6362 15444 6368 15496
rect 6420 15484 6426 15496
rect 6638 15484 6644 15496
rect 6420 15456 6644 15484
rect 6420 15444 6426 15456
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 6880 15456 7205 15484
rect 6880 15444 6886 15456
rect 7193 15453 7205 15456
rect 7239 15484 7251 15487
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7239 15456 7389 15484
rect 7239 15453 7251 15456
rect 7193 15447 7251 15453
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9180 15456 9505 15484
rect 9180 15444 9186 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 5776 15388 6132 15416
rect 5776 15376 5782 15388
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 7745 15419 7803 15425
rect 7745 15416 7757 15419
rect 7524 15388 7757 15416
rect 7524 15376 7530 15388
rect 7745 15385 7757 15388
rect 7791 15385 7803 15419
rect 7745 15379 7803 15385
rect 8294 15376 8300 15428
rect 8352 15376 8358 15428
rect 8389 15419 8447 15425
rect 8389 15385 8401 15419
rect 8435 15416 8447 15419
rect 8573 15419 8631 15425
rect 8573 15416 8585 15419
rect 8435 15388 8585 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 8573 15385 8585 15388
rect 8619 15385 8631 15419
rect 9048 15416 9076 15444
rect 9968 15416 9996 15447
rect 9048 15388 9996 15416
rect 8573 15379 8631 15385
rect 3878 15348 3884 15360
rect 3528 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 5350 15308 5356 15360
rect 5408 15308 5414 15360
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 8938 15308 8944 15360
rect 8996 15308 9002 15360
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 10042 15308 10048 15360
rect 10100 15308 10106 15360
rect 10152 15348 10180 15524
rect 10244 15416 10272 15592
rect 10336 15552 10364 15648
rect 14844 15632 14872 15660
rect 14826 15580 14832 15632
rect 14884 15580 14890 15632
rect 10336 15524 11376 15552
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10594 15444 10600 15496
rect 10652 15444 10658 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11348 15493 11376 15524
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 11333 15447 11391 15453
rect 12406 15456 14197 15484
rect 12406 15416 12434 15456
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 10244 15388 12434 15416
rect 13722 15348 13728 15360
rect 10152 15320 13728 15348
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 3602 15104 3608 15156
rect 3660 15144 3666 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 3660 15116 4261 15144
rect 3660 15104 3666 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 4249 15107 4307 15113
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6089 15147 6147 15153
rect 6089 15144 6101 15147
rect 6052 15116 6101 15144
rect 6052 15104 6058 15116
rect 6089 15113 6101 15116
rect 6135 15113 6147 15147
rect 6089 15107 6147 15113
rect 6362 15104 6368 15156
rect 6420 15104 6426 15156
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8294 15144 8300 15156
rect 8067 15116 8300 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 10134 15144 10140 15156
rect 9539 15116 10140 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 11146 15104 11152 15156
rect 11204 15104 11210 15156
rect 3050 15085 3056 15088
rect 1596 15048 2544 15076
rect 1596 15017 1624 15048
rect 2516 15020 2544 15048
rect 3044 15039 3056 15085
rect 3108 15076 3114 15088
rect 3108 15048 3144 15076
rect 3050 15036 3056 15039
rect 3108 15036 3114 15048
rect 5350 15036 5356 15088
rect 5408 15085 5414 15088
rect 5408 15076 5420 15085
rect 6380 15076 6408 15104
rect 6638 15085 6644 15088
rect 6632 15076 6644 15085
rect 5408 15048 5453 15076
rect 5920 15048 6408 15076
rect 6599 15048 6644 15076
rect 5408 15039 5420 15048
rect 5408 15036 5414 15039
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 2038 15008 2044 15020
rect 1719 14980 2044 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2498 14968 2504 15020
rect 2556 14968 2562 15020
rect 5920 15017 5948 15048
rect 6632 15039 6644 15048
rect 6638 15036 6644 15039
rect 6696 15036 6702 15088
rect 8380 15079 8438 15085
rect 8380 15045 8392 15079
rect 8426 15076 8438 15079
rect 8938 15076 8944 15088
rect 8426 15048 8944 15076
rect 8426 15045 8438 15048
rect 8380 15039 8438 15045
rect 8938 15036 8944 15048
rect 8996 15036 9002 15088
rect 10042 15076 10048 15088
rect 9600 15048 10048 15076
rect 5905 15011 5963 15017
rect 2792 14980 5672 15008
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14909 1915 14943
rect 1857 14903 1915 14909
rect 1489 14875 1547 14881
rect 1489 14841 1501 14875
rect 1535 14872 1547 14875
rect 1872 14872 1900 14903
rect 2406 14900 2412 14952
rect 2464 14900 2470 14952
rect 2792 14949 2820 14980
rect 5644 14952 5672 14980
rect 5905 14977 5917 15011
rect 5951 14977 5963 15011
rect 5905 14971 5963 14977
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 7834 14968 7840 15020
rect 7892 14968 7898 15020
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 9600 15017 9628 15048
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 11164 15076 11192 15104
rect 13354 15076 13360 15088
rect 11164 15048 13360 15076
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 8904 14980 9597 15008
rect 8904 14968 8910 14980
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9585 14971 9643 14977
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9732 14980 9781 15008
rect 9732 14968 9738 14980
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10410 15008 10416 15020
rect 10367 14980 10416 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10410 14968 10416 14980
rect 10468 15008 10474 15020
rect 11256 15017 11284 15048
rect 13354 15036 13360 15048
rect 13412 15036 13418 15088
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10468 14980 11161 15008
rect 10468 14968 10474 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11241 15011 11299 15017
rect 11241 14977 11253 15011
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12124 14980 12449 15008
rect 12124 14968 12130 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 13035 14980 13093 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 1535 14844 1900 14872
rect 1535 14841 1547 14844
rect 1489 14835 1547 14841
rect 2038 14764 2044 14816
rect 2096 14764 2102 14816
rect 2792 14804 2820 14903
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5684 14912 6377 14940
rect 5684 14900 5690 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 8110 14900 8116 14952
rect 8168 14900 8174 14952
rect 10502 14900 10508 14952
rect 10560 14900 10566 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 10704 14912 11529 14940
rect 10704 14881 10732 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 11747 14912 12357 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12710 14900 12716 14952
rect 12768 14900 12774 14952
rect 10229 14875 10287 14881
rect 10229 14841 10241 14875
rect 10275 14872 10287 14875
rect 10689 14875 10747 14881
rect 10689 14872 10701 14875
rect 10275 14844 10701 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 10689 14841 10701 14844
rect 10735 14841 10747 14875
rect 13004 14872 13032 14971
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 10689 14835 10747 14841
rect 12452 14844 13032 14872
rect 12452 14816 12480 14844
rect 3050 14804 3056 14816
rect 2792 14776 3056 14804
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 4154 14764 4160 14816
rect 4212 14764 4218 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 5408 14776 5825 14804
rect 5408 14764 5414 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 5813 14767 5871 14773
rect 7745 14807 7803 14813
rect 7745 14773 7757 14807
rect 7791 14804 7803 14807
rect 8294 14804 8300 14816
rect 7791 14776 8300 14804
rect 7791 14773 7803 14776
rect 7745 14767 7803 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 12158 14764 12164 14816
rect 12216 14764 12222 14816
rect 12434 14764 12440 14816
rect 12492 14764 12498 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 13262 14764 13268 14816
rect 13320 14764 13326 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 2038 14560 2044 14612
rect 2096 14560 2102 14612
rect 2406 14560 2412 14612
rect 2464 14560 2470 14612
rect 5902 14600 5908 14612
rect 2608 14572 5908 14600
rect 2424 14473 2452 14560
rect 2501 14535 2559 14541
rect 2501 14501 2513 14535
rect 2547 14501 2559 14535
rect 2501 14495 2559 14501
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14433 2467 14467
rect 2409 14427 2467 14433
rect 1489 14399 1547 14405
rect 1489 14365 1501 14399
rect 1535 14396 1547 14399
rect 1578 14396 1584 14408
rect 1535 14368 1584 14396
rect 1535 14365 1547 14368
rect 1489 14359 1547 14365
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2516 14396 2544 14495
rect 2271 14368 2544 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 2608 14260 2636 14572
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6641 14603 6699 14609
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 6822 14600 6828 14612
rect 6687 14572 6828 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7892 14572 8125 14600
rect 7892 14560 7898 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8478 14560 8484 14612
rect 8536 14560 8542 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9916 14572 10149 14600
rect 9916 14560 9922 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 10502 14560 10508 14612
rect 10560 14560 10566 14612
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 10652 14572 10793 14600
rect 10652 14560 10658 14572
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 10781 14563 10839 14569
rect 12802 14560 12808 14612
rect 12860 14560 12866 14612
rect 14182 14560 14188 14612
rect 14240 14560 14246 14612
rect 2682 14492 2688 14544
rect 2740 14532 2746 14544
rect 3421 14535 3479 14541
rect 2740 14504 3004 14532
rect 2740 14492 2746 14504
rect 2976 14405 3004 14504
rect 3421 14501 3433 14535
rect 3467 14501 3479 14535
rect 3421 14495 3479 14501
rect 4065 14535 4123 14541
rect 4065 14501 4077 14535
rect 4111 14532 4123 14535
rect 5074 14532 5080 14544
rect 4111 14504 5080 14532
rect 4111 14501 4123 14504
rect 4065 14495 4123 14501
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14396 2743 14399
rect 2961 14399 3019 14405
rect 2731 14368 2820 14396
rect 2731 14365 2743 14368
rect 2685 14359 2743 14365
rect 2792 14269 2820 14368
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 3007 14368 3249 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3237 14365 3249 14368
rect 3283 14365 3295 14399
rect 3436 14396 3464 14495
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4212 14436 4445 14464
rect 4212 14424 4218 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4890 14424 4896 14476
rect 4948 14424 4954 14476
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14464 8079 14467
rect 8110 14464 8116 14476
rect 8067 14436 8116 14464
rect 8067 14433 8079 14436
rect 8021 14427 8079 14433
rect 8110 14424 8116 14436
rect 8168 14464 8174 14476
rect 8478 14464 8484 14476
rect 8168 14436 8484 14464
rect 8168 14424 8174 14436
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 8536 14436 11069 14464
rect 8536 14424 8542 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 12820 14464 12848 14560
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 13219 14504 13645 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 13633 14495 13691 14501
rect 12759 14436 12848 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3436 14368 3893 14396
rect 3237 14359 3295 14365
rect 3881 14365 3893 14368
rect 3927 14365 3939 14399
rect 3881 14359 3939 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4908 14396 4936 14424
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 4387 14368 4936 14396
rect 5644 14368 6561 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 3252 14272 3280 14359
rect 5644 14340 5672 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 7668 14368 7880 14396
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 4982 14328 4988 14340
rect 4295 14300 4988 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 5626 14288 5632 14340
rect 5684 14288 5690 14340
rect 6304 14331 6362 14337
rect 6304 14297 6316 14331
rect 6350 14328 6362 14331
rect 7668 14328 7696 14368
rect 6350 14300 7696 14328
rect 7754 14331 7812 14337
rect 6350 14297 6362 14300
rect 6304 14291 6362 14297
rect 7754 14297 7766 14331
rect 7800 14297 7812 14331
rect 7852 14328 7880 14368
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8352 14368 8585 14396
rect 8352 14356 8358 14368
rect 8573 14365 8585 14368
rect 8619 14396 8631 14399
rect 9122 14396 9128 14408
rect 8619 14368 9128 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 7852 14300 9413 14328
rect 7754 14291 7812 14297
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 1627 14232 2636 14260
rect 2777 14263 2835 14269
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 2777 14229 2789 14263
rect 2823 14229 2835 14263
rect 2777 14223 2835 14229
rect 3234 14220 3240 14272
rect 3292 14220 3298 14272
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 5077 14263 5135 14269
rect 5077 14260 5089 14263
rect 4856 14232 5089 14260
rect 4856 14220 4862 14232
rect 5077 14229 5089 14232
rect 5123 14229 5135 14263
rect 5077 14223 5135 14229
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5994 14260 6000 14272
rect 5224 14232 6000 14260
rect 5224 14220 5230 14232
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 7760 14260 7788 14291
rect 7248 14232 7788 14260
rect 10060 14260 10088 14359
rect 10134 14356 10140 14408
rect 10192 14356 10198 14408
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 10284 14368 10333 14396
rect 10284 14356 10290 14368
rect 10321 14365 10333 14368
rect 10367 14396 10379 14399
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 10367 14368 10609 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10152 14328 10180 14356
rect 10704 14328 10732 14359
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 12216 14368 12541 14396
rect 12216 14356 12222 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12618 14356 12624 14408
rect 12676 14396 12682 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 12676 14368 13277 14396
rect 12676 14356 12682 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 13648 14396 13676 14495
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13648 14368 14105 14396
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 10152 14300 10732 14328
rect 11146 14288 11152 14340
rect 11204 14328 11210 14340
rect 11302 14331 11360 14337
rect 11302 14328 11314 14331
rect 11204 14300 11314 14328
rect 11204 14288 11210 14300
rect 11302 14297 11314 14300
rect 11348 14297 11360 14331
rect 11302 14291 11360 14297
rect 12434 14260 12440 14272
rect 10060 14232 12440 14260
rect 7248 14220 7254 14232
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1670 14016 1676 14068
rect 1728 14016 1734 14068
rect 3513 14059 3571 14065
rect 3513 14025 3525 14059
rect 3559 14056 3571 14059
rect 7101 14059 7159 14065
rect 3559 14028 5764 14056
rect 3559 14025 3571 14028
rect 3513 14019 3571 14025
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1688 13920 1716 14016
rect 3234 13988 3240 14000
rect 1627 13892 1716 13920
rect 2240 13960 2912 13988
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2240 13852 2268 13960
rect 2332 13892 2774 13920
rect 2332 13861 2360 13892
rect 1719 13824 2268 13852
rect 2317 13855 2375 13861
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2501 13855 2559 13861
rect 2501 13852 2513 13855
rect 2317 13815 2375 13821
rect 2424 13824 2513 13852
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 2424 13784 2452 13824
rect 2501 13821 2513 13824
rect 2547 13821 2559 13855
rect 2501 13815 2559 13821
rect 2096 13756 2452 13784
rect 2096 13744 2102 13756
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 1857 13719 1915 13725
rect 1857 13716 1869 13719
rect 1820 13688 1869 13716
rect 1820 13676 1826 13688
rect 1857 13685 1869 13688
rect 1903 13685 1915 13719
rect 1857 13679 1915 13685
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 2593 13719 2651 13725
rect 2593 13716 2605 13719
rect 2556 13688 2605 13716
rect 2556 13676 2562 13688
rect 2593 13685 2605 13688
rect 2639 13685 2651 13719
rect 2746 13716 2774 13892
rect 2884 13784 2912 13960
rect 3160 13960 3240 13988
rect 3160 13929 3188 13960
rect 3234 13948 3240 13960
rect 3292 13988 3298 14000
rect 3528 13988 3556 14019
rect 3292 13960 3556 13988
rect 4648 13991 4706 13997
rect 3292 13948 3298 13960
rect 4648 13957 4660 13991
rect 4694 13988 4706 13991
rect 4798 13988 4804 14000
rect 4694 13960 4804 13988
rect 4694 13957 4706 13960
rect 4648 13951 4706 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 4908 13960 5672 13988
rect 4908 13929 4936 13960
rect 5644 13932 5672 13960
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 4893 13923 4951 13929
rect 3145 13883 3203 13889
rect 3252 13892 4844 13920
rect 3252 13784 3280 13892
rect 4816 13852 4844 13892
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 4982 13880 4988 13932
rect 5040 13880 5046 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 5132 13892 5181 13920
rect 5132 13880 5138 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5626 13880 5632 13932
rect 5684 13880 5690 13932
rect 5736 13929 5764 14028
rect 7101 14025 7113 14059
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14025 7435 14059
rect 7377 14019 7435 14025
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 12161 14059 12219 14065
rect 9539 14028 10364 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 6914 13880 6920 13932
rect 6972 13880 6978 13932
rect 7116 13920 7144 14019
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 7116 13892 7205 13920
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7392 13920 7420 14019
rect 8036 13960 9720 13988
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7392 13892 7941 13920
rect 7193 13883 7251 13889
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8036 13852 8064 13960
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8352 13892 8493 13920
rect 8352 13880 8358 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13920 9367 13923
rect 9355 13910 9444 13920
rect 9355 13892 9536 13910
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 9416 13882 9536 13892
rect 4816 13824 8064 13852
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 8159 13824 8217 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 8205 13821 8217 13824
rect 8251 13821 8263 13855
rect 8205 13815 8263 13821
rect 8680 13824 9444 13852
rect 8680 13793 8708 13824
rect 2884 13756 3280 13784
rect 8665 13787 8723 13793
rect 8665 13753 8677 13787
rect 8711 13753 8723 13787
rect 8665 13747 8723 13753
rect 3142 13716 3148 13728
rect 2746 13688 3148 13716
rect 2593 13679 2651 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 4580 13688 5365 13716
rect 4580 13676 4586 13688
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 5353 13679 5411 13685
rect 5810 13676 5816 13728
rect 5868 13676 5874 13728
rect 7745 13719 7803 13725
rect 7745 13685 7757 13719
rect 7791 13716 7803 13719
rect 7834 13716 7840 13728
rect 7791 13688 7840 13716
rect 7791 13685 7803 13688
rect 7745 13679 7803 13685
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 9416 13716 9444 13824
rect 9508 13784 9536 13882
rect 9692 13852 9720 13960
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10226 13988 10232 14000
rect 10008 13960 10232 13988
rect 10008 13948 10014 13960
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 9968 13920 9996 13948
rect 9815 13892 9996 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9692 13824 9965 13852
rect 9953 13821 9965 13824
rect 9999 13852 10011 13855
rect 9999 13824 10088 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 9585 13787 9643 13793
rect 9585 13784 9597 13787
rect 9508 13756 9597 13784
rect 9585 13753 9597 13756
rect 9631 13753 9643 13787
rect 9585 13747 9643 13753
rect 9858 13716 9864 13728
rect 9416 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 10060 13716 10088 13824
rect 10134 13812 10140 13864
rect 10192 13812 10198 13864
rect 10336 13852 10364 14028
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 12207 14028 12265 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12253 14025 12265 14028
rect 12299 14056 12311 14059
rect 12618 14056 12624 14068
rect 12299 14028 12624 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13446 14056 13452 14068
rect 13219 14028 13452 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10643 13892 11345 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11379 13892 11529 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 12728 13920 12756 14016
rect 13262 13948 13268 14000
rect 13320 13948 13326 14000
rect 13924 13988 13952 14019
rect 14093 13991 14151 13997
rect 14093 13988 14105 13991
rect 13924 13960 14105 13988
rect 14093 13957 14105 13960
rect 14139 13957 14151 13991
rect 14093 13951 14151 13957
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12728 13892 12909 13920
rect 11517 13883 11575 13889
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13920 13047 13923
rect 13280 13920 13308 13948
rect 13035 13892 13308 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 10336 13824 10640 13852
rect 10612 13784 10640 13824
rect 10686 13812 10692 13864
rect 10744 13812 10750 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10796 13824 10885 13852
rect 10796 13784 10824 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 11698 13812 11704 13864
rect 11756 13812 11762 13864
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14458 13852 14464 13864
rect 14415 13824 14464 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 10612 13756 10824 13784
rect 11238 13716 11244 13728
rect 10060 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 1820 13484 2881 13512
rect 1820 13472 1826 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 4522 13472 4528 13524
rect 4580 13472 4586 13524
rect 5810 13512 5816 13524
rect 4724 13484 5816 13512
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13376 2835 13379
rect 3050 13376 3056 13388
rect 2823 13348 3056 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 4540 13376 4568 13472
rect 4724 13385 4752 13484
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10192 13484 10793 13512
rect 10192 13472 10198 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 10781 13475 10839 13481
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11204 13484 11437 13512
rect 11204 13472 11210 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 11756 13484 12265 13512
rect 11756 13472 11762 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12768 13484 12909 13512
rect 12768 13472 12774 13484
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13413 5687 13447
rect 5629 13407 5687 13413
rect 12621 13447 12679 13453
rect 12621 13413 12633 13447
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 3559 13348 4568 13376
rect 4709 13379 4767 13385
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4709 13345 4721 13379
rect 4755 13345 4767 13379
rect 4709 13339 4767 13345
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 5644 13376 5672 13407
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5644 13348 5917 13376
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13376 8263 13379
rect 8294 13376 8300 13388
rect 8251 13348 8300 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 10042 13336 10048 13388
rect 10100 13336 10106 13388
rect 11606 13376 11612 13388
rect 11164 13348 11612 13376
rect 2498 13268 2504 13320
rect 2556 13317 2562 13320
rect 2556 13308 2568 13317
rect 2556 13280 2601 13308
rect 2556 13271 2568 13280
rect 2556 13268 2562 13271
rect 3326 13268 3332 13320
rect 3384 13268 3390 13320
rect 4890 13268 4896 13320
rect 4948 13268 4954 13320
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 5169 13271 5227 13277
rect 5368 13280 5457 13308
rect 3050 13200 3056 13252
rect 3108 13240 3114 13252
rect 5074 13240 5080 13252
rect 3108 13212 5080 13240
rect 3108 13200 3114 13212
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5184 13184 5212 13271
rect 1394 13132 1400 13184
rect 1452 13132 1458 13184
rect 5166 13132 5172 13184
rect 5224 13132 5230 13184
rect 5368 13181 5396 13280
rect 5445 13277 5457 13280
rect 5491 13277 5503 13311
rect 5552 13308 5580 13336
rect 5718 13308 5724 13320
rect 5552 13280 5724 13308
rect 5445 13271 5503 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6380 13280 6469 13308
rect 5353 13175 5411 13181
rect 5353 13141 5365 13175
rect 5399 13141 5411 13175
rect 5353 13135 5411 13141
rect 6178 13132 6184 13184
rect 6236 13172 6242 13184
rect 6380 13181 6408 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6638 13268 6644 13320
rect 6696 13268 6702 13320
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 6972 13280 7757 13308
rect 6972 13268 6978 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11164 13317 11192 13348
rect 11606 13336 11612 13348
rect 11664 13376 11670 13388
rect 12066 13376 12072 13388
rect 11664 13348 12072 13376
rect 11664 13336 11670 13348
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13277 11207 13311
rect 12084 13308 12112 13336
rect 12084 13302 12204 13308
rect 12321 13305 12379 13311
rect 12321 13302 12333 13305
rect 12084 13280 12333 13302
rect 11149 13271 11207 13277
rect 12176 13274 12333 13280
rect 12321 13271 12333 13274
rect 12367 13302 12379 13305
rect 12437 13307 12495 13313
rect 12437 13302 12449 13307
rect 12367 13274 12449 13302
rect 12367 13271 12379 13274
rect 12321 13265 12379 13271
rect 12437 13273 12449 13274
rect 12483 13273 12495 13307
rect 12636 13308 12664 13407
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12636 13280 12725 13308
rect 12437 13267 12495 13273
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13412 13280 13737 13308
rect 13412 13268 13418 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 13725 13271 13783 13277
rect 13924 13280 14197 13308
rect 7101 13243 7159 13249
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 7834 13240 7840 13252
rect 7147 13212 7840 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7834 13200 7840 13212
rect 7892 13240 7898 13252
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 7892 13212 9045 13240
rect 7892 13200 7898 13212
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9033 13203 9091 13209
rect 9122 13200 9128 13252
rect 9180 13200 9186 13252
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6236 13144 6377 13172
rect 6236 13132 6242 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7282 13172 7288 13184
rect 7239 13144 7288 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8754 13132 8760 13184
rect 8812 13132 8818 13184
rect 10594 13132 10600 13184
rect 10652 13132 10658 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11882 13172 11888 13184
rect 11379 13144 11888 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 13924 13181 13952 13280
rect 14185 13277 14197 13280
rect 14231 13277 14243 13311
rect 14185 13271 14243 13277
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13141 13967 13175
rect 13909 13135 13967 13141
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1394 12928 1400 12980
rect 1452 12968 1458 12980
rect 2685 12971 2743 12977
rect 1452 12940 2360 12968
rect 1452 12928 1458 12940
rect 934 12860 940 12912
rect 992 12900 998 12912
rect 992 12872 1900 12900
rect 992 12860 998 12872
rect 1762 12792 1768 12844
rect 1820 12792 1826 12844
rect 1872 12841 1900 12872
rect 2332 12841 2360 12940
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 3326 12968 3332 12980
rect 2731 12940 3332 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 3694 12928 3700 12980
rect 3752 12928 3758 12980
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 6178 12928 6184 12980
rect 6236 12928 6242 12980
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6696 12940 6837 12968
rect 6696 12928 6702 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 8352 12940 8401 12968
rect 8352 12928 8358 12940
rect 8389 12937 8401 12940
rect 8435 12937 8447 12971
rect 8389 12931 8447 12937
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 9180 12940 10885 12968
rect 9180 12928 9186 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11940 12940 12480 12968
rect 11940 12928 11946 12940
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2498 12832 2504 12844
rect 2363 12804 2504 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2498 12792 2504 12804
rect 2556 12832 2562 12844
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 2556 12804 2605 12832
rect 2556 12792 2562 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2593 12795 2651 12801
rect 2746 12804 3065 12832
rect 2501 12699 2559 12705
rect 2501 12665 2513 12699
rect 2547 12696 2559 12699
rect 2746 12696 2774 12804
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3712 12832 3740 12928
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12900 4215 12903
rect 4203 12872 4660 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 4632 12841 4660 12872
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3712 12804 4077 12832
rect 4065 12801 4077 12804
rect 4111 12832 4123 12835
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4111 12804 4353 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4908 12832 4936 12928
rect 9306 12900 9312 12912
rect 7024 12872 9312 12900
rect 4663 12804 4936 12832
rect 5537 12835 5595 12841
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 5902 12832 5908 12844
rect 5583 12804 5908 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6052 12804 6561 12832
rect 6052 12792 6058 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7024 12841 7052 12872
rect 8496 12844 8524 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 9858 12860 9864 12912
rect 9916 12860 9922 12912
rect 12158 12860 12164 12912
rect 12216 12860 12222 12912
rect 12452 12865 12480 12940
rect 7282 12841 7288 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7276 12832 7288 12841
rect 7243 12804 7288 12832
rect 7009 12795 7067 12801
rect 7276 12795 7288 12804
rect 7282 12792 7288 12795
rect 7340 12792 7346 12844
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 8754 12841 8760 12844
rect 8748 12832 8760 12841
rect 8715 12804 8760 12832
rect 8748 12795 8760 12804
rect 8754 12792 8760 12795
rect 8812 12792 8818 12844
rect 9876 12832 9904 12860
rect 12437 12859 12495 12865
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 9876 12804 11069 12832
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11440 12804 12296 12832
rect 12437 12825 12449 12859
rect 12483 12825 12495 12859
rect 12437 12819 12495 12825
rect 4798 12724 4804 12776
rect 4856 12724 4862 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6457 12767 6515 12773
rect 6457 12764 6469 12767
rect 5767 12736 6469 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 6457 12733 6469 12736
rect 6503 12733 6515 12767
rect 6457 12727 6515 12733
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 10008 12736 10701 12764
rect 10008 12724 10014 12736
rect 10689 12733 10701 12736
rect 10735 12764 10747 12767
rect 10870 12764 10876 12776
rect 10735 12736 10876 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 11164 12764 11192 12795
rect 10928 12736 11192 12764
rect 10928 12724 10934 12736
rect 2547 12668 2774 12696
rect 2869 12699 2927 12705
rect 2547 12665 2559 12668
rect 2501 12659 2559 12665
rect 2869 12665 2881 12699
rect 2915 12696 2927 12699
rect 3142 12696 3148 12708
rect 2915 12668 3148 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 11440 12696 11468 12804
rect 11517 12767 11575 12773
rect 11517 12733 11529 12767
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 12268 12764 12296 12804
rect 12268 12736 12434 12764
rect 11701 12727 11759 12733
rect 4540 12668 7052 12696
rect 1670 12588 1676 12640
rect 1728 12588 1734 12640
rect 2038 12588 2044 12640
rect 2096 12588 2102 12640
rect 3418 12588 3424 12640
rect 3476 12588 3482 12640
rect 4540 12637 4568 12668
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12597 4583 12631
rect 4525 12591 4583 12597
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5534 12628 5540 12640
rect 5307 12600 5540 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 7024 12628 7052 12668
rect 9784 12668 11468 12696
rect 9784 12628 9812 12668
rect 7024 12600 9812 12628
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12628 9919 12631
rect 9950 12628 9956 12640
rect 9907 12600 9956 12628
rect 9907 12597 9919 12600
rect 9861 12591 9919 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 11238 12588 11244 12640
rect 11296 12588 11302 12640
rect 11532 12628 11560 12727
rect 11716 12696 11744 12727
rect 12253 12699 12311 12705
rect 12253 12696 12265 12699
rect 11716 12668 12265 12696
rect 12253 12665 12265 12668
rect 12299 12665 12311 12699
rect 12253 12659 12311 12665
rect 11882 12628 11888 12640
rect 11532 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12406 12628 12434 12736
rect 14182 12628 14188 12640
rect 12406 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3234 12424 3240 12436
rect 2915 12396 3240 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4706 12424 4712 12436
rect 4479 12396 4712 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 4798 12384 4804 12436
rect 4856 12384 4862 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 6972 12396 7113 12424
rect 6972 12384 6978 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7101 12387 7159 12393
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3326 12288 3332 12300
rect 3007 12260 3332 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3476 12260 3985 12288
rect 3476 12248 3482 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 5350 12288 5356 12300
rect 3973 12251 4031 12257
rect 5000 12260 5356 12288
rect 5000 12232 5028 12260
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 7116 12288 7144 12387
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 11425 12427 11483 12433
rect 9456 12396 9720 12424
rect 9456 12384 9462 12396
rect 7377 12291 7435 12297
rect 5684 12260 5856 12288
rect 7116 12260 7328 12288
rect 5684 12248 5690 12260
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 992 12192 1409 12220
rect 992 12180 998 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2409 12223 2467 12229
rect 2409 12220 2421 12223
rect 2096 12192 2421 12220
rect 2096 12180 2102 12192
rect 2409 12189 2421 12192
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2677 12223 2735 12229
rect 2677 12189 2689 12223
rect 2723 12216 2735 12223
rect 3050 12220 3056 12232
rect 2792 12216 3056 12220
rect 2723 12192 3056 12216
rect 2723 12189 2820 12192
rect 2677 12188 2820 12189
rect 2677 12183 2735 12188
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 2501 12155 2559 12161
rect 2501 12121 2513 12155
rect 2547 12152 2559 12155
rect 3234 12152 3240 12164
rect 2547 12124 3240 12152
rect 2547 12121 2559 12124
rect 2501 12115 2559 12121
rect 3234 12112 3240 12124
rect 3292 12152 3298 12164
rect 3804 12152 3832 12183
rect 3292 12124 3832 12152
rect 4908 12152 4936 12183
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 5718 12180 5724 12232
rect 5776 12180 5782 12232
rect 5828 12220 5856 12260
rect 7300 12232 7328 12260
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 7423 12260 8033 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 8021 12257 8033 12260
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 5828 12192 7205 12220
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7340 12192 7941 12220
rect 7340 12180 7346 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 8573 12223 8631 12229
rect 8573 12220 8585 12223
rect 8352 12192 8585 12220
rect 8352 12180 8358 12192
rect 8573 12189 8585 12192
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 5988 12155 6046 12161
rect 4908 12124 5120 12152
rect 3292 12112 3298 12124
rect 5092 12096 5120 12124
rect 5988 12121 6000 12155
rect 6034 12152 6046 12155
rect 6730 12152 6736 12164
rect 6034 12124 6736 12152
rect 6034 12121 6046 12124
rect 5988 12115 6046 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 9692 12161 9720 12396
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 11606 12424 11612 12436
rect 11471 12396 11612 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 14415 12396 14872 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 14844 12368 14872 12396
rect 11882 12316 11888 12368
rect 11940 12316 11946 12368
rect 14826 12316 14832 12368
rect 14884 12316 14890 12368
rect 9950 12288 9956 12300
rect 9784 12260 9956 12288
rect 9784 12229 9812 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11296 12260 11713 12288
rect 11296 12248 11302 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9916 12192 10057 12220
rect 9916 12180 9922 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10301 12223 10359 12229
rect 10301 12220 10313 12223
rect 10192 12192 10313 12220
rect 10192 12180 10198 12192
rect 10301 12189 10313 12192
rect 10347 12189 10359 12223
rect 10301 12183 10359 12189
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11790 12220 11796 12232
rect 11563 12192 11796 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 7708 12124 7849 12152
rect 7708 12112 7714 12124
rect 7837 12121 7849 12124
rect 7883 12152 7895 12155
rect 9033 12155 9091 12161
rect 9033 12152 9045 12155
rect 7883 12124 9045 12152
rect 7883 12121 7895 12124
rect 7837 12115 7895 12121
rect 9033 12121 9045 12124
rect 9079 12121 9091 12155
rect 9033 12115 9091 12121
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12121 9183 12155
rect 9125 12115 9183 12121
rect 9677 12155 9735 12161
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 9723 12124 12434 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 1578 12044 1584 12096
rect 1636 12044 1642 12096
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 3878 12084 3884 12096
rect 3651 12056 3884 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 5074 12044 5080 12096
rect 5132 12044 5138 12096
rect 8665 12087 8723 12093
rect 8665 12053 8677 12087
rect 8711 12084 8723 12087
rect 9140 12084 9168 12115
rect 8711 12056 9168 12084
rect 8711 12053 8723 12056
rect 8665 12047 8723 12053
rect 9950 12044 9956 12096
rect 10008 12044 10014 12096
rect 12406 12084 12434 12124
rect 13906 12084 13912 12096
rect 12406 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 1578 11840 1584 11892
rect 1636 11840 1642 11892
rect 2409 11883 2467 11889
rect 2409 11849 2421 11883
rect 2455 11880 2467 11883
rect 3142 11880 3148 11892
rect 2455 11852 3148 11880
rect 2455 11849 2467 11852
rect 2409 11843 2467 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4706 11880 4712 11892
rect 4663 11852 4712 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 4893 11883 4951 11889
rect 4893 11849 4905 11883
rect 4939 11880 4951 11883
rect 5166 11880 5172 11892
rect 4939 11852 5172 11880
rect 4939 11849 4951 11852
rect 4893 11843 4951 11849
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7190 11840 7196 11892
rect 7248 11840 7254 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7650 11880 7656 11892
rect 7515 11852 7656 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 9950 11840 9956 11892
rect 10008 11840 10014 11892
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11882 11880 11888 11892
rect 11011 11852 11888 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11744 1455 11747
rect 1596 11744 1624 11840
rect 1964 11784 2452 11812
rect 1964 11753 1992 11784
rect 1443 11716 1624 11744
rect 1857 11747 1915 11753
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1857 11713 1869 11747
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 1949 11707 2007 11713
rect 2148 11716 2237 11744
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1872 11676 1900 11707
rect 992 11648 1900 11676
rect 992 11636 998 11648
rect 2148 11617 2176 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2424 11676 2452 11784
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 3252 11753 3280 11840
rect 4632 11784 8248 11812
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 3326 11676 3332 11688
rect 2424 11648 3332 11676
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 3510 11636 3516 11688
rect 3568 11676 3574 11688
rect 3973 11679 4031 11685
rect 3973 11676 3985 11679
rect 3568 11648 3985 11676
rect 3568 11636 3574 11648
rect 3973 11645 3985 11648
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 4154 11636 4160 11688
rect 4212 11636 4218 11688
rect 2133 11611 2191 11617
rect 1504 11580 2084 11608
rect 1504 11549 1532 11580
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11509 1547 11543
rect 1489 11503 1547 11509
rect 1670 11500 1676 11552
rect 1728 11500 1734 11552
rect 2056 11540 2084 11580
rect 2133 11577 2145 11611
rect 2179 11577 2191 11611
rect 4632 11608 4660 11784
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4755 11716 5028 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5000 11617 5028 11716
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 5132 11716 5181 11744
rect 5132 11704 5138 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 5169 11707 5227 11713
rect 6656 11716 8125 11744
rect 5184 11676 5212 11707
rect 6549 11679 6607 11685
rect 5184 11648 6040 11676
rect 6012 11620 6040 11648
rect 6549 11645 6561 11679
rect 6595 11645 6607 11679
rect 6549 11639 6607 11645
rect 2133 11571 2191 11577
rect 2746 11580 4660 11608
rect 4985 11611 5043 11617
rect 2746 11540 2774 11580
rect 4985 11577 4997 11611
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 5994 11568 6000 11620
rect 6052 11568 6058 11620
rect 2056 11512 2774 11540
rect 3142 11500 3148 11552
rect 3200 11500 3206 11552
rect 3878 11500 3884 11552
rect 3936 11500 3942 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 6564 11540 6592 11639
rect 6656 11552 6684 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 8220 11676 8248 11784
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 9968 11753 9996 11840
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 10778 11744 10784 11756
rect 9953 11707 10011 11713
rect 10428 11716 10784 11744
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 8220 11648 10333 11676
rect 7929 11639 7987 11645
rect 10321 11645 10333 11648
rect 10367 11676 10379 11679
rect 10428 11676 10456 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 13906 11704 13912 11756
rect 13964 11704 13970 11756
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 14047 11716 14197 11744
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 10367 11648 10456 11676
rect 10505 11679 10563 11685
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10505 11645 10517 11679
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11676 11575 11679
rect 11606 11676 11612 11688
rect 11563 11648 11612 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 7944 11608 7972 11639
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 7944 11580 8217 11608
rect 8205 11577 8217 11580
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 10137 11611 10195 11617
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 10520 11608 10548 11639
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 10183 11580 10548 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 4120 11512 6592 11540
rect 4120 11500 4126 11512
rect 6638 11500 6644 11552
rect 6696 11500 6702 11552
rect 14366 11500 14372 11552
rect 14424 11500 14430 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4154 11296 4160 11348
rect 4212 11296 4218 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 6273 11339 6331 11345
rect 5307 11308 5856 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 1688 11132 1716 11296
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11268 3111 11271
rect 4172 11268 4200 11296
rect 3099 11240 4200 11268
rect 5353 11271 5411 11277
rect 3099 11237 3111 11240
rect 3053 11231 3111 11237
rect 5353 11237 5365 11271
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 1627 11104 1716 11132
rect 2961 11135 3019 11141
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3050 11132 3056 11144
rect 3007 11104 3056 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3384 11104 3525 11132
rect 3384 11092 3390 11104
rect 3513 11101 3525 11104
rect 3559 11132 3571 11135
rect 3970 11132 3976 11144
rect 3559 11104 3976 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5368 11132 5396 11231
rect 5828 11209 5856 11308
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6638 11336 6644 11348
rect 6319 11308 6644 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 8386 11336 8392 11348
rect 7423 11308 8392 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 5813 11203 5871 11209
rect 5123 11104 5396 11132
rect 5460 11172 5764 11200
rect 5460 11132 5488 11172
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5460 11104 5549 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5537 11101 5549 11104
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5736 11132 5764 11172
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 6656 11200 6684 11296
rect 6748 11268 6776 11296
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 6748 11240 7573 11268
rect 7561 11237 7573 11240
rect 7607 11237 7619 11271
rect 7561 11231 7619 11237
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 6656 11172 9321 11200
rect 5813 11163 5871 11169
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9309 11163 9367 11169
rect 9876 11172 10057 11200
rect 9876 11144 9904 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11112 11172 11529 11200
rect 11112 11160 11118 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 6825 11135 6883 11141
rect 5736 11104 6040 11132
rect 5629 11095 5687 11101
rect 1673 11067 1731 11073
rect 1673 11033 1685 11067
rect 1719 11064 1731 11067
rect 5644 11064 5672 11095
rect 6012 11076 6040 11104
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 6914 11132 6920 11144
rect 6871 11104 6920 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7282 11132 7288 11144
rect 7239 11104 7288 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8251 11104 8423 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 1719 11036 5672 11064
rect 1719 11033 1731 11036
rect 1673 11027 1731 11033
rect 5552 11008 5580 11036
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 8395 11064 8423 11104
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8680 11104 9045 11132
rect 6052 11036 8423 11064
rect 6052 11024 6058 11036
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 6730 10956 6736 11008
rect 6788 10956 6794 11008
rect 7098 10956 7104 11008
rect 7156 10956 7162 11008
rect 8294 10956 8300 11008
rect 8352 10956 8358 11008
rect 8395 10996 8423 11036
rect 8680 11008 8708 11104
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9171 11104 9781 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10134 11132 10140 11144
rect 9999 11104 10140 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10312 11135 10370 11141
rect 10312 11101 10324 11135
rect 10358 11132 10370 11135
rect 10594 11132 10600 11144
rect 10358 11104 10600 11132
rect 10358 11101 10370 11104
rect 10312 11095 10370 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11132 11759 11135
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11747 11104 12357 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12452 11064 12480 11095
rect 11440 11036 12480 11064
rect 8662 10996 8668 11008
rect 8395 10968 8668 10996
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11440 11005 11468 11036
rect 11425 10999 11483 11005
rect 11425 10996 11437 10999
rect 11112 10968 11437 10996
rect 11112 10956 11118 10968
rect 11425 10965 11437 10968
rect 11471 10965 11483 10999
rect 11425 10959 11483 10965
rect 12158 10956 12164 11008
rect 12216 10956 12222 11008
rect 12406 10996 12434 11036
rect 13906 10996 13912 11008
rect 12406 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 1026 10684 1032 10736
rect 1084 10724 1090 10736
rect 5902 10724 5908 10736
rect 1084 10696 2084 10724
rect 1084 10684 1090 10696
rect 2056 10665 2084 10696
rect 5552 10696 5908 10724
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 2041 10659 2099 10665
rect 1811 10628 1900 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1872 10529 1900 10628
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 4798 10656 4804 10668
rect 4755 10628 4804 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 5552 10665 5580 10696
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 7558 10684 7564 10736
rect 7616 10724 7622 10736
rect 8478 10724 8484 10736
rect 7616 10696 8484 10724
rect 7616 10684 7622 10696
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 10594 10724 10600 10736
rect 9968 10696 10600 10724
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4856 10628 4997 10656
rect 4856 10616 4862 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5276 10588 5304 10619
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5868 10628 6377 10656
rect 5868 10616 5874 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6730 10656 6736 10668
rect 6595 10628 6736 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7064 10628 7849 10656
rect 7064 10616 7070 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 9968 10665 9996 10696
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 11348 10724 11376 10755
rect 12158 10752 12164 10804
rect 12216 10752 12222 10804
rect 11348 10696 12480 10724
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 4908 10560 5304 10588
rect 5721 10591 5779 10597
rect 4908 10529 4936 10560
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10489 1915 10523
rect 1857 10483 1915 10489
rect 4893 10523 4951 10529
rect 4893 10489 4905 10523
rect 4939 10489 4951 10523
rect 4893 10483 4951 10489
rect 5445 10523 5503 10529
rect 5445 10489 5457 10523
rect 5491 10520 5503 10523
rect 5736 10520 5764 10551
rect 7098 10548 7104 10600
rect 7156 10548 7162 10600
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 8312 10588 8340 10616
rect 7331 10560 8340 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 5491 10492 5764 10520
rect 9692 10520 9720 10619
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 11112 10628 11161 10656
rect 11112 10616 11118 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11606 10656 11612 10668
rect 11563 10628 11612 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12452 10665 12480 10696
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 11701 10591 11759 10597
rect 9815 10560 11468 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 9950 10520 9956 10532
rect 9692 10492 9956 10520
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 9950 10480 9956 10492
rect 10008 10480 10014 10532
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 11330 10520 11336 10532
rect 10091 10492 11336 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 3418 10452 3424 10464
rect 1719 10424 3424 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5626 10452 5632 10464
rect 5123 10424 5632 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5994 10412 6000 10464
rect 6052 10412 6058 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7055 10424 7757 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7745 10421 7757 10424
rect 7791 10452 7803 10455
rect 8294 10452 8300 10464
rect 7791 10424 8300 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 8536 10424 9137 10452
rect 8536 10412 8542 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 11440 10452 11468 10560
rect 11701 10557 11713 10591
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 11716 10520 11744 10551
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11716 10492 12265 10520
rect 12253 10489 12265 10492
rect 12299 10489 12311 10523
rect 12253 10483 12311 10489
rect 14200 10452 14228 10619
rect 11440 10424 14228 10452
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 3436 10220 12081 10248
rect 3436 10112 3464 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 3789 10183 3847 10189
rect 3789 10149 3801 10183
rect 3835 10180 3847 10183
rect 4062 10180 4068 10192
rect 3835 10152 4068 10180
rect 3835 10149 3847 10152
rect 3789 10143 3847 10149
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 8662 10140 8668 10192
rect 8720 10180 8726 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8720 10152 9045 10180
rect 8720 10140 8726 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9033 10143 9091 10149
rect 11149 10183 11207 10189
rect 11149 10149 11161 10183
rect 11195 10180 11207 10183
rect 11606 10180 11612 10192
rect 11195 10152 11612 10180
rect 11195 10149 11207 10152
rect 11149 10143 11207 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 3344 10084 3464 10112
rect 8496 10084 9352 10112
rect 3142 10004 3148 10056
rect 3200 10053 3206 10056
rect 3200 10044 3212 10053
rect 3200 10016 3245 10044
rect 3200 10007 3212 10016
rect 3200 10004 3206 10007
rect 1765 9979 1823 9985
rect 1765 9945 1777 9979
rect 1811 9976 1823 9979
rect 3344 9976 3372 10084
rect 8496 10056 8524 10084
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 3467 10016 5181 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 5169 10013 5181 10016
rect 5215 10044 5227 10047
rect 5718 10044 5724 10056
rect 5215 10016 5724 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5718 10004 5724 10016
rect 5776 10044 5782 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 5776 10016 6837 10044
rect 5776 10004 5782 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 8478 10044 8484 10056
rect 7147 10016 8484 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 9324 10044 9352 10084
rect 10502 10072 10508 10124
rect 10560 10072 10566 10124
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11388 10084 11437 10112
rect 11388 10072 11394 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 9858 10044 9864 10056
rect 9324 10016 9864 10044
rect 8573 10007 8631 10013
rect 1811 9948 3372 9976
rect 1811 9945 1823 9948
rect 1765 9939 1823 9945
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 4902 9979 4960 9985
rect 4902 9976 4914 9979
rect 4764 9948 4914 9976
rect 4764 9936 4770 9948
rect 4902 9945 4914 9948
rect 4948 9945 4960 9979
rect 4902 9939 4960 9945
rect 5261 9979 5319 9985
rect 5261 9945 5273 9979
rect 5307 9976 5319 9979
rect 7006 9976 7012 9988
rect 5307 9948 7012 9976
rect 5307 9945 5319 9948
rect 5261 9939 5319 9945
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7346 9979 7404 9985
rect 7346 9976 7358 9979
rect 7248 9948 7358 9976
rect 7248 9936 7254 9948
rect 7346 9945 7358 9948
rect 7392 9945 7404 9979
rect 8588 9976 8616 10007
rect 9858 10004 9864 10016
rect 9916 10044 9922 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9916 10016 10425 10044
rect 9916 10004 9922 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 12158 10004 12164 10056
rect 12216 10004 12222 10056
rect 8588 9948 9904 9976
rect 7346 9939 7404 9945
rect 9876 9920 9904 9948
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10146 9979 10204 9985
rect 10146 9976 10158 9979
rect 10100 9948 10158 9976
rect 10100 9936 10106 9948
rect 10146 9945 10158 9948
rect 10192 9945 10204 9979
rect 10146 9939 10204 9945
rect 13538 9936 13544 9988
rect 13596 9936 13602 9988
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 3142 9908 3148 9920
rect 2087 9880 3148 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 8478 9868 8484 9920
rect 8536 9868 8542 9920
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9306 9908 9312 9920
rect 8803 9880 9312 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13780 9880 13829 9908
rect 13780 9868 13786 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 13817 9871 13875 9877
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 4525 9707 4583 9713
rect 3068 9676 4384 9704
rect 3068 9636 3096 9676
rect 1780 9608 3096 9636
rect 4356 9636 4384 9676
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 4706 9704 4712 9716
rect 4571 9676 4712 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 6052 9676 6193 9704
rect 6052 9664 6058 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 4356 9608 5396 9636
rect 1780 9577 1808 9608
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 1912 9540 2881 9568
rect 1912 9528 1918 9540
rect 2869 9537 2881 9540
rect 2915 9568 2927 9571
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2915 9540 3065 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3528 9500 3556 9531
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 4062 9568 4068 9580
rect 3660 9540 4068 9568
rect 3660 9528 3666 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5040 9540 5273 9568
rect 5040 9528 5046 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 3694 9500 3700 9512
rect 3528 9472 3700 9500
rect 3694 9460 3700 9472
rect 3752 9500 3758 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3752 9472 3893 9500
rect 3752 9460 3758 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4798 9500 4804 9512
rect 4212 9472 4804 9500
rect 4212 9460 4218 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 5092 9432 5120 9463
rect 3467 9404 5120 9432
rect 5368 9432 5396 9608
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5684 9540 5733 9568
rect 5684 9528 5690 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 6196 9568 6224 9667
rect 10042 9664 10048 9716
rect 10100 9664 10106 9716
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 8536 9608 9536 9636
rect 8536 9596 8542 9608
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 6196 9540 6377 9568
rect 5721 9531 5779 9537
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 7282 9528 7288 9580
rect 7340 9528 7346 9580
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 9508 9577 9536 9608
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10962 9636 10968 9648
rect 10652 9608 10968 9636
rect 10652 9596 10658 9608
rect 10962 9596 10968 9608
rect 11020 9636 11026 9648
rect 11020 9608 11284 9636
rect 11020 9596 11026 9608
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 7892 9540 9137 9568
rect 7892 9528 7898 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 10226 9568 10232 9580
rect 9539 9540 10232 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 11256 9577 11284 9608
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10827 9540 11161 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11606 9568 11612 9580
rect 11563 9540 11612 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6052 9472 6561 9500
rect 6052 9460 6058 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 10965 9503 11023 9509
rect 7064 9472 8616 9500
rect 7064 9460 7070 9472
rect 7466 9432 7472 9444
rect 5368 9404 7472 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 8588 9441 8616 9472
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9401 8631 9435
rect 10980 9432 11008 9463
rect 11698 9460 11704 9512
rect 11756 9460 11762 9512
rect 12250 9460 12256 9512
rect 12308 9460 12314 9512
rect 13814 9432 13820 9444
rect 10980 9404 13820 9432
rect 8573 9395 8631 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 1670 9324 1676 9376
rect 1728 9324 1734 9376
rect 2222 9324 2228 9376
rect 2280 9324 2286 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3510 9364 3516 9376
rect 3191 9336 3516 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4338 9364 4344 9376
rect 3743 9336 4344 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7650 9364 7656 9376
rect 7055 9336 7656 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 9217 9367 9275 9373
rect 9217 9364 9229 9367
rect 8444 9336 9229 9364
rect 8444 9324 8450 9336
rect 9217 9333 9229 9336
rect 9263 9333 9275 9367
rect 9217 9327 9275 9333
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 1670 9120 1676 9172
rect 1728 9120 1734 9172
rect 2222 9120 2228 9172
rect 2280 9120 2286 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 3694 9160 3700 9172
rect 3651 9132 3700 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 4338 9120 4344 9172
rect 4396 9120 4402 9172
rect 4706 9120 4712 9172
rect 4764 9120 4770 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 7291 9132 10333 9160
rect 1688 8956 1716 9120
rect 2240 9024 2268 9120
rect 2240 8996 2360 9024
rect 1765 8959 1823 8965
rect 1765 8956 1777 8959
rect 1688 8928 1777 8956
rect 1765 8925 1777 8928
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2332 8956 2360 8996
rect 2481 8959 2539 8965
rect 2481 8956 2493 8959
rect 2332 8928 2493 8956
rect 2225 8919 2283 8925
rect 2481 8925 2493 8928
rect 2527 8925 2539 8959
rect 2481 8919 2539 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 2240 8888 2268 8919
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3712 8956 3740 9120
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3712 8928 3801 8956
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 3252 8888 3280 8916
rect 2240 8860 3280 8888
rect 4080 8888 4108 8919
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4356 8888 4384 9120
rect 4724 9024 4752 9120
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7291 9092 7319 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10686 9160 10692 9172
rect 10551 9132 10692 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11793 9163 11851 9169
rect 10980 9132 11192 9160
rect 6788 9064 7319 9092
rect 9769 9095 9827 9101
rect 6788 9052 6794 9064
rect 9769 9061 9781 9095
rect 9815 9092 9827 9095
rect 9950 9092 9956 9104
rect 9815 9064 9956 9092
rect 9815 9061 9827 9064
rect 9769 9055 9827 9061
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 10980 9092 11008 9132
rect 10428 9064 11008 9092
rect 11057 9095 11115 9101
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 4724 8996 4905 9024
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 5040 8996 5181 9024
rect 5040 8984 5046 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8352 8996 9229 9024
rect 8352 8984 8358 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 7156 8928 8677 8956
rect 7156 8916 7162 8928
rect 8665 8925 8677 8928
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10226 8956 10232 8968
rect 10183 8928 10232 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 4080 8860 4292 8888
rect 4356 8860 4997 8888
rect 1397 8851 1455 8857
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4154 8820 4160 8832
rect 4019 8792 4160 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4264 8820 4292 8860
rect 4985 8857 4997 8860
rect 5031 8857 5043 8891
rect 4985 8851 5043 8857
rect 5896 8891 5954 8897
rect 5896 8857 5908 8891
rect 5942 8888 5954 8891
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 5942 8860 8125 8888
rect 5942 8857 5954 8860
rect 5896 8851 5954 8857
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 6730 8820 6736 8832
rect 4264 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6972 8792 7021 8820
rect 6972 8780 6978 8792
rect 7009 8789 7021 8792
rect 7055 8820 7067 8823
rect 7834 8820 7840 8832
rect 7055 8792 7840 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8680 8820 8708 8919
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10428 8965 10456 9064
rect 11057 9061 11069 9095
rect 11103 9061 11115 9095
rect 11164 9092 11192 9132
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 11882 9160 11888 9172
rect 11839 9132 11888 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12176 9132 12388 9160
rect 12176 9092 12204 9132
rect 11164 9064 12204 9092
rect 12253 9095 12311 9101
rect 11057 9055 11115 9061
rect 12253 9061 12265 9095
rect 12299 9061 12311 9095
rect 12360 9092 12388 9132
rect 12452 9132 13492 9160
rect 12452 9092 12480 9132
rect 12360 9064 12480 9092
rect 12529 9095 12587 9101
rect 12253 9055 12311 9061
rect 12529 9061 12541 9095
rect 12575 9092 12587 9095
rect 12575 9064 12664 9092
rect 12575 9061 12587 9064
rect 12529 9055 12587 9061
rect 11072 9024 11100 9055
rect 10704 8996 11100 9024
rect 11977 9027 12035 9033
rect 10704 8965 10732 8996
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 12268 9024 12296 9055
rect 12023 8996 12296 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 9306 8848 9312 8900
rect 9364 8848 9370 8900
rect 10428 8888 10456 8919
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11020 8928 11253 8956
rect 11020 8916 11026 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12250 8956 12256 8968
rect 12207 8928 12256 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 12636 8956 12664 9064
rect 12483 8928 12664 8956
rect 12713 8959 12771 8965
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 13464 8956 13492 9132
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13596 9132 13737 9160
rect 13596 9120 13602 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 14369 9163 14427 9169
rect 14369 9129 14381 9163
rect 14415 9160 14427 9163
rect 14415 9132 14872 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 14844 9104 14872 9132
rect 14826 9052 14832 9104
rect 14884 9052 14890 9104
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 12759 8928 12848 8956
rect 13464 8928 13921 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 9646 8860 10088 8888
rect 9646 8820 9674 8860
rect 10060 8832 10088 8860
rect 10244 8860 10456 8888
rect 10244 8832 10272 8860
rect 8680 8792 9674 8820
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 9916 8792 9965 8820
rect 9916 8780 9922 8792
rect 9953 8789 9965 8792
rect 9999 8789 10011 8823
rect 9953 8783 10011 8789
rect 10042 8780 10048 8832
rect 10100 8780 10106 8832
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 10560 8792 10793 8820
rect 10560 8780 10566 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 10781 8783 10839 8789
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 12820 8820 12848 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 13909 8919 13967 8925
rect 14182 8916 14188 8968
rect 14240 8916 14246 8968
rect 11664 8792 12848 8820
rect 11664 8780 11670 8792
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1854 8576 1860 8628
rect 1912 8576 1918 8628
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8585 3755 8619
rect 3697 8579 3755 8585
rect 2958 8440 2964 8492
rect 3016 8489 3022 8492
rect 3016 8480 3028 8489
rect 3513 8483 3571 8489
rect 3016 8452 3061 8480
rect 3016 8443 3028 8452
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 3620 8480 3648 8576
rect 3559 8452 3648 8480
rect 3712 8480 3740 8579
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 5902 8616 5908 8628
rect 4571 8588 5908 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4080 8489 4108 8576
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3712 8452 3801 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4264 8480 4292 8579
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7708 8588 7941 8616
rect 7708 8576 7714 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 9600 8588 10364 8616
rect 4801 8551 4859 8557
rect 4801 8548 4813 8551
rect 4448 8520 4813 8548
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4264 8452 4353 8480
rect 4065 8443 4123 8449
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 3016 8440 3022 8443
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 3694 8412 3700 8424
rect 3292 8384 3700 8412
rect 3292 8372 3298 8384
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4448 8412 4476 8520
rect 4801 8517 4813 8520
rect 4847 8517 4859 8551
rect 4801 8511 4859 8517
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 7098 8548 7104 8560
rect 4948 8520 7104 8548
rect 4948 8508 4954 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 7944 8548 7972 8579
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 7944 8520 9045 8548
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 9033 8511 9091 8517
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 9600 8548 9628 8588
rect 10336 8560 10364 8588
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11698 8616 11704 8628
rect 11195 8588 11704 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 11940 8588 13124 8616
rect 11940 8576 11946 8588
rect 9171 8520 9628 8548
rect 9677 8551 9735 8557
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 9677 8517 9689 8551
rect 9723 8548 9735 8551
rect 9950 8548 9956 8560
rect 9723 8520 9956 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10318 8508 10324 8560
rect 10376 8508 10382 8560
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 13096 8557 13124 8588
rect 13081 8551 13139 8557
rect 10652 8520 12940 8548
rect 10652 8508 10658 8520
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7650 8480 7656 8492
rect 6779 8452 7656 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 9692 8452 10517 8480
rect 4356 8400 4476 8412
rect 4172 8384 4476 8400
rect 4172 8372 4384 8384
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8412 6607 8415
rect 6822 8412 6828 8424
rect 6595 8384 6828 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4172 8344 4200 8372
rect 4019 8316 4200 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 5000 8344 5028 8372
rect 4488 8316 5028 8344
rect 6104 8344 6132 8375
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7248 8384 7297 8412
rect 7248 8372 7254 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 8404 8412 8432 8440
rect 7515 8384 8432 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 8662 8372 8668 8424
rect 8720 8372 8726 8424
rect 6104 8316 6592 8344
rect 4488 8304 4494 8316
rect 6564 8288 6592 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 3016 8248 5457 8276
rect 3016 8236 3022 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5445 8239 5503 8245
rect 6546 8236 6552 8288
rect 6604 8236 6610 8288
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 8168 8248 8217 8276
rect 8168 8236 8174 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9692 8276 9720 8452
rect 10505 8449 10517 8452
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10744 8452 10793 8480
rect 10744 8440 10750 8452
rect 10781 8449 10793 8452
rect 10827 8480 10839 8483
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10827 8452 11069 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11057 8449 11069 8452
rect 11103 8480 11115 8483
rect 11606 8480 11612 8492
rect 11103 8452 11612 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 12641 8483 12699 8489
rect 12641 8449 12653 8483
rect 12687 8480 12699 8483
rect 12802 8480 12808 8492
rect 12687 8452 12808 8480
rect 12687 8449 12699 8452
rect 12641 8443 12699 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 12912 8489 12940 8520
rect 13081 8517 13093 8551
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 13173 8551 13231 8557
rect 13173 8517 13185 8551
rect 13219 8548 13231 8551
rect 13814 8548 13820 8560
rect 13219 8520 13820 8548
rect 13219 8517 13231 8520
rect 13173 8511 13231 8517
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 9784 8344 9812 8375
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 10100 8384 11560 8412
rect 10100 8372 10106 8384
rect 10778 8344 10784 8356
rect 9784 8316 10784 8344
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11238 8344 11244 8356
rect 11011 8316 11244 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 11532 8353 11560 8384
rect 13280 8384 13369 8412
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 13280 8288 13308 8384
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14458 8344 14464 8356
rect 14415 8316 14464 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 9180 8248 9720 8276
rect 9180 8236 9186 8248
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 10100 8248 10149 8276
rect 10100 8236 10106 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 10137 8239 10195 8245
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 13262 8276 13268 8288
rect 12676 8248 13268 8276
rect 12676 8236 12682 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1854 8032 1860 8084
rect 1912 8032 1918 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6914 8072 6920 8084
rect 6696 8044 6920 8072
rect 6696 8032 6702 8044
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8720 8044 9045 8072
rect 8720 8032 8726 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 12802 8032 12808 8084
rect 12860 8032 12866 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 1872 7936 1900 8032
rect 3694 7964 3700 8016
rect 3752 8004 3758 8016
rect 6273 8007 6331 8013
rect 3752 7976 4936 8004
rect 3752 7964 3758 7976
rect 1872 7908 2360 7936
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 2332 7877 2360 7908
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 3568 7908 4261 7936
rect 3568 7896 3574 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 4706 7936 4712 7948
rect 4663 7908 4712 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 992 7840 1409 7868
rect 992 7828 998 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2823 7840 2881 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 1765 7803 1823 7809
rect 1765 7769 1777 7803
rect 1811 7800 1823 7803
rect 2041 7803 2099 7809
rect 2041 7800 2053 7803
rect 1811 7772 2053 7800
rect 1811 7769 1823 7772
rect 1765 7763 1823 7769
rect 2041 7769 2053 7772
rect 2087 7769 2099 7803
rect 2148 7800 2176 7831
rect 3050 7828 3056 7880
rect 3108 7828 3114 7880
rect 4908 7877 4936 7976
rect 6273 7973 6285 8007
rect 6319 8004 6331 8007
rect 6546 8004 6552 8016
rect 6319 7976 6552 8004
rect 6319 7973 6331 7976
rect 6273 7967 6331 7973
rect 6546 7964 6552 7976
rect 6604 8004 6610 8016
rect 6604 7976 7880 8004
rect 6604 7964 6610 7976
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 5960 7908 6929 7936
rect 5960 7896 5966 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7156 7908 7788 7936
rect 7156 7896 7162 7908
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 5626 7868 5632 7880
rect 4939 7840 5632 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 4338 7800 4344 7812
rect 2148 7772 4344 7800
rect 2041 7763 2099 7769
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 2498 7692 2504 7744
rect 2556 7692 2562 7744
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3568 7704 3801 7732
rect 3568 7692 3574 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 4448 7732 4476 7831
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 6638 7828 6644 7880
rect 6696 7828 6702 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7760 7877 7788 7908
rect 7852 7877 7880 7976
rect 10042 7964 10048 8016
rect 10100 7964 10106 8016
rect 11333 8007 11391 8013
rect 11333 8004 11345 8007
rect 10796 7976 11345 8004
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9030 7936 9036 7948
rect 8803 7908 9036 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9030 7896 9036 7908
rect 9088 7936 9094 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9088 7908 9413 7936
rect 9088 7896 9094 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 10060 7936 10088 7964
rect 10796 7945 10824 7976
rect 11333 7973 11345 7976
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 12618 7964 12624 8016
rect 12676 7964 12682 8016
rect 13725 8007 13783 8013
rect 13725 7973 13737 8007
rect 13771 7973 13783 8007
rect 13725 7967 13783 7973
rect 10597 7939 10655 7945
rect 10597 7936 10609 7939
rect 10060 7908 10609 7936
rect 9401 7899 9459 7905
rect 10597 7905 10609 7908
rect 10643 7905 10655 7939
rect 10597 7899 10655 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 11900 7908 13369 7936
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7883 7840 8248 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 5160 7803 5218 7809
rect 5160 7769 5172 7803
rect 5206 7800 5218 7803
rect 5258 7800 5264 7812
rect 5206 7772 5264 7800
rect 5206 7769 5218 7772
rect 5160 7763 5218 7769
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 8110 7800 8116 7812
rect 6380 7772 6592 7800
rect 6380 7732 6408 7772
rect 4448 7704 6408 7732
rect 3789 7695 3847 7701
rect 6454 7692 6460 7744
rect 6512 7692 6518 7744
rect 6564 7732 6592 7772
rect 6932 7772 8116 7800
rect 6932 7732 6960 7772
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8220 7800 8248 7840
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 8956 7800 8984 7831
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10502 7868 10508 7880
rect 10367 7840 10508 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11256 7868 11284 7896
rect 11900 7880 11928 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11256 7840 11529 7868
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 13372 7868 13400 7899
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13372 7840 13553 7868
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13740 7868 13768 7967
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13740 7840 14289 7868
rect 13541 7831 13599 7837
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 8220 7772 8984 7800
rect 11241 7803 11299 7809
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 12066 7800 12072 7812
rect 11287 7772 12072 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7769 12219 7803
rect 12161 7763 12219 7769
rect 6564 7704 6960 7732
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8202 7732 8208 7744
rect 8067 7704 8208 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 11793 7735 11851 7741
rect 11793 7701 11805 7735
rect 11839 7732 11851 7735
rect 12176 7732 12204 7763
rect 11839 7704 12204 7732
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 3050 7528 3056 7540
rect 2746 7500 3056 7528
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2516 7392 2544 7488
rect 2363 7364 2544 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2222 7284 2228 7336
rect 2280 7284 2286 7336
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2464 7296 2605 7324
rect 2464 7284 2470 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 2746 7256 2774 7500
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 5258 7488 5264 7540
rect 5316 7488 5322 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6052 7500 6193 7528
rect 6052 7488 6058 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6181 7491 6239 7497
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7558 7528 7564 7540
rect 7331 7500 7564 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 8570 7488 8576 7540
rect 8628 7488 8634 7540
rect 9030 7488 9036 7540
rect 9088 7488 9094 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 9640 7500 10885 7528
rect 9640 7488 9646 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 12124 7500 12434 7528
rect 12124 7488 12130 7500
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 3936 7432 6684 7460
rect 3936 7420 3942 7432
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3476 7364 3525 7392
rect 3476 7352 3482 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4304 7364 4445 7392
rect 4304 7352 4310 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4939 7364 4997 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5350 7392 5356 7404
rect 5031 7364 5356 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5350 7352 5356 7364
rect 5408 7392 5414 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5408 7364 5825 7392
rect 5408 7352 5414 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6454 7392 6460 7404
rect 6043 7364 6460 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 3694 7284 3700 7336
rect 3752 7284 3758 7336
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 6546 7284 6552 7336
rect 6604 7284 6610 7336
rect 6656 7324 6684 7432
rect 6932 7392 6960 7488
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 6932 7364 7113 7392
rect 7101 7361 7113 7364
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8220 7392 8248 7488
rect 12406 7460 12434 7500
rect 13262 7488 13268 7540
rect 13320 7488 13326 7540
rect 12897 7463 12955 7469
rect 12897 7460 12909 7463
rect 12406 7432 12909 7460
rect 12897 7429 12909 7432
rect 12943 7429 12955 7463
rect 12897 7423 12955 7429
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8220 7364 8401 7392
rect 8113 7355 8171 7361
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 8895 7364 8984 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6656 7296 7389 7324
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 2547 7228 2774 7256
rect 4801 7259 4859 7265
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 4801 7225 4813 7259
rect 4847 7256 4859 7259
rect 5626 7256 5632 7268
rect 4847 7228 5632 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 8128 7256 8156 7355
rect 8956 7336 8984 7364
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9576 7395 9634 7401
rect 9576 7361 9588 7395
rect 9622 7392 9634 7395
rect 9858 7392 9864 7404
rect 9622 7364 9864 7392
rect 9622 7361 9634 7364
rect 9576 7355 9634 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 10928 7364 10977 7392
rect 10928 7352 10934 7364
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 11195 7364 12449 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 12437 7361 12449 7364
rect 12483 7361 12495 7395
rect 13280 7392 13308 7488
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13280 7364 13921 7392
rect 12437 7355 12495 7361
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 14047 7364 14197 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 11072 7324 11100 7355
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 10704 7296 12081 7324
rect 10704 7268 10732 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 7392 7228 8156 7256
rect 8220 7228 8769 7256
rect 7392 7200 7420 7228
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 992 7160 1501 7188
rect 992 7148 998 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 4154 7148 4160 7200
rect 4212 7148 4218 7200
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 6454 7188 6460 7200
rect 5215 7160 6460 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6914 7148 6920 7200
rect 6972 7148 6978 7200
rect 7374 7148 7380 7200
rect 7432 7148 7438 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7524 7160 7757 7188
rect 7524 7148 7530 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8220 7188 8248 7228
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 10410 7216 10416 7268
rect 10468 7216 10474 7268
rect 10686 7216 10692 7268
rect 10744 7216 10750 7268
rect 12268 7256 12296 7287
rect 11164 7228 12296 7256
rect 7892 7160 8248 7188
rect 7892 7148 7898 7160
rect 8294 7148 8300 7200
rect 8352 7148 8358 7200
rect 10428 7188 10456 7216
rect 11164 7188 11192 7228
rect 10428 7160 11192 7188
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11296 7160 11529 7188
rect 11296 7148 11302 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 14366 7148 14372 7200
rect 14424 7148 14430 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 1762 6984 1768 6996
rect 1719 6956 1768 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3694 6984 3700 6996
rect 3559 6956 3700 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 4212 6956 5304 6984
rect 4212 6944 4218 6956
rect 5276 6916 5304 6956
rect 5350 6944 5356 6996
rect 5408 6944 5414 6996
rect 8294 6944 8300 6996
rect 8352 6944 8358 6996
rect 9858 6944 9864 6996
rect 9916 6944 9922 6996
rect 10612 6956 12434 6984
rect 7285 6919 7343 6925
rect 7285 6916 7297 6919
rect 5276 6888 7297 6916
rect 7285 6885 7297 6888
rect 7331 6916 7343 6919
rect 8312 6916 8340 6944
rect 10612 6916 10640 6956
rect 7331 6888 8064 6916
rect 8312 6888 10640 6916
rect 7331 6885 7343 6888
rect 7285 6879 7343 6885
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2280 6820 2605 6848
rect 2280 6808 2286 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3844 6820 3985 6848
rect 3844 6808 3850 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 8036 6857 8064 6888
rect 11882 6876 11888 6928
rect 11940 6916 11946 6928
rect 11977 6919 12035 6925
rect 11977 6916 11989 6919
rect 11940 6888 11989 6916
rect 11940 6876 11946 6888
rect 11977 6885 11989 6888
rect 12023 6885 12035 6919
rect 12406 6916 12434 6956
rect 14090 6916 14096 6928
rect 12406 6888 14096 6916
rect 11977 6879 12035 6885
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6788 6820 6929 6848
rect 6788 6808 6794 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6848 7159 6851
rect 8021 6851 8079 6857
rect 7147 6820 7604 6848
rect 7147 6817 7159 6820
rect 7101 6811 7159 6817
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 1780 6712 1808 6743
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2406 6740 2412 6792
rect 2464 6780 2470 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2464 6752 2789 6780
rect 2464 6740 2470 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7024 6780 7144 6782
rect 6871 6754 7420 6780
rect 6871 6752 7052 6754
rect 7116 6752 7420 6754
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 3510 6712 3516 6724
rect 1780 6684 3516 6712
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 4246 6721 4252 6724
rect 4240 6675 4252 6721
rect 4246 6672 4252 6675
rect 4304 6672 4310 6724
rect 5445 6715 5503 6721
rect 5445 6712 5457 6715
rect 4908 6684 5457 6712
rect 4908 6656 4936 6684
rect 5445 6681 5457 6684
rect 5491 6681 5503 6715
rect 5445 6675 5503 6681
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5684 6684 6009 6712
rect 5684 6672 5690 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 6089 6715 6147 6721
rect 6089 6681 6101 6715
rect 6135 6712 6147 6715
rect 6914 6712 6920 6724
rect 6135 6684 6920 6712
rect 6135 6681 6147 6684
rect 6089 6675 6147 6681
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 7392 6656 7420 6752
rect 7576 6712 7604 6820
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 10594 6848 10600 6860
rect 9364 6820 10600 6848
rect 9364 6808 9370 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 12805 6851 12863 6857
rect 12805 6817 12817 6851
rect 12851 6848 12863 6851
rect 13173 6851 13231 6857
rect 13173 6848 13185 6851
rect 12851 6820 13185 6848
rect 12851 6817 12863 6820
rect 12805 6811 12863 6817
rect 13173 6817 13185 6820
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7708 6752 7757 6780
rect 7708 6740 7714 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10864 6783 10922 6789
rect 10551 6752 10824 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 7834 6712 7840 6724
rect 7576 6684 7840 6712
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8220 6712 8248 6743
rect 10796 6724 10824 6752
rect 10864 6749 10876 6783
rect 10910 6780 10922 6783
rect 11238 6780 11244 6792
rect 10910 6752 11244 6780
rect 10910 6749 10922 6752
rect 10864 6743 10922 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12989 6783 13047 6789
rect 12989 6780 13001 6783
rect 12584 6752 13001 6780
rect 12584 6740 12590 6752
rect 12989 6749 13001 6752
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 7944 6684 8248 6712
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 2556 6616 3249 6644
rect 2556 6604 2562 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 4890 6604 4896 6656
rect 4948 6604 4954 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6638 6644 6644 6656
rect 6595 6616 6644 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 7944 6653 7972 6684
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 13096 6712 13124 6743
rect 14182 6740 14188 6792
rect 14240 6740 14246 6792
rect 12820 6684 13124 6712
rect 12820 6656 12848 6684
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 9272 6616 12357 6644
rect 9272 6604 9278 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 14366 6604 14372 6656
rect 14424 6604 14430 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 3326 6400 3332 6452
rect 3384 6400 3390 6452
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 3620 6412 3893 6440
rect 2148 6344 2728 6372
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 2148 6313 2176 6344
rect 2700 6313 2728 6344
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3142 6304 3148 6316
rect 2731 6276 3148 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2240 6168 2268 6267
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3620 6313 3648 6412
rect 3881 6409 3893 6412
rect 3927 6409 3939 6443
rect 3881 6403 3939 6409
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4246 6440 4252 6452
rect 4203 6412 4252 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6362 6440 6368 6452
rect 6227 6412 6368 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6457 6443 6515 6449
rect 6457 6409 6469 6443
rect 6503 6440 6515 6443
rect 6546 6440 6552 6452
rect 6503 6412 6552 6440
rect 6503 6409 6515 6412
rect 6457 6403 6515 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7285 6443 7343 6449
rect 7285 6440 7297 6443
rect 6972 6412 7297 6440
rect 6972 6400 6978 6412
rect 7285 6409 7297 6412
rect 7331 6409 7343 6443
rect 7285 6403 7343 6409
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7708 6412 7941 6440
rect 7708 6400 7714 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8720 6412 8861 6440
rect 8720 6400 8726 6412
rect 8849 6409 8861 6412
rect 8895 6440 8907 6443
rect 9858 6440 9864 6452
rect 8895 6412 9864 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10468 6412 10701 6440
rect 10468 6400 10474 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 10689 6403 10747 6409
rect 4890 6372 4896 6384
rect 4448 6344 4896 6372
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3605 6267 3663 6273
rect 3988 6276 4077 6304
rect 3528 6236 3556 6267
rect 3988 6248 4016 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 3970 6236 3976 6248
rect 3528 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 2501 6171 2559 6177
rect 2501 6168 2513 6171
rect 2240 6140 2513 6168
rect 2501 6137 2513 6140
rect 2547 6137 2559 6171
rect 4448 6168 4476 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 5445 6375 5503 6381
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 5491 6344 6500 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6043 6276 6377 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5583 6208 5733 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 2501 6131 2559 6137
rect 2746 6140 4476 6168
rect 4816 6168 4844 6199
rect 6012 6180 6040 6267
rect 5994 6168 6000 6180
rect 4816 6140 6000 6168
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 2746 6100 2774 6140
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 6472 6168 6500 6344
rect 6656 6304 6684 6400
rect 7576 6372 7604 6400
rect 7745 6375 7803 6381
rect 7745 6372 7757 6375
rect 7576 6344 7757 6372
rect 7745 6341 7757 6344
rect 7791 6341 7803 6375
rect 7745 6335 7803 6341
rect 8938 6332 8944 6384
rect 8996 6372 9002 6384
rect 12802 6372 12808 6384
rect 8996 6344 12808 6372
rect 8996 6332 9002 6344
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6656 6276 6837 6304
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 7883 6276 8125 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8113 6273 8125 6276
rect 8159 6304 8171 6307
rect 8754 6304 8760 6316
rect 8159 6276 8760 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6730 6236 6736 6248
rect 6687 6208 6736 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7377 6171 7435 6177
rect 7377 6168 7389 6171
rect 6472 6140 7389 6168
rect 7377 6137 7389 6140
rect 7423 6137 7435 6171
rect 7377 6131 7435 6137
rect 2188 6072 2774 6100
rect 3789 6103 3847 6109
rect 2188 6060 2194 6072
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4062 6100 4068 6112
rect 3835 6072 4068 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 7576 6100 7604 6267
rect 8754 6264 8760 6276
rect 8812 6304 8818 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8812 6276 9137 6304
rect 8812 6264 8818 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9953 6307 10011 6313
rect 9539 6276 9812 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8389 6239 8447 6245
rect 8251 6208 8340 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8312 6180 8340 6208
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8435 6208 9045 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 9232 6168 9260 6264
rect 9784 6177 9812 6276
rect 9953 6273 9965 6307
rect 9999 6304 10011 6307
rect 10318 6304 10324 6316
rect 9999 6276 10324 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 10318 6264 10324 6276
rect 10376 6304 10382 6316
rect 10778 6304 10784 6316
rect 10376 6276 10784 6304
rect 10376 6264 10382 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 8352 6140 9260 6168
rect 9769 6171 9827 6177
rect 8352 6128 8358 6140
rect 9769 6137 9781 6171
rect 9815 6137 9827 6171
rect 9769 6131 9827 6137
rect 6512 6072 7604 6100
rect 9677 6103 9735 6109
rect 6512 6060 6518 6072
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 10244 6100 10272 6199
rect 9723 6072 10272 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2041 5899 2099 5905
rect 2041 5896 2053 5899
rect 1820 5868 2053 5896
rect 1820 5856 1826 5868
rect 2041 5865 2053 5868
rect 2087 5865 2099 5899
rect 2041 5859 2099 5865
rect 2498 5856 2504 5908
rect 2556 5856 2562 5908
rect 3786 5856 3792 5908
rect 3844 5856 3850 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4028 5868 6040 5896
rect 4028 5856 4034 5868
rect 2516 5769 2544 5856
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 3329 5831 3387 5837
rect 3329 5828 3341 5831
rect 2648 5800 3341 5828
rect 2648 5788 2654 5800
rect 3329 5797 3341 5800
rect 3375 5797 3387 5831
rect 3329 5791 3387 5797
rect 2501 5763 2559 5769
rect 2501 5729 2513 5763
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 3142 5720 3148 5772
rect 3200 5720 3206 5772
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 3804 5760 3832 5856
rect 6012 5828 6040 5868
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 6144 5868 6469 5896
rect 6144 5856 6150 5868
rect 6457 5865 6469 5868
rect 6503 5865 6515 5899
rect 6457 5859 6515 5865
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 6822 5896 6828 5908
rect 6779 5868 6828 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8846 5856 8852 5908
rect 8904 5856 8910 5908
rect 9306 5896 9312 5908
rect 8956 5868 9312 5896
rect 8864 5828 8892 5856
rect 6012 5800 8892 5828
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 3660 5732 5089 5760
rect 3660 5720 3666 5732
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 8294 5760 8300 5772
rect 5077 5723 5135 5729
rect 6748 5732 8300 5760
rect 2130 5652 2136 5704
rect 2188 5652 2194 5704
rect 3160 5692 3188 5720
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 3160 5664 3525 5692
rect 3513 5661 3525 5664
rect 3559 5692 3571 5695
rect 3694 5692 3700 5704
rect 3559 5664 3700 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 4120 5664 4169 5692
rect 4120 5652 4126 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 6748 5692 6776 5732
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8956 5769 8984 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14240 5868 14289 5896
rect 14240 5856 14246 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 4663 5664 6776 5692
rect 6825 5695 6883 5701
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 6871 5664 8340 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5593 1823 5627
rect 1765 5587 1823 5593
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 1780 5556 1808 5587
rect 2590 5584 2596 5636
rect 2648 5584 2654 5636
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 3326 5624 3332 5636
rect 3191 5596 3332 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 5350 5633 5356 5636
rect 5344 5587 5356 5633
rect 5350 5584 5356 5587
rect 5408 5584 5414 5636
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 6840 5624 6868 5655
rect 6052 5596 6868 5624
rect 6052 5584 6058 5596
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 7524 5596 7941 5624
rect 7524 5584 7530 5596
rect 7668 5568 7696 5596
rect 7929 5593 7941 5596
rect 7975 5593 7987 5627
rect 7929 5587 7987 5593
rect 3234 5556 3240 5568
rect 1780 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5534 5556 5540 5568
rect 5031 5528 5540 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 8312 5556 8340 5664
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 10594 5692 10600 5704
rect 8619 5664 10600 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 12406 5664 14105 5692
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9186 5627 9244 5633
rect 9186 5624 9198 5627
rect 9088 5596 9198 5624
rect 9088 5584 9094 5596
rect 9186 5593 9198 5596
rect 9232 5593 9244 5627
rect 9186 5587 9244 5593
rect 12406 5556 12434 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 13538 5584 13544 5636
rect 13596 5584 13602 5636
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 15010 5624 15016 5636
rect 13955 5596 15016 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 8312 5528 12434 5556
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2590 5352 2596 5364
rect 2271 5324 2596 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3602 5352 3608 5364
rect 3108 5324 3608 5352
rect 3108 5312 3114 5324
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 7006 5352 7012 5364
rect 4356 5324 7012 5352
rect 2409 5287 2467 5293
rect 2409 5253 2421 5287
rect 2455 5284 2467 5287
rect 3786 5284 3792 5296
rect 2455 5256 3792 5284
rect 2455 5253 2467 5256
rect 2409 5247 2467 5253
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 4356 5293 4384 5324
rect 7006 5312 7012 5324
rect 7064 5352 7070 5364
rect 7064 5324 7880 5352
rect 7064 5312 7070 5324
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5253 4399 5287
rect 4341 5247 4399 5253
rect 5350 5244 5356 5296
rect 5408 5244 5414 5296
rect 5534 5244 5540 5296
rect 5592 5244 5598 5296
rect 5626 5244 5632 5296
rect 5684 5244 5690 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 7852 5293 7880 5324
rect 9306 5312 9312 5364
rect 9364 5312 9370 5364
rect 9416 5324 12434 5352
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5253 7895 5287
rect 7837 5247 7895 5253
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 9416 5284 9444 5324
rect 8076 5256 9444 5284
rect 8076 5244 8082 5256
rect 9766 5244 9772 5296
rect 9824 5244 9830 5296
rect 9858 5244 9864 5296
rect 9916 5244 9922 5296
rect 10686 5244 10692 5296
rect 10744 5244 10750 5296
rect 1762 5176 1768 5228
rect 1820 5176 1826 5228
rect 2038 5176 2044 5228
rect 2096 5176 2102 5228
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 2501 5219 2559 5225
rect 2501 5216 2513 5219
rect 2280 5188 2513 5216
rect 2280 5176 2286 5188
rect 2501 5185 2513 5188
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 8478 5216 8484 5228
rect 7331 5188 8484 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 4448 5148 4476 5179
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 12406 5216 12434 5324
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 12406 5188 14197 5216
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 4706 5148 4712 5160
rect 4448 5120 4712 5148
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5859 5120 6377 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5148 7067 5151
rect 7190 5148 7196 5160
rect 7055 5120 7196 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 5828 5080 5856 5111
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 8386 5108 8392 5160
rect 8444 5108 8450 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 8496 5120 10609 5148
rect 3160 5052 5856 5080
rect 7469 5083 7527 5089
rect 3160 5024 3188 5052
rect 7469 5049 7481 5083
rect 7515 5080 7527 5083
rect 8404 5080 8432 5108
rect 7515 5052 8432 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 3142 4972 3148 5024
rect 3200 4972 3206 5024
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 4798 5012 4804 5024
rect 4663 4984 4804 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 8496 5012 8524 5120
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10888 5080 10916 5111
rect 10367 5052 11008 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 7708 4984 8524 5012
rect 10980 5012 11008 5052
rect 14090 5012 14096 5024
rect 10980 4984 14096 5012
rect 7708 4972 7714 4984
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3234 4808 3240 4820
rect 3099 4780 3240 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 8018 4808 8024 4820
rect 3651 4780 8024 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9030 4768 9036 4820
rect 9088 4768 9094 4820
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10686 4808 10692 4820
rect 10551 4780 10692 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 13538 4808 13544 4820
rect 11103 4780 13544 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 4154 4700 4160 4752
rect 4212 4700 4218 4752
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 8803 4712 9628 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3050 4672 3056 4684
rect 2915 4644 3056 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 9600 4681 9628 4712
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 2222 4564 2228 4616
rect 2280 4564 2286 4616
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2602 4607 2660 4613
rect 2602 4604 2614 4607
rect 2372 4576 2614 4604
rect 2372 4564 2378 4576
rect 2602 4573 2614 4576
rect 2648 4573 2660 4607
rect 2602 4567 2660 4573
rect 3142 4564 3148 4616
rect 3200 4564 3206 4616
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 2240 4536 2268 4564
rect 3436 4536 3464 4567
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4246 4604 4252 4616
rect 4019 4576 4252 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 2240 4508 3464 4536
rect 5752 4539 5810 4545
rect 5752 4505 5764 4539
rect 5798 4536 5810 4539
rect 6012 4536 6040 4567
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6696 4576 6837 4604
rect 6696 4564 6702 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 9324 4604 9352 4632
rect 7423 4576 9352 4604
rect 9600 4604 9628 4635
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9600 4576 9965 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 9953 4573 9965 4576
rect 9999 4604 10011 4607
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9999 4576 10057 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10045 4567 10103 4573
rect 10244 4576 10333 4604
rect 6730 4536 6736 4548
rect 5798 4508 5948 4536
rect 6012 4508 6736 4536
rect 5798 4505 5810 4508
rect 5752 4499 5810 4505
rect 1489 4471 1547 4477
rect 1489 4437 1501 4471
rect 1535 4468 1547 4471
rect 2130 4468 2136 4480
rect 1535 4440 2136 4468
rect 1535 4437 1547 4440
rect 1489 4431 1547 4437
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 4706 4468 4712 4480
rect 4663 4440 4712 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 4706 4428 4712 4440
rect 4764 4468 4770 4480
rect 5534 4468 5540 4480
rect 4764 4440 5540 4468
rect 4764 4428 4770 4440
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5920 4468 5948 4508
rect 6730 4496 6736 4508
rect 6788 4536 6794 4548
rect 7392 4536 7420 4567
rect 7650 4545 7656 4548
rect 6788 4508 7420 4536
rect 6788 4496 6794 4508
rect 7644 4499 7656 4545
rect 7650 4496 7656 4499
rect 7708 4496 7714 4548
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5920 4440 6101 4468
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 6914 4428 6920 4480
rect 6972 4428 6978 4480
rect 10244 4477 10272 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 10870 4564 10876 4616
rect 10928 4564 10934 4616
rect 14090 4564 14096 4616
rect 14148 4564 14154 4616
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4437 10287 4471
rect 10229 4431 10287 4437
rect 14182 4428 14188 4480
rect 14240 4428 14246 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 4304 4236 4629 4264
rect 4304 4224 4310 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 4617 4227 4675 4233
rect 4798 4224 4804 4276
rect 4856 4224 4862 4276
rect 5077 4267 5135 4273
rect 5077 4233 5089 4267
rect 5123 4264 5135 4267
rect 5442 4264 5448 4276
rect 5123 4236 5448 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5592 4236 6408 4264
rect 5592 4224 5598 4236
rect 2406 4156 2412 4208
rect 2464 4196 2470 4208
rect 3421 4199 3479 4205
rect 3421 4196 3433 4199
rect 2464 4168 3433 4196
rect 2464 4156 2470 4168
rect 3421 4165 3433 4168
rect 3467 4165 3479 4199
rect 3421 4159 3479 4165
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 1946 4128 1952 4140
rect 1811 4100 1952 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2130 4088 2136 4140
rect 2188 4088 2194 4140
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 3752 4100 4537 4128
rect 3752 4088 3758 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4816 4128 4844 4224
rect 5810 4156 5816 4208
rect 5868 4156 5874 4208
rect 6380 4137 6408 4236
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 8113 4267 8171 4273
rect 8113 4264 8125 4267
rect 7708 4236 8125 4264
rect 7708 4224 7714 4236
rect 8113 4233 8125 4236
rect 8159 4233 8171 4267
rect 8113 4227 8171 4233
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 8536 4236 9597 4264
rect 8536 4224 8542 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 8772 4168 9674 4196
rect 8772 4140 8800 4168
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4816 4100 4905 4128
rect 4525 4091 4583 4097
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6730 4128 6736 4140
rect 6687 4100 6736 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6908 4131 6966 4137
rect 6908 4097 6920 4131
rect 6954 4128 6966 4131
rect 6954 4112 8616 4128
rect 6954 4100 8708 4112
rect 6954 4097 6966 4100
rect 6908 4091 6966 4097
rect 8588 4084 8708 4100
rect 8754 4088 8760 4140
rect 8812 4088 8818 4140
rect 9646 4128 9674 4168
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9646 4100 9781 4128
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3326 4060 3332 4072
rect 3283 4032 3332 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 4154 4060 4160 4072
rect 3559 4032 4160 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4246 4020 4252 4072
rect 4304 4020 4310 4072
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4706 4060 4712 4072
rect 4479 4032 4712 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5307 4032 5396 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4172 3992 4200 4020
rect 4111 3964 4200 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 5368 3936 5396 4032
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5592 4032 5917 4060
rect 5592 4020 5598 4032
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 8680 3992 8708 4084
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 8996 4032 9321 4060
rect 8996 4020 9002 4032
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 10502 4060 10508 4072
rect 9539 4032 10508 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 12802 4060 12808 4072
rect 10643 4032 12808 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 8680 3964 9965 3992
rect 9953 3961 9965 3964
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 992 3896 1501 3924
rect 992 3884 998 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 2556 3896 2789 3924
rect 2556 3884 2562 3896
rect 2777 3893 2789 3896
rect 2823 3893 2835 3927
rect 2777 3887 2835 3893
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 7006 3924 7012 3936
rect 6503 3896 7012 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8754 3924 8760 3936
rect 8067 3896 8760 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8846 3884 8852 3936
rect 8904 3884 8910 3936
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 4246 3720 4252 3732
rect 2179 3692 4252 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6638 3720 6644 3732
rect 6319 3692 6644 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7745 3723 7803 3729
rect 7248 3692 7696 3720
rect 7248 3680 7254 3692
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 7668 3652 7696 3692
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8938 3720 8944 3732
rect 7791 3692 8944 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 10042 3720 10048 3732
rect 9815 3692 10048 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 8846 3652 8852 3664
rect 5960 3624 7328 3652
rect 7668 3624 8852 3652
rect 5960 3612 5966 3624
rect 3970 3584 3976 3596
rect 3804 3556 3976 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1728 3488 1777 3516
rect 1728 3476 1734 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 3050 3516 3056 3528
rect 2271 3488 3056 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 992 3420 1409 3448
rect 992 3408 998 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 1964 3448 1992 3479
rect 3050 3476 3056 3488
rect 3108 3516 3114 3528
rect 3804 3516 3832 3556
rect 3970 3544 3976 3556
rect 4028 3584 4034 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4028 3556 4905 3584
rect 4028 3544 4034 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 6914 3584 6920 3596
rect 6779 3556 6920 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 3108 3488 3832 3516
rect 4525 3519 4583 3525
rect 3108 3476 3114 3488
rect 4525 3485 4537 3519
rect 4571 3516 4583 3519
rect 6549 3519 6607 3525
rect 4571 3488 6500 3516
rect 4571 3485 4583 3488
rect 4525 3479 4583 3485
rect 2314 3448 2320 3460
rect 1964 3420 2320 3448
rect 1397 3411 1455 3417
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 2498 3457 2504 3460
rect 2492 3448 2504 3457
rect 2459 3420 2504 3448
rect 2492 3411 2504 3420
rect 2498 3408 2504 3411
rect 2556 3408 2562 3460
rect 4540 3448 4568 3479
rect 3620 3420 4568 3448
rect 5160 3451 5218 3457
rect 3620 3389 3648 3420
rect 5160 3417 5172 3451
rect 5206 3448 5218 3451
rect 5258 3448 5264 3460
rect 5206 3420 5264 3448
rect 5206 3417 5218 3420
rect 5160 3411 5218 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 6472 3448 6500 3488
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6822 3516 6828 3528
rect 6595 3488 6828 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7300 3525 7328 3624
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 9784 3584 9812 3683
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 10560 3692 12081 3720
rect 10560 3680 10566 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 10870 3612 10876 3664
rect 10928 3612 10934 3664
rect 9631 3556 9812 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8159 3488 8401 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 8527 3488 9413 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 8128 3448 8156 3479
rect 9858 3476 9864 3528
rect 9916 3516 9922 3528
rect 10888 3516 10916 3612
rect 9916 3488 10916 3516
rect 12161 3519 12219 3525
rect 9916 3476 9922 3488
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12526 3516 12532 3528
rect 12207 3488 12532 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 14185 3519 14243 3525
rect 14185 3516 14197 3519
rect 13964 3488 14197 3516
rect 13964 3476 13970 3488
rect 14185 3485 14197 3488
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 6472 3420 8156 3448
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11790 3448 11796 3460
rect 11204 3420 11796 3448
rect 11204 3408 11210 3420
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3349 3663 3383
rect 3605 3343 3663 3349
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4062 3380 4068 3392
rect 4019 3352 4068 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 8294 3340 8300 3392
rect 8352 3340 8358 3392
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 14366 3340 14372 3392
rect 14424 3340 14430 3392
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 1762 3176 1768 3188
rect 1719 3148 1768 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 1946 3136 1952 3188
rect 2004 3136 2010 3188
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 2096 3148 2145 3176
rect 2096 3136 2102 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 2133 3139 2191 3145
rect 3712 3148 5365 3176
rect 1964 3108 1992 3136
rect 2501 3111 2559 3117
rect 2501 3108 2513 3111
rect 1964 3080 2513 3108
rect 2501 3077 2513 3080
rect 2547 3077 2559 3111
rect 2501 3071 2559 3077
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2130 3040 2136 3052
rect 1903 3012 2136 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 1780 2904 1808 3003
rect 2130 3000 2136 3012
rect 2188 3040 2194 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2188 3012 2329 3040
rect 2188 3000 2194 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 3326 3040 3332 3052
rect 2639 3012 3332 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3712 3049 3740 3148
rect 5353 3145 5365 3148
rect 5399 3176 5411 3179
rect 5718 3176 5724 3188
rect 5399 3148 5724 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5718 3136 5724 3148
rect 5776 3176 5782 3188
rect 5902 3176 5908 3188
rect 5776 3148 5908 3176
rect 5776 3136 5782 3148
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 7374 3176 7380 3188
rect 6012 3148 7380 3176
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 6012 3117 6040 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 8938 3176 8944 3188
rect 8711 3148 8944 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 4218 3111 4276 3117
rect 4218 3108 4230 3111
rect 4120 3080 4230 3108
rect 4120 3068 4126 3080
rect 4218 3077 4230 3080
rect 4264 3077 4276 3111
rect 4218 3071 4276 3077
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3077 6055 3111
rect 5997 3071 6055 3077
rect 6638 3068 6644 3120
rect 6696 3068 6702 3120
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 3970 3000 3976 3052
rect 4028 3000 4034 3052
rect 5350 3040 5356 3052
rect 4080 3012 5356 3040
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2424 2972 2452 3000
rect 4080 2972 4108 3012
rect 5350 3000 5356 3012
rect 5408 3040 5414 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5408 3012 5457 3040
rect 5408 3000 5414 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6656 3040 6684 3068
rect 6595 3012 6684 3040
rect 8312 3040 8340 3136
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8312 3012 8401 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 1995 2944 2452 2972
rect 2746 2944 4108 2972
rect 6089 2975 6147 2981
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2746 2904 2774 2944
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 8680 2972 8708 3139
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9364 3148 10916 3176
rect 9364 3136 9370 3148
rect 10888 3108 10916 3148
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 11020 3148 14289 3176
rect 11020 3136 11026 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14277 3139 14335 3145
rect 10888 3080 11560 3108
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10686 3040 10692 3052
rect 9999 3012 10692 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 11238 3040 11244 3052
rect 10919 3012 11244 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11532 3049 11560 3080
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11784 3043 11842 3049
rect 11784 3009 11796 3043
rect 11830 3040 11842 3043
rect 13722 3040 13728 3052
rect 11830 3012 13728 3040
rect 11830 3009 11842 3012
rect 11784 3003 11842 3009
rect 6135 2944 8708 2972
rect 9125 2975 9183 2981
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 9355 2944 10793 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 6733 2907 6791 2913
rect 1780 2876 2774 2904
rect 5276 2876 5488 2904
rect 3881 2839 3939 2845
rect 3881 2805 3893 2839
rect 3927 2836 3939 2839
rect 5276 2836 5304 2876
rect 3927 2808 5304 2836
rect 5460 2836 5488 2876
rect 6733 2873 6745 2907
rect 6779 2904 6791 2907
rect 7558 2904 7564 2916
rect 6779 2876 7564 2904
rect 6779 2873 6791 2876
rect 6733 2867 6791 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2904 8631 2907
rect 9140 2904 9168 2935
rect 11146 2932 11152 2984
rect 11204 2932 11210 2984
rect 8619 2876 9168 2904
rect 9861 2907 9919 2913
rect 8619 2873 8631 2876
rect 8573 2867 8631 2873
rect 9861 2873 9873 2907
rect 9907 2904 9919 2907
rect 10134 2904 10140 2916
rect 9907 2876 10140 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 10134 2864 10140 2876
rect 10192 2864 10198 2916
rect 11164 2904 11192 2932
rect 11241 2907 11299 2913
rect 11241 2904 11253 2907
rect 11164 2876 11253 2904
rect 11241 2873 11253 2876
rect 11287 2873 11299 2907
rect 11241 2867 11299 2873
rect 5626 2836 5632 2848
rect 5460 2808 5632 2836
rect 3927 2805 3939 2808
rect 3881 2799 3939 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 11348 2836 11376 3003
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 15010 3040 15016 3052
rect 14507 3012 15016 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 12820 2876 14136 2904
rect 12820 2836 12848 2876
rect 14108 2848 14136 2876
rect 11348 2808 12848 2836
rect 12894 2796 12900 2848
rect 12952 2796 12958 2848
rect 14090 2796 14096 2848
rect 14148 2796 14154 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2280 2604 2421 2632
rect 2280 2592 2286 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4706 2632 4712 2644
rect 4663 2604 4712 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5258 2592 5264 2644
rect 5316 2592 5322 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5868 2604 6009 2632
rect 5868 2592 5874 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 7558 2592 7564 2644
rect 7616 2592 7622 2644
rect 9122 2592 9128 2644
rect 9180 2592 9186 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10226 2632 10232 2644
rect 10183 2604 10232 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11296 2604 11529 2632
rect 11296 2592 11302 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 12526 2592 12532 2644
rect 12584 2592 12590 2644
rect 13722 2592 13728 2644
rect 13780 2592 13786 2644
rect 14090 2592 14096 2644
rect 14148 2592 14154 2644
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2564 4491 2567
rect 5902 2564 5908 2576
rect 4479 2536 5908 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 7282 2496 7288 2508
rect 4120 2468 7288 2496
rect 4120 2456 4126 2468
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 13924 2468 14688 2496
rect 2222 2388 2228 2440
rect 2280 2388 2286 2440
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3476 2400 3801 2428
rect 3476 2388 3482 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4522 2428 4528 2440
rect 4295 2400 4528 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5534 2428 5540 2440
rect 5031 2400 5540 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 3970 2252 3976 2304
rect 4028 2252 4034 2304
rect 4724 2292 4752 2391
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5920 2400 6193 2428
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 5920 2360 5948 2400
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 5684 2332 5948 2360
rect 5684 2320 5690 2332
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 6564 2360 6592 2391
rect 7374 2388 7380 2440
rect 7432 2388 7438 2440
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8628 2400 8953 2428
rect 8628 2388 8634 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11204 2400 11713 2428
rect 11204 2388 11210 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13924 2437 13952 2468
rect 14660 2440 14688 2468
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12492 2400 12725 2428
rect 12492 2388 12498 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 6052 2332 6592 2360
rect 6052 2320 6058 2332
rect 6365 2295 6423 2301
rect 6365 2292 6377 2295
rect 4724 2264 6377 2292
rect 6365 2261 6377 2264
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 9766 2088 9772 2100
rect 4028 2060 9772 2088
rect 4028 2048 4034 2060
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
<< via1 >>
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 1032 17280 1084 17332
rect 1124 17280 1176 17332
rect 940 17144 992 17196
rect 2412 17280 2464 17332
rect 3792 17280 3844 17332
rect 5172 17280 5224 17332
rect 6552 17280 6604 17332
rect 8208 17280 8260 17332
rect 9312 17280 9364 17332
rect 10692 17280 10744 17332
rect 12072 17280 12124 17332
rect 14464 17280 14516 17332
rect 14556 17280 14608 17332
rect 4160 17144 4212 17196
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 14004 17144 14056 17196
rect 14096 17144 14148 17196
rect 2780 17076 2832 17128
rect 3700 17008 3752 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2136 16940 2188 16992
rect 11152 17076 11204 17128
rect 4252 16940 4304 16992
rect 4896 16940 4948 16992
rect 5724 16940 5776 16992
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 7196 16940 7248 16992
rect 9036 16940 9088 16992
rect 9864 16940 9916 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 13268 16983 13320 16992
rect 13268 16949 13277 16983
rect 13277 16949 13311 16983
rect 13311 16949 13320 16983
rect 13268 16940 13320 16949
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 1584 16736 1636 16788
rect 5632 16779 5684 16788
rect 5632 16745 5641 16779
rect 5641 16745 5675 16779
rect 5675 16745 5684 16779
rect 5632 16736 5684 16745
rect 1952 16600 2004 16652
rect 5816 16600 5868 16652
rect 940 16464 992 16516
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 3516 16396 3568 16448
rect 3884 16396 3936 16448
rect 4712 16507 4764 16516
rect 4712 16473 4721 16507
rect 4721 16473 4755 16507
rect 4755 16473 4764 16507
rect 4712 16464 4764 16473
rect 4804 16507 4856 16516
rect 4804 16473 4813 16507
rect 4813 16473 4847 16507
rect 4847 16473 4856 16507
rect 4804 16464 4856 16473
rect 5356 16507 5408 16516
rect 5356 16473 5365 16507
rect 5365 16473 5399 16507
rect 5399 16473 5408 16507
rect 5356 16464 5408 16473
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7196 16532 7248 16541
rect 7472 16532 7524 16584
rect 12164 16736 12216 16788
rect 13268 16736 13320 16788
rect 13360 16711 13412 16720
rect 13360 16677 13369 16711
rect 13369 16677 13403 16711
rect 13403 16677 13412 16711
rect 13360 16668 13412 16677
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10600 16532 10652 16584
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 10784 16532 10836 16541
rect 13360 16532 13412 16584
rect 13452 16532 13504 16584
rect 13912 16532 13964 16584
rect 5264 16396 5316 16448
rect 5816 16396 5868 16448
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 6828 16396 6880 16448
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 14096 16464 14148 16516
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 12532 16396 12584 16448
rect 13820 16439 13872 16448
rect 13820 16405 13829 16439
rect 13829 16405 13863 16439
rect 13863 16405 13872 16439
rect 13820 16396 13872 16405
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 2780 16192 2832 16244
rect 3056 16192 3108 16244
rect 3516 16192 3568 16244
rect 5908 16192 5960 16244
rect 6920 16192 6972 16244
rect 7288 16192 7340 16244
rect 7472 16235 7524 16244
rect 7472 16201 7481 16235
rect 7481 16201 7515 16235
rect 7515 16201 7524 16235
rect 7472 16192 7524 16201
rect 13912 16192 13964 16244
rect 14004 16192 14056 16244
rect 1032 16124 1084 16176
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 4252 16124 4304 16176
rect 5356 16124 5408 16176
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2412 15852 2464 15904
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 4712 15988 4764 16040
rect 6000 16031 6052 16040
rect 6000 15997 6009 16031
rect 6009 15997 6043 16031
rect 6043 15997 6052 16031
rect 6000 15988 6052 15997
rect 3884 15920 3936 15972
rect 6736 16031 6788 16040
rect 6736 15997 6745 16031
rect 6745 15997 6779 16031
rect 6779 15997 6788 16031
rect 6736 15988 6788 15997
rect 8484 16124 8536 16176
rect 9036 16124 9088 16176
rect 10692 16124 10744 16176
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 4528 15852 4580 15904
rect 5540 15852 5592 15904
rect 6460 15852 6512 15904
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 7472 15920 7524 15972
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 1676 15648 1728 15700
rect 3148 15648 3200 15700
rect 4160 15648 4212 15700
rect 4712 15691 4764 15700
rect 4712 15657 4721 15691
rect 4721 15657 4755 15691
rect 4755 15657 4764 15691
rect 4712 15648 4764 15657
rect 4804 15648 4856 15700
rect 5908 15648 5960 15700
rect 6460 15648 6512 15700
rect 6736 15648 6788 15700
rect 10324 15648 10376 15700
rect 10784 15648 10836 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 3424 15444 3476 15496
rect 3608 15487 3660 15496
rect 3608 15453 3617 15487
rect 3617 15453 3651 15487
rect 3651 15453 3660 15487
rect 3608 15444 3660 15453
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 3056 15308 3108 15360
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 5724 15376 5776 15428
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 6644 15444 6696 15496
rect 6828 15444 6880 15496
rect 9036 15444 9088 15496
rect 9128 15444 9180 15496
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 7472 15376 7524 15428
rect 8300 15419 8352 15428
rect 8300 15385 8309 15419
rect 8309 15385 8343 15419
rect 8343 15385 8352 15419
rect 8300 15376 8352 15385
rect 3884 15308 3936 15360
rect 4160 15308 4212 15360
rect 5356 15351 5408 15360
rect 5356 15317 5365 15351
rect 5365 15317 5399 15351
rect 5399 15317 5408 15351
rect 5356 15308 5408 15317
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 10048 15351 10100 15360
rect 10048 15317 10057 15351
rect 10057 15317 10091 15351
rect 10091 15317 10100 15351
rect 10048 15308 10100 15317
rect 14832 15580 14884 15632
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 13728 15308 13780 15360
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 3608 15104 3660 15156
rect 6000 15104 6052 15156
rect 6368 15104 6420 15156
rect 8300 15104 8352 15156
rect 10140 15104 10192 15156
rect 11152 15104 11204 15156
rect 3056 15079 3108 15088
rect 3056 15045 3090 15079
rect 3090 15045 3108 15079
rect 3056 15036 3108 15045
rect 5356 15079 5408 15088
rect 5356 15045 5374 15079
rect 5374 15045 5408 15079
rect 6644 15079 6696 15088
rect 5356 15036 5408 15045
rect 2044 14968 2096 15020
rect 2504 14968 2556 15020
rect 6644 15045 6678 15079
rect 6678 15045 6696 15079
rect 6644 15036 6696 15045
rect 8944 15036 8996 15088
rect 2412 14943 2464 14952
rect 2412 14909 2421 14943
rect 2421 14909 2455 14943
rect 2455 14909 2464 14943
rect 2412 14900 2464 14909
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 8852 14968 8904 15020
rect 10048 15036 10100 15088
rect 9680 14968 9732 15020
rect 10416 14968 10468 15020
rect 13360 15036 13412 15088
rect 12072 14968 12124 15020
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 5632 14943 5684 14952
rect 5632 14909 5641 14943
rect 5641 14909 5675 14943
rect 5675 14909 5684 14943
rect 5632 14900 5684 14909
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 10508 14943 10560 14952
rect 10508 14909 10517 14943
rect 10517 14909 10551 14943
rect 10551 14909 10560 14943
rect 10508 14900 10560 14909
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 3056 14764 3108 14816
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5356 14764 5408 14816
rect 8300 14764 8352 14816
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 12440 14764 12492 14816
rect 12808 14764 12860 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 2044 14603 2096 14612
rect 2044 14569 2053 14603
rect 2053 14569 2087 14603
rect 2087 14569 2096 14603
rect 2044 14560 2096 14569
rect 2412 14560 2464 14612
rect 1584 14356 1636 14408
rect 5908 14560 5960 14612
rect 6828 14560 6880 14612
rect 7840 14560 7892 14612
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 9864 14560 9916 14612
rect 10508 14603 10560 14612
rect 10508 14569 10517 14603
rect 10517 14569 10551 14603
rect 10551 14569 10560 14603
rect 10508 14560 10560 14569
rect 10600 14560 10652 14612
rect 12808 14560 12860 14612
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 2688 14492 2740 14544
rect 5080 14492 5132 14544
rect 4160 14424 4212 14476
rect 4896 14424 4948 14476
rect 8116 14424 8168 14476
rect 8484 14424 8536 14476
rect 4988 14288 5040 14340
rect 5632 14288 5684 14340
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 9128 14356 9180 14408
rect 3240 14220 3292 14272
rect 4804 14220 4856 14272
rect 5172 14263 5224 14272
rect 5172 14229 5181 14263
rect 5181 14229 5215 14263
rect 5215 14229 5224 14263
rect 5172 14220 5224 14229
rect 6000 14220 6052 14272
rect 7196 14220 7248 14272
rect 10140 14356 10192 14408
rect 10232 14356 10284 14408
rect 12164 14356 12216 14408
rect 12624 14356 12676 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 11152 14288 11204 14340
rect 12440 14263 12492 14272
rect 12440 14229 12449 14263
rect 12449 14229 12483 14263
rect 12483 14229 12492 14263
rect 12440 14220 12492 14229
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 1676 14016 1728 14068
rect 2044 13744 2096 13796
rect 1768 13676 1820 13728
rect 2504 13676 2556 13728
rect 3240 13948 3292 14000
rect 4804 13948 4856 14000
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 5080 13880 5132 13932
rect 5632 13880 5684 13932
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 8300 13880 8352 13932
rect 3148 13676 3200 13728
rect 4528 13676 4580 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 7840 13676 7892 13728
rect 9956 13948 10008 14000
rect 10232 13948 10284 14000
rect 9864 13676 9916 13728
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 12624 14016 12676 14068
rect 12716 14016 12768 14068
rect 13452 14016 13504 14068
rect 13268 13948 13320 14000
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 14464 13812 14516 13864
rect 11244 13676 11296 13728
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 1768 13472 1820 13524
rect 4528 13515 4580 13524
rect 4528 13481 4537 13515
rect 4537 13481 4571 13515
rect 4571 13481 4580 13515
rect 4528 13472 4580 13481
rect 3056 13336 3108 13388
rect 5816 13472 5868 13524
rect 10140 13472 10192 13524
rect 11152 13472 11204 13524
rect 11704 13472 11756 13524
rect 12716 13472 12768 13524
rect 5540 13336 5592 13388
rect 8300 13336 8352 13388
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 2504 13311 2556 13320
rect 2504 13277 2522 13311
rect 2522 13277 2556 13311
rect 2504 13268 2556 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 3056 13200 3108 13252
rect 5080 13200 5132 13252
rect 1400 13175 1452 13184
rect 1400 13141 1409 13175
rect 1409 13141 1443 13175
rect 1443 13141 1452 13175
rect 1400 13132 1452 13141
rect 5172 13132 5224 13184
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 6184 13132 6236 13184
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 6920 13268 6972 13320
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 11612 13336 11664 13388
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 13360 13268 13412 13320
rect 7840 13200 7892 13252
rect 9128 13243 9180 13252
rect 9128 13209 9137 13243
rect 9137 13209 9171 13243
rect 9171 13209 9180 13243
rect 9128 13200 9180 13209
rect 7288 13132 7340 13184
rect 8760 13175 8812 13184
rect 8760 13141 8769 13175
rect 8769 13141 8803 13175
rect 8803 13141 8812 13175
rect 8760 13132 8812 13141
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 11888 13132 11940 13184
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 1400 12928 1452 12980
rect 940 12860 992 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 3332 12928 3384 12980
rect 3700 12928 3752 12980
rect 4896 12928 4948 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 6644 12928 6696 12980
rect 8300 12928 8352 12980
rect 9128 12928 9180 12980
rect 11888 12928 11940 12980
rect 2504 12792 2556 12844
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 5908 12792 5960 12844
rect 6000 12792 6052 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 9312 12860 9364 12912
rect 9864 12860 9916 12912
rect 12164 12903 12216 12912
rect 12164 12869 12173 12903
rect 12173 12869 12207 12903
rect 12207 12869 12216 12903
rect 12164 12860 12216 12869
rect 7288 12835 7340 12844
rect 7288 12801 7322 12835
rect 7322 12801 7340 12835
rect 7288 12792 7340 12801
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8760 12835 8812 12844
rect 8760 12801 8794 12835
rect 8794 12801 8812 12835
rect 8760 12792 8812 12801
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 9956 12724 10008 12776
rect 10876 12724 10928 12776
rect 3148 12656 3200 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 5540 12588 5592 12640
rect 9956 12588 10008 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 11888 12588 11940 12640
rect 14188 12588 14240 12640
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 3240 12384 3292 12436
rect 4712 12384 4764 12436
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 6920 12384 6972 12436
rect 3332 12248 3384 12300
rect 3424 12248 3476 12300
rect 5356 12248 5408 12300
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 9404 12384 9456 12436
rect 5632 12248 5684 12257
rect 940 12180 992 12232
rect 2044 12180 2096 12232
rect 3056 12180 3108 12232
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3240 12112 3292 12164
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 7288 12180 7340 12232
rect 8300 12180 8352 12232
rect 6736 12112 6788 12164
rect 7656 12112 7708 12164
rect 11612 12384 11664 12436
rect 11888 12359 11940 12368
rect 11888 12325 11897 12359
rect 11897 12325 11931 12359
rect 11931 12325 11940 12359
rect 11888 12316 11940 12325
rect 14832 12316 14884 12368
rect 9956 12248 10008 12300
rect 11244 12248 11296 12300
rect 9864 12180 9916 12232
rect 10140 12180 10192 12232
rect 11796 12180 11848 12232
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 3884 12044 3936 12096
rect 5080 12044 5132 12096
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 13912 12044 13964 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 1584 11840 1636 11892
rect 3148 11840 3200 11892
rect 3240 11840 3292 11892
rect 4712 11840 4764 11892
rect 5172 11840 5224 11892
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 7656 11840 7708 11892
rect 9956 11840 10008 11892
rect 11888 11840 11940 11892
rect 940 11636 992 11688
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 3332 11636 3384 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 3516 11636 3568 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 5080 11704 5132 11756
rect 6000 11568 6052 11620
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4068 11500 4120 11552
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 10784 11704 10836 11756
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 11612 11636 11664 11688
rect 6644 11500 6696 11552
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 1676 11296 1728 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4160 11296 4212 11348
rect 3056 11092 3108 11144
rect 3332 11092 3384 11144
rect 3976 11092 4028 11144
rect 6644 11296 6696 11348
rect 6736 11296 6788 11348
rect 8392 11296 8444 11348
rect 11060 11160 11112 11212
rect 6920 11092 6972 11144
rect 7288 11092 7340 11144
rect 6000 11024 6052 11076
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 5540 10956 5592 11008
rect 6736 10999 6788 11008
rect 6736 10965 6745 10999
rect 6745 10965 6779 10999
rect 6779 10965 6788 10999
rect 6736 10956 6788 10965
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 9864 11092 9916 11144
rect 10140 11092 10192 11144
rect 10600 11092 10652 11144
rect 8668 10956 8720 11008
rect 11060 10956 11112 11008
rect 12164 10999 12216 11008
rect 12164 10965 12173 10999
rect 12173 10965 12207 10999
rect 12207 10965 12216 10999
rect 12164 10956 12216 10965
rect 13912 10956 13964 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 1032 10684 1084 10736
rect 4804 10616 4856 10668
rect 5908 10684 5960 10736
rect 7564 10684 7616 10736
rect 8484 10684 8536 10736
rect 5816 10616 5868 10668
rect 6736 10616 6788 10668
rect 7012 10616 7064 10668
rect 8300 10616 8352 10668
rect 10600 10684 10652 10736
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 10232 10659 10284 10668
rect 10232 10625 10241 10659
rect 10241 10625 10275 10659
rect 10275 10625 10284 10659
rect 10232 10616 10284 10625
rect 11060 10616 11112 10668
rect 11612 10616 11664 10668
rect 9956 10480 10008 10532
rect 11336 10480 11388 10532
rect 3424 10412 3476 10464
rect 5632 10412 5684 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 8300 10412 8352 10464
rect 8484 10412 8536 10464
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 4068 10140 4120 10192
rect 8668 10140 8720 10192
rect 11612 10183 11664 10192
rect 11612 10149 11621 10183
rect 11621 10149 11655 10183
rect 11655 10149 11664 10183
rect 11612 10140 11664 10149
rect 3148 10047 3200 10056
rect 3148 10013 3166 10047
rect 3166 10013 3200 10047
rect 3148 10004 3200 10013
rect 5724 10004 5776 10056
rect 8484 10004 8536 10056
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11336 10072 11388 10124
rect 4712 9936 4764 9988
rect 7012 9936 7064 9988
rect 7196 9936 7248 9988
rect 9864 10004 9916 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 10048 9936 10100 9988
rect 13544 9979 13596 9988
rect 13544 9945 13553 9979
rect 13553 9945 13587 9979
rect 13587 9945 13596 9979
rect 13544 9936 13596 9945
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 3148 9868 3200 9920
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 9312 9868 9364 9920
rect 9864 9868 9916 9920
rect 13728 9868 13780 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 4712 9664 4764 9716
rect 6000 9664 6052 9716
rect 1860 9528 1912 9580
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 4068 9528 4120 9580
rect 4988 9528 5040 9580
rect 3700 9460 3752 9512
rect 4160 9460 4212 9512
rect 4804 9460 4856 9512
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 5632 9528 5684 9580
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 8484 9596 8536 9648
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7840 9528 7892 9580
rect 10600 9596 10652 9648
rect 10968 9596 11020 9648
rect 10232 9528 10284 9580
rect 11612 9528 11664 9580
rect 6000 9460 6052 9512
rect 7012 9460 7064 9512
rect 7472 9392 7524 9444
rect 11704 9503 11756 9512
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 13820 9392 13872 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 3516 9324 3568 9376
rect 4344 9324 4396 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 7656 9324 7708 9376
rect 8392 9324 8444 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 1676 9120 1728 9172
rect 2228 9120 2280 9172
rect 3700 9120 3752 9172
rect 4344 9120 4396 9172
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 940 8848 992 8900
rect 3240 8916 3292 8968
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 6736 9052 6788 9104
rect 10692 9120 10744 9172
rect 9956 9052 10008 9104
rect 4988 8984 5040 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8300 8984 8352 9036
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 7104 8916 7156 8968
rect 4160 8780 4212 8832
rect 6736 8780 6788 8832
rect 6920 8780 6972 8832
rect 7840 8780 7892 8832
rect 10232 8916 10284 8968
rect 11888 9120 11940 9172
rect 9312 8891 9364 8900
rect 9312 8857 9321 8891
rect 9321 8857 9355 8891
rect 9355 8857 9364 8891
rect 9312 8848 9364 8857
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 12256 8916 12308 8968
rect 13544 9120 13596 9172
rect 14832 9052 14884 9104
rect 9864 8780 9916 8832
rect 10048 8780 10100 8832
rect 10232 8780 10284 8832
rect 10508 8780 10560 8832
rect 11612 8780 11664 8832
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 3608 8576 3660 8628
rect 2964 8483 3016 8492
rect 2964 8449 2982 8483
rect 2982 8449 3016 8483
rect 2964 8440 3016 8449
rect 4068 8576 4120 8628
rect 5908 8576 5960 8628
rect 7656 8576 7708 8628
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 3700 8372 3752 8424
rect 4896 8508 4948 8560
rect 7104 8508 7156 8560
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 11704 8576 11756 8628
rect 11888 8576 11940 8628
rect 9956 8508 10008 8560
rect 10324 8508 10376 8560
rect 10600 8508 10652 8560
rect 7656 8440 7708 8492
rect 8392 8440 8444 8492
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 4436 8304 4488 8356
rect 6828 8372 6880 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 2964 8236 3016 8288
rect 6552 8236 6604 8288
rect 8116 8236 8168 8288
rect 9128 8236 9180 8288
rect 10692 8440 10744 8492
rect 11612 8440 11664 8492
rect 12808 8440 12860 8492
rect 13820 8508 13872 8560
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10048 8372 10100 8424
rect 10784 8304 10836 8356
rect 11244 8304 11296 8356
rect 14464 8304 14516 8356
rect 10048 8236 10100 8288
rect 12624 8236 12676 8288
rect 13268 8236 13320 8288
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 1860 8032 1912 8084
rect 6644 8032 6696 8084
rect 6920 8032 6972 8084
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 8668 8032 8720 8084
rect 9956 8032 10008 8084
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 13820 8032 13872 8084
rect 3700 7964 3752 8016
rect 940 7828 992 7880
rect 3516 7896 3568 7948
rect 4712 7896 4764 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 6552 7964 6604 8016
rect 5908 7896 5960 7948
rect 7104 7896 7156 7948
rect 4344 7760 4396 7812
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 5632 7828 5684 7880
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 10048 8007 10100 8016
rect 10048 7973 10057 8007
rect 10057 7973 10091 8007
rect 10091 7973 10100 8007
rect 10048 7964 10100 7973
rect 9036 7896 9088 7948
rect 12624 8007 12676 8016
rect 12624 7973 12633 8007
rect 12633 7973 12667 8007
rect 12667 7973 12676 8007
rect 12624 7964 12676 7973
rect 11244 7896 11296 7948
rect 5264 7760 5316 7812
rect 8116 7803 8168 7812
rect 6460 7735 6512 7744
rect 6460 7701 6469 7735
rect 6469 7701 6503 7735
rect 6503 7701 6512 7735
rect 6460 7692 6512 7701
rect 8116 7769 8125 7803
rect 8125 7769 8159 7803
rect 8159 7769 8168 7803
rect 8116 7760 8168 7769
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 10508 7828 10560 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12072 7803 12124 7812
rect 12072 7769 12081 7803
rect 12081 7769 12115 7803
rect 12115 7769 12124 7803
rect 12072 7760 12124 7769
rect 8208 7692 8260 7744
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2504 7488 2556 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2412 7284 2464 7336
rect 3056 7488 3108 7540
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 6000 7488 6052 7540
rect 6920 7488 6972 7540
rect 7564 7488 7616 7540
rect 8208 7488 8260 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 9036 7531 9088 7540
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 9588 7488 9640 7540
rect 12072 7488 12124 7540
rect 3884 7420 3936 7472
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3424 7352 3476 7404
rect 4252 7352 4304 7404
rect 5356 7352 5408 7404
rect 6460 7352 6512 7404
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 13268 7488 13320 7540
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 5632 7216 5684 7268
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9864 7352 9916 7404
rect 10876 7352 10928 7404
rect 8944 7284 8996 7336
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 940 7148 992 7200
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 6460 7148 6512 7200
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 7380 7148 7432 7200
rect 7472 7148 7524 7200
rect 7840 7148 7892 7200
rect 10416 7216 10468 7268
rect 10692 7259 10744 7268
rect 10692 7225 10701 7259
rect 10701 7225 10735 7259
rect 10735 7225 10744 7259
rect 10692 7216 10744 7225
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 11244 7148 11296 7200
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 1768 6944 1820 6996
rect 3700 6944 3752 6996
rect 4160 6944 4212 6996
rect 5356 6987 5408 6996
rect 5356 6953 5365 6987
rect 5365 6953 5399 6987
rect 5399 6953 5408 6987
rect 5356 6944 5408 6953
rect 8300 6944 8352 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 2228 6808 2280 6860
rect 3792 6808 3844 6860
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 11888 6876 11940 6928
rect 14096 6876 14148 6928
rect 6736 6808 6788 6817
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2412 6740 2464 6792
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 3516 6672 3568 6724
rect 4252 6715 4304 6724
rect 4252 6681 4286 6715
rect 4286 6681 4304 6715
rect 4252 6672 4304 6681
rect 5632 6672 5684 6724
rect 6920 6672 6972 6724
rect 9312 6808 9364 6860
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 7656 6740 7708 6792
rect 7840 6672 7892 6724
rect 11244 6740 11296 6792
rect 12532 6740 12584 6792
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 4896 6604 4948 6656
rect 6644 6604 6696 6656
rect 7380 6604 7432 6656
rect 10784 6672 10836 6724
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 9220 6604 9272 6656
rect 12808 6604 12860 6656
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 940 6264 992 6316
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 3148 6264 3200 6316
rect 4252 6400 4304 6452
rect 6368 6400 6420 6452
rect 6552 6400 6604 6452
rect 6644 6400 6696 6452
rect 6920 6400 6972 6452
rect 7564 6400 7616 6452
rect 7656 6400 7708 6452
rect 8668 6400 8720 6452
rect 9864 6400 9916 6452
rect 10416 6400 10468 6452
rect 4896 6375 4948 6384
rect 3976 6196 4028 6248
rect 4896 6341 4905 6375
rect 4905 6341 4939 6375
rect 4939 6341 4948 6375
rect 4896 6332 4948 6341
rect 2136 6060 2188 6112
rect 6000 6128 6052 6180
rect 8944 6332 8996 6384
rect 12808 6332 12860 6384
rect 6736 6196 6788 6248
rect 4068 6060 4120 6112
rect 6460 6060 6512 6112
rect 8760 6264 8812 6316
rect 9220 6264 9272 6316
rect 8300 6128 8352 6180
rect 10324 6264 10376 6316
rect 10784 6264 10836 6316
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 1768 5856 1820 5908
rect 2504 5856 2556 5908
rect 3792 5856 3844 5908
rect 3976 5856 4028 5908
rect 2596 5788 2648 5840
rect 3148 5720 3200 5772
rect 3608 5720 3660 5772
rect 6092 5856 6144 5908
rect 6828 5856 6880 5908
rect 8852 5856 8904 5908
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 3700 5652 3752 5704
rect 3792 5652 3844 5704
rect 4068 5652 4120 5704
rect 8300 5720 8352 5772
rect 9312 5856 9364 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 14188 5856 14240 5908
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2596 5627 2648 5636
rect 2596 5593 2605 5627
rect 2605 5593 2639 5627
rect 2639 5593 2648 5627
rect 2596 5584 2648 5593
rect 3332 5584 3384 5636
rect 5356 5627 5408 5636
rect 5356 5593 5390 5627
rect 5390 5593 5408 5627
rect 5356 5584 5408 5593
rect 6000 5584 6052 5636
rect 7472 5584 7524 5636
rect 3240 5516 3292 5568
rect 5540 5516 5592 5568
rect 7656 5516 7708 5568
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 10600 5652 10652 5704
rect 9036 5584 9088 5636
rect 13544 5627 13596 5636
rect 13544 5593 13553 5627
rect 13553 5593 13587 5627
rect 13587 5593 13596 5627
rect 13544 5584 13596 5593
rect 15016 5584 15068 5636
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 2596 5312 2648 5364
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3608 5312 3660 5364
rect 3792 5244 3844 5296
rect 7012 5312 7064 5364
rect 5356 5287 5408 5296
rect 5356 5253 5365 5287
rect 5365 5253 5399 5287
rect 5399 5253 5408 5287
rect 5356 5244 5408 5253
rect 5540 5287 5592 5296
rect 5540 5253 5549 5287
rect 5549 5253 5583 5287
rect 5583 5253 5592 5287
rect 5540 5244 5592 5253
rect 5632 5287 5684 5296
rect 5632 5253 5641 5287
rect 5641 5253 5675 5287
rect 5675 5253 5684 5287
rect 5632 5244 5684 5253
rect 6920 5287 6972 5296
rect 6920 5253 6929 5287
rect 6929 5253 6963 5287
rect 6963 5253 6972 5287
rect 6920 5244 6972 5253
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 8024 5244 8076 5296
rect 9772 5287 9824 5296
rect 9772 5253 9781 5287
rect 9781 5253 9815 5287
rect 9815 5253 9824 5287
rect 9772 5244 9824 5253
rect 9864 5287 9916 5296
rect 9864 5253 9873 5287
rect 9873 5253 9907 5287
rect 9907 5253 9916 5287
rect 9864 5244 9916 5253
rect 10692 5287 10744 5296
rect 10692 5253 10701 5287
rect 10701 5253 10735 5287
rect 10735 5253 10744 5287
rect 10692 5244 10744 5253
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2228 5176 2280 5228
rect 8484 5176 8536 5228
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 7196 5108 7248 5160
rect 8392 5108 8444 5160
rect 940 4972 992 5024
rect 3148 4972 3200 5024
rect 4804 4972 4856 5024
rect 7656 4972 7708 5024
rect 14096 4972 14148 5024
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 3240 4768 3292 4820
rect 8024 4768 8076 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10692 4768 10744 4820
rect 13544 4768 13596 4820
rect 4160 4743 4212 4752
rect 4160 4709 4169 4743
rect 4169 4709 4203 4743
rect 4203 4709 4212 4743
rect 4160 4700 4212 4709
rect 3056 4632 3108 4684
rect 9312 4632 9364 4684
rect 2228 4564 2280 4616
rect 2320 4564 2372 4616
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4252 4564 4304 4616
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 2136 4428 2188 4480
rect 4712 4428 4764 4480
rect 5540 4428 5592 4480
rect 6736 4496 6788 4548
rect 7656 4539 7708 4548
rect 7656 4505 7690 4539
rect 7690 4505 7708 4539
rect 7656 4496 7708 4505
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 4252 4224 4304 4276
rect 4804 4224 4856 4276
rect 5448 4224 5500 4276
rect 5540 4224 5592 4276
rect 2412 4156 2464 4208
rect 1952 4088 2004 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 3700 4088 3752 4140
rect 5816 4199 5868 4208
rect 5816 4165 5825 4199
rect 5825 4165 5859 4199
rect 5859 4165 5868 4199
rect 5816 4156 5868 4165
rect 7656 4224 7708 4276
rect 8484 4224 8536 4276
rect 6736 4088 6788 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 3332 4020 3384 4072
rect 4160 4020 4212 4072
rect 4252 4063 4304 4072
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 4712 4020 4764 4072
rect 5540 4020 5592 4072
rect 8944 4020 8996 4072
rect 10508 4020 10560 4072
rect 12808 4020 12860 4072
rect 940 3884 992 3936
rect 2504 3884 2556 3936
rect 5356 3884 5408 3936
rect 7012 3884 7064 3936
rect 8760 3884 8812 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 4252 3680 4304 3732
rect 6644 3680 6696 3732
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 5908 3612 5960 3664
rect 8944 3680 8996 3732
rect 1676 3476 1728 3528
rect 940 3408 992 3460
rect 3056 3476 3108 3528
rect 3976 3544 4028 3596
rect 6920 3544 6972 3596
rect 2320 3408 2372 3460
rect 2504 3451 2556 3460
rect 2504 3417 2538 3451
rect 2538 3417 2556 3451
rect 2504 3408 2556 3417
rect 5264 3408 5316 3460
rect 6828 3476 6880 3528
rect 8852 3612 8904 3664
rect 10048 3680 10100 3732
rect 10508 3680 10560 3732
rect 10876 3612 10928 3664
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 12532 3476 12584 3528
rect 13912 3476 13964 3528
rect 11152 3408 11204 3460
rect 11796 3408 11848 3460
rect 4068 3340 4120 3392
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 1768 3136 1820 3188
rect 1952 3136 2004 3188
rect 2044 3136 2096 3188
rect 2136 3000 2188 3052
rect 2412 3000 2464 3052
rect 3332 3000 3384 3052
rect 5724 3136 5776 3188
rect 5908 3136 5960 3188
rect 4068 3068 4120 3120
rect 7380 3136 7432 3188
rect 8300 3136 8352 3188
rect 6644 3068 6696 3120
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 5356 3000 5408 3052
rect 8944 3136 8996 3188
rect 9312 3136 9364 3188
rect 10968 3136 11020 3188
rect 10692 3000 10744 3052
rect 11244 3000 11296 3052
rect 7564 2864 7616 2916
rect 11152 2932 11204 2984
rect 10140 2864 10192 2916
rect 5632 2796 5684 2848
rect 13728 3000 13780 3052
rect 15016 3000 15068 3052
rect 12900 2839 12952 2848
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 14096 2796 14148 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 2228 2592 2280 2644
rect 4712 2592 4764 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 5816 2592 5868 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 10232 2592 10284 2644
rect 11244 2592 11296 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 5908 2524 5960 2576
rect 4068 2456 4120 2508
rect 7288 2456 7340 2508
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 3424 2388 3476 2440
rect 4528 2388 4580 2440
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 5540 2388 5592 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 5632 2320 5684 2372
rect 6000 2320 6052 2372
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 8576 2388 8628 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 11152 2388 11204 2440
rect 12440 2388 12492 2440
rect 14004 2388 14056 2440
rect 14648 2388 14700 2440
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 3976 2048 4028 2100
rect 9772 2048 9824 2100
<< metal2 >>
rect 1030 19200 1086 20000
rect 2410 19200 2466 20000
rect 3790 19200 3846 20000
rect 5170 19200 5226 20000
rect 6550 19200 6606 20000
rect 7930 19200 7986 20000
rect 8036 19230 8248 19258
rect 1044 17338 1072 19200
rect 1122 17776 1178 17785
rect 1122 17711 1178 17720
rect 1136 17338 1164 17711
rect 2424 17338 2452 19200
rect 2778 18592 2834 18601
rect 2778 18527 2834 18536
rect 1032 17332 1084 17338
rect 1032 17274 1084 17280
rect 1124 17332 1176 17338
rect 1124 17274 1176 17280
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 16969 980 17138
rect 2792 17134 2820 18527
rect 3804 17338 3832 19200
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 5184 17338 5212 19200
rect 6564 17338 6592 19200
rect 7944 19122 7972 19200
rect 8036 19122 8064 19230
rect 7944 19094 8064 19122
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 8220 17338 8248 19230
rect 9310 19200 9366 20000
rect 10690 19200 10746 20000
rect 12070 19200 12126 20000
rect 13450 19200 13506 20000
rect 14568 19230 14780 19258
rect 9324 17338 9352 19200
rect 10704 17338 10732 19200
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 12084 17338 12112 19200
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 1584 16992 1636 16998
rect 938 16960 994 16969
rect 1584 16934 1636 16940
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 938 16895 994 16904
rect 1596 16794 1624 16934
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1964 16658 1992 16934
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16153 980 16458
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1032 16176 1084 16182
rect 938 16144 994 16153
rect 1032 16118 1084 16124
rect 938 16079 994 16088
rect 1044 15337 1072 16118
rect 1688 15994 1716 16390
rect 1688 15966 1808 15994
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15706 1716 15846
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1030 15328 1086 15337
rect 1030 15263 1086 15272
rect 1412 13705 1440 15438
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1596 14414 1624 15302
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1688 14074 1716 15302
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1780 13852 1808 15966
rect 2148 15502 2176 16934
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2792 16250 2820 16526
rect 3068 16250 3096 16526
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 16250 3556 16390
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 2424 15570 2452 15846
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 3160 15706 3188 15846
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 3424 15496 3476 15502
rect 3528 15484 3556 16050
rect 3608 15496 3660 15502
rect 3528 15456 3608 15484
rect 3424 15438 3476 15444
rect 3608 15438 3660 15444
rect 1872 14657 1900 15438
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2056 15026 2084 15302
rect 3068 15094 3096 15302
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1858 14648 1914 14657
rect 2056 14618 2084 14758
rect 2424 14618 2452 14894
rect 1858 14583 1914 14592
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 1780 13824 1900 13852
rect 1768 13728 1820 13734
rect 1398 13696 1454 13705
rect 1768 13670 1820 13676
rect 1398 13631 1454 13640
rect 1780 13530 1808 13670
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 12986 1440 13126
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 940 12912 992 12918
rect 938 12880 940 12889
rect 992 12880 994 12889
rect 1780 12850 1808 13466
rect 938 12815 994 12824
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 952 12073 980 12174
rect 1584 12096 1636 12102
rect 938 12064 994 12073
rect 1584 12038 1636 12044
rect 938 11999 994 12008
rect 1596 11898 1624 12038
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 940 11688 992 11694
rect 1688 11642 1716 12582
rect 1872 12434 1900 13824
rect 2056 13802 2084 14554
rect 2516 14532 2544 14962
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2688 14544 2740 14550
rect 2516 14504 2688 14532
rect 2688 14486 2740 14492
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13326 2544 13670
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 3068 13394 3096 14758
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3252 14006 3280 14214
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 940 11630 992 11636
rect 952 11257 980 11630
rect 1596 11614 1716 11642
rect 1780 12406 1900 12434
rect 938 11248 994 11257
rect 938 11183 994 11192
rect 1032 10736 1084 10742
rect 1032 10678 1084 10684
rect 1044 10441 1072 10678
rect 1030 10432 1086 10441
rect 1030 10367 1086 10376
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8809 980 8842
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 938 7984 994 7993
rect 938 7919 994 7928
rect 952 7886 980 7919
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 940 7200 992 7206
rect 938 7168 940 7177
rect 992 7168 994 7177
rect 938 7103 994 7112
rect 1596 6914 1624 11614
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9178 1716 9318
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1780 7970 1808 12406
rect 2056 12238 2084 12582
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2516 11762 2544 12786
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 3068 12238 3096 13194
rect 3160 12714 3188 13670
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12986 3372 13262
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3436 12866 3464 15438
rect 3620 15162 3648 15438
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3712 12986 3740 17002
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3896 15978 3924 16390
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3896 15366 3924 15914
rect 4172 15706 4200 17138
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4264 16182 4292 16934
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4724 16046 4752 16458
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4528 15904 4580 15910
rect 4580 15864 4660 15892
rect 4528 15846 4580 15852
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4632 15450 4660 15864
rect 4724 15706 4752 15982
rect 4816 15706 4844 16458
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4632 15422 4752 15450
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 14822 4200 15302
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14482 4200 14758
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13530 4568 13670
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3344 12838 3464 12866
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3252 12442 3280 12786
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 12306 3372 12838
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12306 3464 12582
rect 4724 12442 4752 15422
rect 4908 14482 4936 16934
rect 5644 16794 5672 17138
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 16114 5304 16390
rect 5368 16182 5396 16458
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 15094 5396 15302
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14006 4844 14214
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 5000 13938 5028 14282
rect 5092 13938 5120 14486
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5184 13818 5212 14214
rect 5092 13790 5212 13818
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12986 4936 13262
rect 5092 13258 5120 13790
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12442 4844 12718
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 3068 11150 3096 12174
rect 3160 11898 3188 12174
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3252 11898 3280 12106
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 3160 10062 3188 11494
rect 3344 11150 3372 11630
rect 3436 11354 3464 11630
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11234 3556 11630
rect 3896 11558 3924 12038
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4724 11898 4752 12378
rect 5184 12322 5212 13126
rect 5092 12294 5212 12322
rect 5368 12306 5396 14758
rect 5552 13394 5580 15846
rect 5736 15434 5764 16934
rect 5828 16658 5856 16934
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5828 15484 5856 16390
rect 5920 16250 5948 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5920 15706 5948 16186
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5908 15496 5960 15502
rect 5828 15456 5908 15484
rect 5908 15438 5960 15444
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5920 15008 5948 15438
rect 6012 15162 6040 15982
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 6472 15706 6500 15846
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6380 15162 6408 15438
rect 6564 15178 6592 16526
rect 6656 15502 6684 16934
rect 7208 16590 7236 16934
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6748 15706 6776 15982
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6840 15502 6868 16390
rect 6932 16250 6960 16390
rect 7300 16250 7328 16390
rect 7484 16250 7512 16526
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 9048 16182 9076 16934
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9876 16590 9904 16934
rect 10796 16590 10824 16934
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6472 15150 6592 15178
rect 6000 15020 6052 15026
rect 5920 14980 6000 15008
rect 6000 14962 6052 14968
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5644 14346 5672 14894
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5644 13938 5672 14282
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12322 5580 12582
rect 5644 12434 5672 13874
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 13530 5856 13670
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5724 13320 5776 13326
rect 5776 13280 5856 13308
rect 5724 13262 5776 13268
rect 5644 12406 5764 12434
rect 5552 12306 5672 12322
rect 5356 12300 5408 12306
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3436 11206 3556 11234
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3436 10470 3464 11206
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1872 8634 1900 9522
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9178 2268 9318
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1872 8090 1900 8570
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 8294 3004 8434
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1780 7942 1900 7970
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 7002 1808 7346
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1596 6886 1716 6914
rect 938 6352 994 6361
rect 938 6287 940 6296
rect 992 6287 994 6296
rect 940 6258 992 6264
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4729 980 4966
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 3936 992 3942
rect 938 3904 940 3913
rect 992 3904 994 3913
rect 938 3839 994 3848
rect 1688 3534 1716 6886
rect 1872 6866 1900 7942
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7546 2544 7686
rect 3068 7546 3096 7822
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3160 7410 3188 9862
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8430 3280 8910
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3436 7410 3464 10406
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 7954 3556 9318
rect 3620 8634 3648 9522
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3712 9178 3740 9454
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 8022 3740 8366
rect 3700 8016 3752 8022
rect 3752 7976 3832 8004
rect 3700 7958 3752 7964
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 2228 7336 2280 7342
rect 2412 7336 2464 7342
rect 2228 7278 2280 7284
rect 2332 7284 2412 7290
rect 2332 7278 2464 7284
rect 2240 6866 2268 7278
rect 2332 7262 2452 7278
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 6458 2084 6734
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1780 5914 1808 6258
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 2148 5710 2176 6054
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 1780 3194 1808 5170
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1964 3194 1992 4082
rect 2056 3194 2084 5170
rect 2240 4622 2268 5170
rect 2332 4622 2360 7262
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2424 6458 2452 6734
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2516 5914 2544 6598
rect 3160 6322 3188 7346
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 6458 3372 6734
rect 3528 6730 3556 7686
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3712 7002 3740 7278
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3804 6866 3832 7976
rect 3896 7478 3924 11494
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2596 5840 2648 5846
rect 2424 5788 2596 5794
rect 2424 5782 2648 5788
rect 2424 5766 2636 5782
rect 3160 5778 3188 6258
rect 3804 5914 3832 6802
rect 3988 6254 4016 11086
rect 4080 10198 4108 11494
rect 4172 11354 4200 11630
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4080 9586 4108 10134
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4724 9722 4752 9930
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4816 9518 4844 10610
rect 5000 9586 5028 12174
rect 5092 12102 5120 12294
rect 5552 12300 5684 12306
rect 5552 12294 5632 12300
rect 5356 12242 5408 12248
rect 5632 12242 5684 12248
rect 5736 12238 5764 12406
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11762 5120 12038
rect 5184 11898 5212 12174
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 9586 5580 10950
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 9586 5672 10406
rect 5736 10062 5764 12174
rect 5828 10674 5856 13280
rect 5920 12850 5948 14554
rect 6012 14278 6040 14962
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12986 6224 13126
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5920 10742 5948 12786
rect 6012 11626 6040 12786
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6012 11082 6040 11562
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 6012 9722 6040 10406
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4804 9512 4856 9518
rect 6000 9512 6052 9518
rect 4856 9472 4936 9500
rect 4804 9454 4856 9460
rect 4172 8922 4200 9454
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4356 9178 4384 9318
rect 4724 9178 4752 9318
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4080 8894 4200 8922
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4080 8634 4108 8894
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4172 7426 4200 8774
rect 4264 7546 4292 8910
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4908 8566 4936 9472
rect 6000 9454 6052 9460
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5000 8430 5028 8978
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4436 8356 4488 8362
rect 4356 8316 4436 8344
rect 4356 7818 4384 8316
rect 4436 8298 4488 8304
rect 4724 7954 4752 8366
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 5644 7886 5672 8910
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5920 7954 5948 8570
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 5276 7546 5304 7754
rect 6012 7546 6040 9454
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6472 8072 6500 15150
rect 6656 15094 6684 15302
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6840 14618 6868 15438
rect 7484 15434 7512 15914
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13326 6960 13874
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6656 12986 6684 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6932 12850 6960 13262
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12442 6960 12786
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11354 6684 11494
rect 6748 11354 6776 12106
rect 7208 11898 7236 14214
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12850 7328 13126
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7300 11150 7328 12174
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10674 6776 10950
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6748 8838 6776 9046
rect 6932 8838 6960 11086
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7024 9994 7052 10610
rect 7116 10606 7144 10950
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7024 9518 7052 9930
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6380 8044 6500 8072
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 4172 7410 4292 7426
rect 4172 7404 4304 7410
rect 4172 7398 4252 7404
rect 4252 7346 4304 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 7002 4200 7142
rect 5368 7002 5396 7346
rect 6380 7342 6408 8044
rect 6564 8022 6592 8230
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6656 7886 6684 8026
rect 6748 7886 6776 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6472 7410 6500 7686
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5644 6730 5672 7210
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 4264 6458 4292 6666
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4908 6390 4936 6598
rect 6380 6458 6408 6734
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5914 4016 6190
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3148 5772 3200 5778
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4146 2176 4422
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 938 3088 994 3097
rect 2148 3058 2176 4082
rect 938 3023 994 3032
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2240 2650 2268 4558
rect 2424 4298 2452 5766
rect 3148 5714 3200 5720
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 2608 5370 2636 5578
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 3068 4690 3096 5306
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2332 4270 2452 4298
rect 2332 3466 2360 4270
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2424 3058 2452 4150
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2516 3466 2544 3878
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 3068 3534 3096 4626
rect 3160 4622 3188 4966
rect 3252 4826 3280 5510
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3344 4078 3372 5578
rect 3620 5370 3648 5714
rect 4080 5710 4108 6054
rect 6012 5896 6040 6122
rect 6472 6118 6500 7142
rect 6564 6458 6592 7278
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 6458 6684 6598
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6254 6776 6802
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6840 5914 6868 8366
rect 6932 8090 6960 8774
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6932 7546 6960 8026
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 6730 6960 7142
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6458 6960 6666
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6092 5908 6144 5914
rect 6012 5868 6092 5896
rect 6092 5850 6144 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3712 4146 3740 5646
rect 3804 5302 3832 5646
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 5368 5302 5396 5578
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5302 5580 5510
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 3804 4622 3832 5238
rect 4712 5160 4764 5166
rect 5644 5114 5672 5238
rect 4712 5102 4764 5108
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 4172 4078 4200 4694
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4282 4292 4558
rect 4724 4486 4752 5102
rect 5460 5086 5672 5114
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4816 4282 4844 4966
rect 5460 4282 5488 5086
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 3344 3058 3372 4014
rect 4264 3738 4292 4014
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3988 3058 4016 3538
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3126 4108 3334
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 4724 2650 4752 4014
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 2650 5304 3402
rect 5368 3058 5396 3878
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 2240 1306 2268 2382
rect 2148 1278 2268 1306
rect 2148 800 2176 1278
rect 3436 800 3464 2382
rect 3976 2304 4028 2310
rect 4080 2281 4108 2450
rect 5552 2446 5580 4014
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4528 2440 4580 2446
rect 5540 2440 5592 2446
rect 4580 2400 4752 2428
rect 4528 2382 4580 2388
rect 3976 2246 4028 2252
rect 4066 2272 4122 2281
rect 3988 2106 4016 2246
rect 4066 2207 4122 2216
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4724 800 4752 2400
rect 5540 2382 5592 2388
rect 5644 2378 5672 2790
rect 5736 2428 5764 3130
rect 5828 2650 5856 4150
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3194 5948 3606
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6012 2774 6040 5578
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6656 3738 6684 4558
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6748 4146 6776 4490
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6656 3126 6684 3674
rect 6840 3534 6868 5850
rect 7024 5370 7052 9454
rect 7208 9178 7236 9930
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8566 7144 8910
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7116 7954 7144 8502
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 8090 7236 8366
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4570 6960 5238
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 6932 4542 7052 4570
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 3602 6960 4422
rect 7024 3942 7052 4542
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7208 3738 7236 5102
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 5920 2746 6040 2774
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2582 5948 2746
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 7300 2514 7328 9522
rect 7484 9450 7512 15370
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 8312 15162 8340 15370
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7852 14618 7880 14962
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 8128 14482 8156 14894
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8312 14414 8340 14758
rect 8496 14618 8524 16118
rect 9048 15502 9076 16118
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15094 8984 15302
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13258 7880 13670
rect 8312 13394 8340 13874
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 8312 12986 8340 13330
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12238 8340 12922
rect 8496 12850 8524 14418
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12850 8800 13126
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11898 7696 12106
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8404 11354 8432 11698
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7576 7546 7604 10678
rect 8312 10674 8340 10950
rect 8496 10742 8524 11086
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8634 7696 9318
rect 7852 9042 7880 9522
rect 8312 9042 8340 10406
rect 8496 10062 8524 10406
rect 8680 10198 8708 10950
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9654 8524 9862
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7852 8838 7880 8978
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 8404 8498 8432 9318
rect 8864 8498 8892 14962
rect 9140 14414 9168 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15026 9720 15302
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9876 14618 9904 15438
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 15094 10088 15302
rect 10152 15162 10180 16050
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15706 10364 15846
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10612 15586 10640 16526
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16182 10732 16390
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10796 15706 10824 15982
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10612 15558 10732 15586
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 10152 14414 10180 15098
rect 10428 15026 10456 15438
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10520 14618 10548 14894
rect 10612 14618 10640 15438
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 9128 14408 9180 14414
rect 10140 14408 10192 14414
rect 9128 14350 9180 14356
rect 10060 14368 10140 14396
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12986 9168 13194
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9324 12322 9352 12854
rect 9416 12442 9444 13330
rect 9876 12918 9904 13670
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9968 12782 9996 13942
rect 10060 13394 10088 14368
rect 10140 14350 10192 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 14006 10272 14350
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10704 13870 10732 15558
rect 11072 15502 11100 15846
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10140 13864 10192 13870
rect 10692 13864 10744 13870
rect 10140 13806 10192 13812
rect 10520 13824 10692 13852
rect 10152 13530 10180 13806
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9968 12646 9996 12718
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9324 12294 9904 12322
rect 9968 12306 9996 12582
rect 9876 12238 9904 12294
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10152 12238 10180 12582
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 9876 11150 9904 12174
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11898 9996 12038
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9876 10062 9904 11086
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9324 8906 9352 9862
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9876 8838 9904 9862
rect 9968 9110 9996 10474
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 9722 10088 9930
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9968 8566 9996 9046
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 7668 8090 7696 8434
rect 10060 8430 10088 8774
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8128 7818 8156 8230
rect 8680 8090 8708 8366
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 8220 7546 8248 7686
rect 8588 7546 8616 7822
rect 9048 7546 9076 7890
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9140 7410 9168 8230
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9968 8090 9996 8366
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 8022 10088 8230
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7546 9628 7822
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7392 6662 7420 7142
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 5522 7420 6598
rect 7484 5642 7512 7142
rect 7576 6458 7604 7278
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6458 7696 6734
rect 7852 6730 7880 7142
rect 8312 7002 8340 7142
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 8680 6458 8708 6598
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8956 6390 8984 7278
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5778 8340 6122
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7656 5568 7708 5574
rect 7392 5494 7512 5522
rect 7656 5510 7708 5516
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3194 7420 3334
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7484 2774 7512 5494
rect 7668 5030 7696 5510
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 8036 4826 8064 5238
rect 8404 5166 8432 5646
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7668 4282 7696 4490
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 8496 4282 8524 5170
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8772 4146 8800 6258
rect 8852 5908 8904 5914
rect 8956 5896 8984 6326
rect 8904 5868 8984 5896
rect 8852 5850 8904 5856
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 4826 9076 5578
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8772 3942 8800 4082
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3670 8892 3878
rect 8956 3738 8984 4014
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7576 2922 7604 3470
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 8312 3194 8340 3334
rect 8956 3194 8984 3334
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7484 2746 7604 2774
rect 7576 2650 7604 2746
rect 9140 2650 9168 7346
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6866 9352 7278
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9876 7002 9904 7346
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6322 9260 6598
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9324 5914 9352 6802
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9312 5908 9364 5914
rect 9876 5896 9904 6394
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9312 5850 9364 5856
rect 9784 5868 9904 5896
rect 9324 5370 9352 5850
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9324 4690 9352 5306
rect 9784 5302 9812 5868
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9876 4826 9904 5238
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9324 3194 9352 4626
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 10060 3738 10088 6190
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 9128 2644 9180 2650
rect 9876 2632 9904 3470
rect 10152 2922 10180 11086
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 9586 10272 10610
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 8974 10272 9522
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10244 2650 10272 8774
rect 10336 8566 10364 10406
rect 10520 10130 10548 13824
rect 10692 13806 10744 13812
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 11150 10640 13126
rect 10888 12782 10916 13262
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10612 9654 10640 10678
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10428 7274 10456 9318
rect 10704 9178 10732 9998
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10690 8936 10746 8945
rect 10690 8871 10746 8880
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 7886 10548 8774
rect 10704 8634 10732 8871
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10428 6458 10456 7210
rect 10612 6866 10640 8502
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 7274 10732 8434
rect 10796 8362 10824 11698
rect 11072 11218 11100 15438
rect 11164 15162 11192 17070
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12176 16794 12204 16934
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 13280 16794 13308 16934
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13372 16590 13400 16662
rect 13464 16590 13492 19200
rect 14462 17776 14518 17785
rect 14462 17711 14518 17720
rect 14476 17338 14504 17711
rect 14568 17338 14596 19230
rect 14752 19122 14780 19230
rect 14830 19200 14886 20000
rect 14844 19122 14872 19200
rect 14752 19094 14872 19122
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11164 13530 11192 14282
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11256 13410 11284 13670
rect 11716 13530 11744 13806
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11164 13382 11284 13410
rect 12084 13394 12112 14962
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12176 14414 12204 14758
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11612 13388 11664 13394
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10674 11100 10950
rect 11164 10690 11192 13382
rect 11612 13330 11664 13336
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12306 11284 12582
rect 11624 12442 11652 13330
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12986 11928 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12176 12918 12204 14350
rect 12452 14278 12480 14758
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11900 12374 11928 12582
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11060 10668 11112 10674
rect 11164 10662 11284 10690
rect 11624 10674 11652 11630
rect 11060 10610 11112 10616
rect 11256 10130 11284 10662
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 10130 11376 10474
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 8974 11008 9590
rect 11624 9586 11652 10134
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 10968 8968 11020 8974
rect 10888 8916 10968 8922
rect 10888 8910 11020 8916
rect 10888 8894 11008 8910
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10888 7410 10916 8894
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11624 8498 11652 8774
rect 11716 8634 11744 9454
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 7954 11284 8298
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10888 6746 10916 7346
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6798 11284 7142
rect 10796 6730 10916 6746
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10784 6724 10916 6730
rect 10836 6718 10916 6724
rect 10784 6666 10836 6672
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10796 6322 10824 6666
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10336 5914 10364 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10612 4690 10640 5646
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10704 4826 10732 5238
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10520 3738 10548 4014
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10888 3670 10916 4558
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 11808 3466 11836 12174
rect 11900 11898 11928 12310
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10810 12204 10950
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12176 10062 12204 10746
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11900 8634 11928 9114
rect 12268 8974 12296 9454
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 6934 11928 7822
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7546 12112 7754
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 12544 6798 12572 16390
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14074 12664 14350
rect 12728 14074 12756 14894
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12820 14618 12848 14758
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13280 14006 13308 14758
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13530 12756 13806
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 13372 13326 13400 15030
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13464 14074 13492 14350
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13740 13938 13768 15302
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 13556 9178 13584 9930
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9625 13768 9862
rect 13726 9616 13782 9625
rect 13726 9551 13782 9560
rect 13832 9450 13860 16390
rect 13924 16250 13952 16526
rect 14016 16250 14044 17138
rect 14108 16522 14136 17138
rect 14372 16992 14424 16998
rect 14370 16960 14372 16969
rect 14424 16960 14426 16969
rect 14370 16895 14426 16904
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14384 16153 14412 16390
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14844 15473 14872 15574
rect 14830 15464 14886 15473
rect 14830 15399 14886 15408
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14200 14618 14228 14962
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14384 14521 14412 14758
rect 14370 14512 14426 14521
rect 14370 14447 14426 14456
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13705 14504 13806
rect 14462 13696 14518 13705
rect 14462 13631 14518 13640
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12889 14412 13126
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12238 14228 12582
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14188 12232 14240 12238
rect 14844 12209 14872 12310
rect 14188 12174 14240 12180
rect 14830 12200 14886 12209
rect 14830 12135 14886 12144
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11762 13952 12038
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11257 14412 11494
rect 14370 11248 14426 11257
rect 14370 11183 14426 11192
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8022 12664 8230
rect 12820 8090 12848 8434
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 13280 7546 13308 8230
rect 13832 8090 13860 8502
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6390 12848 6598
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12820 4078 12848 6326
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 13556 4826 13584 5578
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12820 3618 12848 4014
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 12820 3590 12940 3618
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 10968 3188 11020 3194
rect 10704 3148 10968 3176
rect 10704 3058 10732 3148
rect 10968 3130 11020 3136
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 11164 2990 11192 3402
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11256 2650 11284 2994
rect 12544 2650 12572 3470
rect 12912 2854 12940 3590
rect 13924 3534 13952 10950
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14372 10464 14424 10470
rect 14370 10432 14372 10441
rect 14424 10432 14426 10441
rect 14370 10367 14426 10376
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14188 8968 14240 8974
rect 14186 8936 14188 8945
rect 14844 8945 14872 9046
rect 14240 8936 14242 8945
rect 14186 8871 14242 8880
rect 14830 8936 14886 8945
rect 14830 8871 14886 8880
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14108 6934 14136 8434
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 7993 14504 8298
rect 14462 7984 14518 7993
rect 14462 7919 14518 7928
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14372 7200 14424 7206
rect 14370 7168 14372 7177
rect 14424 7168 14426 7177
rect 14370 7103 14426 7112
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 5914 14228 6734
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6361 14412 6598
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14370 6352 14426 6361
rect 14370 6287 14426 6296
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 15014 5672 15070 5681
rect 15014 5607 15016 5616
rect 15068 5607 15070 5616
rect 15016 5578 15068 5584
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14108 4622 14136 4966
rect 14384 4729 14412 4966
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4146 14228 4422
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14372 3936 14424 3942
rect 14370 3904 14372 3913
rect 14424 3904 14426 3913
rect 14370 3839 14426 3848
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 3097 14412 3334
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14370 3088 14426 3097
rect 13728 3052 13780 3058
rect 14370 3023 14426 3032
rect 15016 3052 15068 3058
rect 13728 2994 13780 3000
rect 15016 2994 15068 3000
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 13740 2650 13768 2994
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14108 2650 14136 2790
rect 9128 2586 9180 2592
rect 9784 2604 9904 2632
rect 10232 2644 10284 2650
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 5816 2440 5868 2446
rect 5736 2400 5816 2428
rect 5816 2382 5868 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 800 6040 2314
rect 7392 1306 7420 2382
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 7300 1278 7420 1306
rect 7300 800 7328 1278
rect 8588 800 8616 2382
rect 9784 2106 9812 2604
rect 10232 2586 10284 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 9956 2440 10008 2446
rect 9876 2400 9956 2428
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9876 800 9904 2400
rect 9956 2382 10008 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14004 2440 14056 2446
rect 14648 2440 14700 2446
rect 14004 2382 14056 2388
rect 14646 2408 14648 2417
rect 14700 2408 14702 2417
rect 11164 800 11192 2382
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 12452 800 12480 2382
rect 14016 1442 14044 2382
rect 14646 2343 14702 2352
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 13740 1414 14044 1442
rect 13740 800 13768 1414
rect 15028 800 15056 2994
rect 2134 0 2190 800
rect 3422 0 3478 800
rect 4710 0 4766 800
rect 5998 0 6054 800
rect 7286 0 7342 800
rect 8574 0 8630 800
rect 9862 0 9918 800
rect 11150 0 11206 800
rect 12438 0 12494 800
rect 13726 0 13782 800
rect 15014 0 15070 800
<< via2 >>
rect 1122 17720 1178 17776
rect 2778 18536 2834 18592
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 938 16904 994 16960
rect 938 16088 994 16144
rect 1030 15272 1086 15328
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 1858 14592 1914 14648
rect 1398 13640 1454 13696
rect 938 12860 940 12880
rect 940 12860 992 12880
rect 992 12860 994 12880
rect 938 12824 994 12860
rect 938 12008 994 12064
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 938 11192 994 11248
rect 1030 10376 1086 10432
rect 1490 9560 1546 9616
rect 938 8744 994 8800
rect 938 7928 994 7984
rect 938 7148 940 7168
rect 940 7148 992 7168
rect 992 7148 994 7168
rect 938 7112 994 7148
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 938 6316 994 6352
rect 938 6296 940 6316
rect 940 6296 992 6316
rect 992 6296 994 6316
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 938 4664 994 4720
rect 938 3884 940 3904
rect 940 3884 992 3904
rect 992 3884 994 3904
rect 938 3848 994 3884
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 938 3032 994 3088
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4066 2216 4122 2272
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 10690 8880 10746 8936
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 14462 17720 14518 17776
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 13726 9560 13782 9616
rect 14370 16940 14372 16960
rect 14372 16940 14424 16960
rect 14424 16940 14426 16960
rect 14370 16904 14426 16940
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14370 16088 14426 16144
rect 14830 15408 14886 15464
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14370 14456 14426 14512
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14462 13640 14518 13696
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14370 12824 14426 12880
rect 14830 12144 14886 12200
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14370 11192 14426 11248
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14370 10412 14372 10432
rect 14372 10412 14424 10432
rect 14424 10412 14426 10432
rect 14370 10376 14426 10412
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14186 8916 14188 8936
rect 14188 8916 14240 8936
rect 14240 8916 14242 8936
rect 14186 8880 14242 8916
rect 14830 8880 14886 8936
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14462 7928 14518 7984
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14370 7148 14372 7168
rect 14372 7148 14424 7168
rect 14424 7148 14426 7168
rect 14370 7112 14426 7148
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14370 6296 14426 6352
rect 15014 5636 15070 5672
rect 15014 5616 15016 5636
rect 15016 5616 15068 5636
rect 15068 5616 15070 5636
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14370 4664 14426 4720
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14370 3884 14372 3904
rect 14372 3884 14424 3904
rect 14424 3884 14426 3904
rect 14370 3848 14426 3884
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 14370 3032 14426 3088
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 14646 2388 14648 2408
rect 14648 2388 14700 2408
rect 14700 2388 14702 2408
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14646 2352 14702 2388
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
<< metal3 >>
rect 0 18594 800 18624
rect 2773 18594 2839 18597
rect 0 18592 2839 18594
rect 0 18536 2778 18592
rect 2834 18536 2839 18592
rect 0 18534 2839 18536
rect 0 18504 800 18534
rect 2773 18531 2839 18534
rect 0 17778 800 17808
rect 1117 17778 1183 17781
rect 0 17776 1183 17778
rect 0 17720 1122 17776
rect 1178 17720 1183 17776
rect 0 17718 1183 17720
rect 0 17688 800 17718
rect 1117 17715 1183 17718
rect 14457 17778 14523 17781
rect 15200 17778 16000 17808
rect 14457 17776 16000 17778
rect 14457 17720 14462 17776
rect 14518 17720 16000 17776
rect 14457 17718 16000 17720
rect 14457 17715 14523 17718
rect 15200 17688 16000 17718
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 0 16962 800 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 800 16902
rect 933 16899 999 16902
rect 14365 16962 14431 16965
rect 15200 16962 16000 16992
rect 14365 16960 16000 16962
rect 14365 16904 14370 16960
rect 14426 16904 16000 16960
rect 14365 16902 16000 16904
rect 14365 16899 14431 16902
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 15200 16872 16000 16902
rect 12940 16831 13256 16832
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 14365 16146 14431 16149
rect 15200 16146 16000 16176
rect 14365 16144 16000 16146
rect 14365 16088 14370 16144
rect 14426 16088 16000 16144
rect 14365 16086 16000 16088
rect 14365 16083 14431 16086
rect 15200 16056 16000 16086
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 14825 15466 14891 15469
rect 14825 15464 15210 15466
rect 14825 15408 14830 15464
rect 14886 15408 15210 15464
rect 14825 15406 15210 15408
rect 14825 15403 14891 15406
rect 15150 15360 15210 15406
rect 0 15330 800 15360
rect 1025 15330 1091 15333
rect 0 15328 1091 15330
rect 0 15272 1030 15328
rect 1086 15272 1091 15328
rect 0 15270 1091 15272
rect 15150 15270 16000 15360
rect 0 15240 800 15270
rect 1025 15267 1091 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 15200 15240 16000 15270
rect 14653 15199 14969 15200
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 1853 14650 1919 14653
rect 936 14648 1919 14650
rect 936 14592 1858 14648
rect 1914 14592 1919 14648
rect 936 14590 1919 14592
rect 0 14514 800 14544
rect 936 14514 996 14590
rect 1853 14587 1919 14590
rect 0 14454 996 14514
rect 14365 14514 14431 14517
rect 15200 14514 16000 14544
rect 14365 14512 16000 14514
rect 14365 14456 14370 14512
rect 14426 14456 16000 14512
rect 14365 14454 16000 14456
rect 0 14424 800 14454
rect 14365 14451 14431 14454
rect 15200 14424 16000 14454
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 14457 13698 14523 13701
rect 15200 13698 16000 13728
rect 14457 13696 16000 13698
rect 14457 13640 14462 13696
rect 14518 13640 16000 13696
rect 14457 13638 16000 13640
rect 14457 13635 14523 13638
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 15200 13608 16000 13638
rect 12940 13567 13256 13568
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 14365 12882 14431 12885
rect 15200 12882 16000 12912
rect 14365 12880 16000 12882
rect 14365 12824 14370 12880
rect 14426 12824 16000 12880
rect 14365 12822 16000 12824
rect 14365 12819 14431 12822
rect 15200 12792 16000 12822
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 14825 12202 14891 12205
rect 14825 12200 15210 12202
rect 14825 12144 14830 12200
rect 14886 12144 15210 12200
rect 14825 12142 15210 12144
rect 14825 12139 14891 12142
rect 15150 12096 15210 12142
rect 0 12066 800 12096
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 15150 12006 16000 12096
rect 0 11976 800 12006
rect 933 12003 999 12006
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 15200 11976 16000 12006
rect 14653 11935 14969 11936
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 0 11250 800 11280
rect 933 11250 999 11253
rect 0 11248 999 11250
rect 0 11192 938 11248
rect 994 11192 999 11248
rect 0 11190 999 11192
rect 0 11160 800 11190
rect 933 11187 999 11190
rect 14365 11250 14431 11253
rect 15200 11250 16000 11280
rect 14365 11248 16000 11250
rect 14365 11192 14370 11248
rect 14426 11192 16000 11248
rect 14365 11190 16000 11192
rect 14365 11187 14431 11190
rect 15200 11160 16000 11190
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 0 10434 800 10464
rect 1025 10434 1091 10437
rect 0 10432 1091 10434
rect 0 10376 1030 10432
rect 1086 10376 1091 10432
rect 0 10374 1091 10376
rect 0 10344 800 10374
rect 1025 10371 1091 10374
rect 14365 10434 14431 10437
rect 15200 10434 16000 10464
rect 14365 10432 16000 10434
rect 14365 10376 14370 10432
rect 14426 10376 16000 10432
rect 14365 10374 16000 10376
rect 14365 10371 14431 10374
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 15200 10344 16000 10374
rect 12940 10303 13256 10304
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 13721 9618 13787 9621
rect 15200 9618 16000 9648
rect 13721 9616 16000 9618
rect 13721 9560 13726 9616
rect 13782 9560 16000 9616
rect 13721 9558 16000 9560
rect 13721 9555 13787 9558
rect 15200 9528 16000 9558
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 10685 8938 10751 8941
rect 14181 8938 14247 8941
rect 10685 8936 14247 8938
rect 10685 8880 10690 8936
rect 10746 8880 14186 8936
rect 14242 8880 14247 8936
rect 10685 8878 14247 8880
rect 10685 8875 10751 8878
rect 14181 8875 14247 8878
rect 14825 8938 14891 8941
rect 14825 8936 15210 8938
rect 14825 8880 14830 8936
rect 14886 8880 15210 8936
rect 14825 8878 15210 8880
rect 14825 8875 14891 8878
rect 15150 8832 15210 8878
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 15150 8742 16000 8832
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 15200 8712 16000 8742
rect 14653 8671 14969 8672
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 0 7986 800 8016
rect 933 7986 999 7989
rect 0 7984 999 7986
rect 0 7928 938 7984
rect 994 7928 999 7984
rect 0 7926 999 7928
rect 0 7896 800 7926
rect 933 7923 999 7926
rect 14457 7986 14523 7989
rect 15200 7986 16000 8016
rect 14457 7984 16000 7986
rect 14457 7928 14462 7984
rect 14518 7928 16000 7984
rect 14457 7926 16000 7928
rect 14457 7923 14523 7926
rect 15200 7896 16000 7926
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 0 7170 800 7200
rect 933 7170 999 7173
rect 0 7168 999 7170
rect 0 7112 938 7168
rect 994 7112 999 7168
rect 0 7110 999 7112
rect 0 7080 800 7110
rect 933 7107 999 7110
rect 14365 7170 14431 7173
rect 15200 7170 16000 7200
rect 14365 7168 16000 7170
rect 14365 7112 14370 7168
rect 14426 7112 16000 7168
rect 14365 7110 16000 7112
rect 14365 7107 14431 7110
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 15200 7080 16000 7110
rect 12940 7039 13256 7040
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 14365 6354 14431 6357
rect 15200 6354 16000 6384
rect 14365 6352 16000 6354
rect 14365 6296 14370 6352
rect 14426 6296 16000 6352
rect 14365 6294 16000 6296
rect 14365 6291 14431 6294
rect 15200 6264 16000 6294
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 15009 5674 15075 5677
rect 15009 5672 15210 5674
rect 15009 5616 15014 5672
rect 15070 5616 15210 5672
rect 15009 5614 15210 5616
rect 15009 5611 15075 5614
rect 15150 5568 15210 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 15150 5478 16000 5568
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 15200 5448 16000 5478
rect 14653 5407 14969 5408
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 14365 4722 14431 4725
rect 15200 4722 16000 4752
rect 14365 4720 16000 4722
rect 14365 4664 14370 4720
rect 14426 4664 16000 4720
rect 14365 4662 16000 4664
rect 14365 4659 14431 4662
rect 15200 4632 16000 4662
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 14365 3906 14431 3909
rect 15200 3906 16000 3936
rect 14365 3904 16000 3906
rect 14365 3848 14370 3904
rect 14426 3848 16000 3904
rect 14365 3846 16000 3848
rect 14365 3843 14431 3846
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 15200 3816 16000 3846
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 14365 3090 14431 3093
rect 15200 3090 16000 3120
rect 14365 3088 16000 3090
rect 14365 3032 14370 3088
rect 14426 3032 16000 3088
rect 14365 3030 16000 3032
rect 14365 3027 14431 3030
rect 15200 3000 16000 3030
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 14641 2410 14707 2413
rect 14641 2408 15210 2410
rect 14641 2352 14646 2408
rect 14702 2352 15210 2408
rect 14641 2350 15210 2352
rect 14641 2347 14707 2350
rect 15150 2304 15210 2350
rect 0 2274 800 2304
rect 4061 2274 4127 2277
rect 0 2272 4127 2274
rect 0 2216 4066 2272
rect 4122 2216 4127 2272
rect 0 2214 4127 2216
rect 15150 2214 16000 2304
rect 0 2184 800 2214
rect 4061 2211 4127 2214
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 15200 2184 16000 2214
rect 14653 2143 14969 2144
<< via3 >>
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 16896 2977 17456
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 17440 4690 17456
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 16896 6404 17456
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 17440 8117 17456
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 16896 9831 17456
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 17440 11544 17456
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 16896 13258 17456
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 17440 14971 17456
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__inv_2  _177_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _178_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1688980957
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1688980957
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1688980957
transform 1 0 7360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1688980957
transform -1 0 6992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1688980957
transform -1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1688980957
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1688980957
transform -1 0 8096 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1688980957
transform -1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1688980957
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1688980957
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1688980957
transform -1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1688980957
transform -1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform -1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1688980957
transform -1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1688980957
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1688980957
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1688980957
transform -1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1688980957
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform -1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1688980957
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1688980957
transform -1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1688980957
transform -1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1688980957
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1688980957
transform 1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1688980957
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1688980957
transform -1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1688980957
transform -1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1688980957
transform -1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1688980957
transform 1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1688980957
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1688980957
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1688980957
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1688980957
transform -1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1688980957
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1688980957
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1688980957
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1688980957
transform -1 0 3496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1688980957
transform -1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1688980957
transform -1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1688980957
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1688980957
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1688980957
transform 1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1688980957
transform -1 0 5704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1688980957
transform -1 0 5888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1688980957
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform -1 0 3312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1688980957
transform -1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1688980957
transform -1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform -1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform -1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1688980957
transform -1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform -1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1688980957
transform -1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1688980957
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1688980957
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1688980957
transform -1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1688980957
transform -1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1688980957
transform 1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1688980957
transform -1 0 6256 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1688980957
transform -1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1688980957
transform -1 0 5520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1688980957
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1688980957
transform -1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1688980957
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1688980957
transform -1 0 13064 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1688980957
transform -1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1688980957
transform -1 0 10672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1688980957
transform 1 0 10120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1688980957
transform -1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1688980957
transform -1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1688980957
transform -1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1688980957
transform -1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1688980957
transform -1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1688980957
transform -1 0 12420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1688980957
transform -1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1688980957
transform -1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1688980957
transform -1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1688980957
transform -1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1688980957
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1688980957
transform 1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1688980957
transform -1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1688980957
transform -1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1688980957
transform -1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1688980957
transform 1 0 9016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1688980957
transform 1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1688980957
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1688980957
transform -1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1688980957
transform -1 0 6992 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1688980957
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1688980957
transform -1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1688980957
transform -1 0 5704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1688980957
transform -1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1688980957
transform -1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1688980957
transform -1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1688980957
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1688980957
transform -1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1688980957
transform -1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1688980957
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1688980957
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1688980957
transform 1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1688980957
transform 1 0 11040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1688980957
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1688980957
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1688980957
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1688980957
transform -1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1688980957
transform -1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1688980957
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1688980957
transform -1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1688980957
transform -1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1688980957
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1688980957
transform -1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1688980957
transform -1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1688980957
transform -1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1688980957
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1688980957
transform -1 0 2208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1688980957
transform -1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1688980957
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1688980957
transform -1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform -1 0 13156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1688980957
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1688980957
transform 1 0 1472 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1688980957
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1688980957
transform -1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1688980957
transform -1 0 11408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1688980957
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1688980957
transform -1 0 11316 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1688980957
transform 1 0 9384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1688980957
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1688980957
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1688980957
transform -1 0 7268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1688980957
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1688980957
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1688980957
transform -1 0 4416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1688980957
transform -1 0 2208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1688980957
transform -1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1688980957
transform -1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1688980957
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1688980957
transform -1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1688980957
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1688980957
transform -1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1688980957
transform -1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1688980957
transform -1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1688980957
transform -1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1688980957
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1688980957
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1688980957
transform -1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1688980957
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1688980957
transform -1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1688980957
transform -1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1688980957
transform -1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1688980957
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1688980957
transform -1 0 11868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1688980957
transform -1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1688980957
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1688980957
transform -1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _387_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1688980957
transform 1 0 6624 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _389_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1688980957
transform 1 0 10580 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1688980957
transform 1 0 9292 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _392_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1688980957
transform 1 0 6992 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _395_
timestamp 1688980957
transform -1 0 10488 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1688980957
transform 1 0 11040 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _398_
timestamp 1688980957
transform 1 0 8464 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1688980957
transform -1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1688980957
transform -1 0 5704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1688980957
transform -1 0 6624 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1688980957
transform -1 0 2852 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1688980957
transform -1 0 4968 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1688980957
transform -1 0 2944 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1688980957
transform -1 0 3496 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1688980957
transform 1 0 3956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1688980957
transform -1 0 6072 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1688980957
transform 1 0 3956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1688980957
transform -1 0 3312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1688980957
transform -1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1688980957
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1688980957
transform -1 0 8096 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _421_
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1688980957
transform 1 0 8096 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1688980957
transform -1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1688980957
transform -1 0 9384 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1688980957
transform -1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _441_
timestamp 1688980957
transform -1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1688980957
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _443_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1688980957
transform -1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1688980957
transform -1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _447_
timestamp 1688980957
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1688980957
transform -1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _449_
timestamp 1688980957
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _450_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _451_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _452_
timestamp 1688980957
transform 1 0 3496 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _453_
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _454_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _455_
timestamp 1688980957
transform -1 0 8648 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _455__63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _456_
timestamp 1688980957
transform 1 0 3220 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _457_
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _458_
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _459_
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _460_
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _461_
timestamp 1688980957
transform -1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _462_
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _463__64
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _463_
timestamp 1688980957
transform -1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _464_
timestamp 1688980957
transform 1 0 10580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _465_
timestamp 1688980957
transform 1 0 10488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _466_
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _467_
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _468_
timestamp 1688980957
transform 1 0 11960 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _469_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _470_
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _471_
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _472_
timestamp 1688980957
transform 1 0 9384 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _473_
timestamp 1688980957
transform -1 0 11040 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _474_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _475__65
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _475_
timestamp 1688980957
transform -1 0 8188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _476_
timestamp 1688980957
transform -1 0 8188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _477_
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _478_
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _479_
timestamp 1688980957
transform 1 0 4968 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _480_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _481_
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _482_
timestamp 1688980957
transform 1 0 7176 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _483_
timestamp 1688980957
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _484_
timestamp 1688980957
transform -1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _485_
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _486_
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _487__66
timestamp 1688980957
transform -1 0 12788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _487_
timestamp 1688980957
transform -1 0 12972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _488_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _489_
timestamp 1688980957
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _490_
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _491_
timestamp 1688980957
transform 1 0 9568 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _492_
timestamp 1688980957
transform 1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _493_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _494_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _495_
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _496_
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _497_
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _498_
timestamp 1688980957
transform 1 0 9108 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _499__67
timestamp 1688980957
transform -1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _499_
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _500_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _501_
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _502_
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _503_
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _504_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _505_
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _506_
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _507_
timestamp 1688980957
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _508_
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _509_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _509__68
timestamp 1688980957
transform -1 0 3588 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _510_
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _511_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _512_
timestamp 1688980957
transform -1 0 6624 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _513_
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _514_
timestamp 1688980957
transform 1 0 2208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _515_
timestamp 1688980957
transform -1 0 5152 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _516_
timestamp 1688980957
transform 1 0 3956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _517_
timestamp 1688980957
transform -1 0 6256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _518_
timestamp 1688980957
transform -1 0 2576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__69
timestamp 1688980957
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _519_
timestamp 1688980957
transform -1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _520_
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _521_
timestamp 1688980957
transform -1 0 3588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _522_
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _523_
timestamp 1688980957
transform -1 0 4968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _524_
timestamp 1688980957
transform 1 0 2392 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _525__70
timestamp 1688980957
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _525_
timestamp 1688980957
transform 1 0 2576 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _526_
timestamp 1688980957
transform -1 0 4508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _527_
timestamp 1688980957
transform -1 0 3680 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _528_
timestamp 1688980957
transform 1 0 1840 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _529_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _530_
timestamp 1688980957
transform -1 0 6072 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _530__71
timestamp 1688980957
transform -1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _531_
timestamp 1688980957
transform -1 0 9384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _532_
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _533_
timestamp 1688980957
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _534__72
timestamp 1688980957
transform -1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _534_
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _535_
timestamp 1688980957
transform -1 0 9568 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _536_
timestamp 1688980957
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _537_
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _538__73
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _538_
timestamp 1688980957
transform -1 0 5704 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _539_
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _540_
timestamp 1688980957
transform -1 0 6256 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _541_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _542__74
timestamp 1688980957
transform -1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _542_
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _543_
timestamp 1688980957
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _544_
timestamp 1688980957
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _545_
timestamp 1688980957
transform -1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _546_
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _546__75
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _547_
timestamp 1688980957
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _548_
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _549_
timestamp 1688980957
transform -1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _550__76
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _550_
timestamp 1688980957
transform -1 0 8556 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _551_
timestamp 1688980957
transform -1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _552_
timestamp 1688980957
transform -1 0 8372 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _553_
timestamp 1688980957
transform 1 0 6532 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _554__77
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _554_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _555_
timestamp 1688980957
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _556_
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _557_
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_43
timestamp 1688980957
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_88
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_116
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_17
timestamp 1688980957
transform 1 0 2668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_78
timestamp 1688980957
transform 1 0 8280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_103
timestamp 1688980957
transform 1 0 10580 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_107
timestamp 1688980957
transform 1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_130
timestamp 1688980957
transform 1 0 13064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_142
timestamp 1688980957
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_39
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_57
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_96
timestamp 1688980957
transform 1 0 9936 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_108
timestamp 1688980957
transform 1 0 11040 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_116
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_28
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_40
timestamp 1688980957
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_44
timestamp 1688980957
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_95
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_104
timestamp 1688980957
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_23
timestamp 1688980957
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_144
timestamp 1688980957
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_66
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_70
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_12
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_23
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_39
timestamp 1688980957
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_59
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_63
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_71
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_102
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_114
timestamp 1688980957
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_126
timestamp 1688980957
transform 1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_18
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_88
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_56
timestamp 1688980957
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_119
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_24
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_37
timestamp 1688980957
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_88
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_129
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_12
timestamp 1688980957
transform 1 0 2208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_57
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_69
timestamp 1688980957
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_88
timestamp 1688980957
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_114
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_144
timestamp 1688980957
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1688980957
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_138
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_74
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_111
timestamp 1688980957
transform 1 0 11316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_127
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_8
timestamp 1688980957
transform 1 0 1840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_20
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_46
timestamp 1688980957
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_98
timestamp 1688980957
transform 1 0 10120 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_136
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_144
timestamp 1688980957
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_9
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_145
timestamp 1688980957
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_11
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_23
timestamp 1688980957
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_35
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_102
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_124
timestamp 1688980957
transform 1 0 12512 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_136
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_8
timestamp 1688980957
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_57
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_69
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_124
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1688980957
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_67
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_80
timestamp 1688980957
transform 1 0 8464 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_92
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_99
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1688980957
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_128
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_6
timestamp 1688980957
transform 1 0 1656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_22
timestamp 1688980957
transform 1 0 3128 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_26
timestamp 1688980957
transform 1 0 3496 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_46
timestamp 1688980957
transform 1 0 5336 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_60
timestamp 1688980957
transform 1 0 6624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_97
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_124
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_136
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_144
timestamp 1688980957
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_42
timestamp 1688980957
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_74
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_94
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_107
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_24
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_95
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_132
timestamp 1688980957
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_136
timestamp 1688980957
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_21
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_89
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_107
timestamp 1688980957
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_144
timestamp 1688980957
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_17
timestamp 1688980957
transform 1 0 2668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_133
timestamp 1688980957
transform 1 0 13340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_44
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_71
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_99
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_112
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_124
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_11
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_20
timestamp 1688980957
transform 1 0 2944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_44
timestamp 1688980957
transform 1 0 5152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_79
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_90
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_101
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_144
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_11
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_17
timestamp 1688980957
transform 1 0 2668 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_50
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_60
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 1688980957
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_89
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_98
timestamp 1688980957
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_102
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_117
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_125
timestamp 1688980957
transform 1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_131
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_136
timestamp 1688980957
transform 1 0 13616 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_18
timestamp 1688980957
transform 1 0 2760 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_26
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_29
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_33
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_37
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_48
timestamp 1688980957
transform 1 0 5520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_63
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_78
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_123
timestamp 1688980957
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_129
timestamp 1688980957
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 9660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 5980 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 13524 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 10120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 4416 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 4876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 5980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 4692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 9936 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 8280 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 8832 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 10856 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 3680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 8832 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 6072 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform -1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 13340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output36 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform -1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1688980957
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1688980957
transform 1 0 14168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1688980957
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output53
timestamp 1688980957
transform -1 0 13984 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1688980957
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1688980957
transform 1 0 14168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1688980957
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1688980957
transform 1 0 14168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 0 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal input
flabel metal3 s 15200 2184 16000 2304 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 15200 3000 16000 3120 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 5 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 6 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 7 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 8 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 9 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 10 nsew signal input
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 11 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 12 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 13 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 14 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 15 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 16 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 17 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 18 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 19 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 20 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 21 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 22 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 23 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 24 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 25 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 26 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 27 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 28 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 29 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 30 nsew signal input
flabel metal3 s 15200 11160 16000 11280 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 31 nsew signal tristate
flabel metal3 s 15200 11976 16000 12096 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 32 nsew signal tristate
flabel metal3 s 15200 12792 16000 12912 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 33 nsew signal tristate
flabel metal3 s 15200 13608 16000 13728 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 34 nsew signal tristate
flabel metal3 s 15200 14424 16000 14544 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 35 nsew signal tristate
flabel metal3 s 15200 15240 16000 15360 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 36 nsew signal tristate
flabel metal3 s 15200 16056 16000 16176 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 37 nsew signal tristate
flabel metal3 s 15200 16872 16000 16992 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 38 nsew signal tristate
flabel metal3 s 15200 17688 16000 17808 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 39 nsew signal tristate
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 2410 19200 2466 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 41 nsew signal input
flabel metal2 s 3790 19200 3846 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 42 nsew signal input
flabel metal2 s 5170 19200 5226 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 43 nsew signal input
flabel metal2 s 6550 19200 6606 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 44 nsew signal input
flabel metal2 s 7930 19200 7986 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 45 nsew signal input
flabel metal2 s 9310 19200 9366 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 46 nsew signal input
flabel metal2 s 10690 19200 10746 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 47 nsew signal input
flabel metal2 s 12070 19200 12126 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 48 nsew signal input
flabel metal3 s 15200 3816 16000 3936 0 FreeSans 480 0 0 0 chany_top_out[0]
port 49 nsew signal tristate
flabel metal3 s 15200 4632 16000 4752 0 FreeSans 480 0 0 0 chany_top_out[1]
port 50 nsew signal tristate
flabel metal3 s 15200 5448 16000 5568 0 FreeSans 480 0 0 0 chany_top_out[2]
port 51 nsew signal tristate
flabel metal3 s 15200 6264 16000 6384 0 FreeSans 480 0 0 0 chany_top_out[3]
port 52 nsew signal tristate
flabel metal3 s 15200 7080 16000 7200 0 FreeSans 480 0 0 0 chany_top_out[4]
port 53 nsew signal tristate
flabel metal3 s 15200 7896 16000 8016 0 FreeSans 480 0 0 0 chany_top_out[5]
port 54 nsew signal tristate
flabel metal3 s 15200 8712 16000 8832 0 FreeSans 480 0 0 0 chany_top_out[6]
port 55 nsew signal tristate
flabel metal3 s 15200 9528 16000 9648 0 FreeSans 480 0 0 0 chany_top_out[7]
port 56 nsew signal tristate
flabel metal3 s 15200 10344 16000 10464 0 FreeSans 480 0 0 0 chany_top_out[8]
port 57 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 58 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 59 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 prog_clk
port 60 nsew signal input
flabel metal2 s 13450 19200 13506 20000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 61 nsew signal input
flabel metal2 s 14830 19200 14886 20000 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 62 nsew signal input
flabel metal4 s 2657 2128 2977 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 6084 2128 6404 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 9511 2128 9831 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 12938 2128 13258 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 4370 2128 4690 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
rlabel metal1 7958 16864 7958 16864 0 vdd
rlabel via1 8037 17408 8037 17408 0 vss
rlabel metal1 11362 15504 11362 15504 0 _000_
rlabel metal1 12466 10676 12466 10676 0 _001_
rlabel metal1 7130 16082 7130 16082 0 _002_
rlabel metal1 8004 14586 8004 14586 0 _003_
rlabel metal1 4370 7378 4370 7378 0 _004_
rlabel metal1 3772 8466 3772 8466 0 _005_
rlabel metal1 8326 7378 8326 7378 0 _006_
rlabel metal1 2438 7378 2438 7378 0 _007_
rlabel metal1 6302 6426 6302 6426 0 _008_
rlabel metal1 7590 6188 7590 6188 0 _009_
rlabel metal1 7176 2890 7176 2890 0 _010_
rlabel metal1 4876 4114 4876 4114 0 _011_
rlabel metal1 8372 3026 8372 3026 0 _012_
rlabel metal1 5796 2346 5796 2346 0 _013_
rlabel metal1 1978 3468 1978 3468 0 _014_
rlabel metal1 2116 3162 2116 3162 0 _015_
rlabel metal1 2254 6222 2254 6222 0 _016_
rlabel metal1 3680 14382 3680 14382 0 _017_
rlabel metal1 2645 12682 2645 12682 0 _018_
rlabel metal1 2806 14314 2806 14314 0 _019_
rlabel metal2 5658 16966 5658 16966 0 _020_
rlabel metal1 3220 16218 3220 16218 0 _021_
rlabel metal1 3082 12410 3082 12410 0 _022_
rlabel metal1 4140 15674 4140 15674 0 _023_
rlabel metal2 2806 16388 2806 16388 0 _024_
rlabel metal1 4324 8466 4324 8466 0 _025_
rlabel metal1 6256 7378 6256 7378 0 _026_
rlabel metal1 5290 10608 5290 10608 0 _027_
rlabel metal1 9936 8806 9936 8806 0 _028_
rlabel metal1 7452 7514 7452 7514 0 _029_
rlabel metal1 10028 14586 10028 14586 0 _030_
rlabel metal1 12466 12898 12466 12898 0 _031_
rlabel metal1 9982 11798 9982 11798 0 _032_
rlabel metal1 13156 13906 13156 13906 0 _033_
rlabel metal1 9384 13906 9384 13906 0 _034_
rlabel metal1 12696 13294 12696 13294 0 _035_
rlabel metal1 4876 11730 4876 11730 0 _036_
rlabel metal1 7912 11322 7912 11322 0 _037_
rlabel metal1 5244 11118 5244 11118 0 _038_
rlabel metal1 10488 12818 10488 12818 0 _039_
rlabel metal1 5428 13294 5428 13294 0 _040_
rlabel metal1 7176 13906 7176 13906 0 _041_
rlabel metal1 9660 6290 9660 6290 0 _042_
rlabel metal1 11408 7854 11408 7854 0 _043_
rlabel metal1 10442 7854 10442 7854 0 _044_
rlabel metal1 14030 7854 14030 7854 0 _045_
rlabel metal1 10718 8976 10718 8976 0 _046_
rlabel metal1 12558 8942 12558 8942 0 _047_
rlabel metal1 3634 6358 3634 6358 0 _048_
rlabel metal1 7820 6426 7820 6426 0 _049_
rlabel metal2 3358 6596 3358 6596 0 _050_
rlabel metal1 10304 4590 10304 4590 0 _051_
rlabel metal1 2208 11730 2208 11730 0 _052_
rlabel metal1 9062 4250 9062 4250 0 _053_
rlabel metal1 4140 5678 4140 5678 0 _054_
rlabel metal1 10626 4794 10626 4794 0 _055_
rlabel metal1 3634 6970 3634 6970 0 _056_
rlabel metal2 3174 12036 3174 12036 0 _057_
rlabel metal1 8234 6732 8234 6732 0 _058_
rlabel metal1 7958 5066 7958 5066 0 _059_
rlabel metal2 3450 11492 3450 11492 0 _060_
rlabel metal1 8740 6222 8740 6222 0 _061_
rlabel metal1 7682 6358 7682 6358 0 _062_
rlabel metal2 9890 5032 9890 5032 0 _063_
rlabel metal1 7360 6834 7360 6834 0 _064_
rlabel metal1 13018 6834 13018 6834 0 _065_
rlabel metal1 13984 8058 13984 8058 0 _066_
rlabel metal1 12144 9010 12144 9010 0 _067_
rlabel metal1 10810 7956 10810 7956 0 _068_
rlabel metal1 10626 9146 10626 9146 0 _069_
rlabel metal1 10074 8058 10074 8058 0 _070_
rlabel metal1 10258 6154 10258 6154 0 _071_
rlabel metal1 12190 7752 12190 7752 0 _072_
rlabel metal1 11454 8602 11454 8602 0 _073_
rlabel metal1 11822 7378 11822 7378 0 _074_
rlabel metal1 11408 10098 11408 10098 0 _075_
rlabel metal1 10258 7514 10258 7514 0 _076_
rlabel metal1 10994 9554 10994 9554 0 _077_
rlabel metal1 10028 12954 10028 12954 0 _078_
rlabel metal1 7682 13906 7682 13906 0 _079_
rlabel metal1 7958 11628 7958 11628 0 _080_
rlabel metal1 5796 13362 5796 13362 0 _081_
rlabel metal1 5842 11254 5842 11254 0 _082_
rlabel metal1 5060 11866 5060 11866 0 _083_
rlabel metal1 9154 12104 9154 12104 0 _084_
rlabel metal1 6762 12954 6762 12954 0 _085_
rlabel metal1 7728 12274 7728 12274 0 _086_
rlabel metal1 6118 12750 6118 12750 0 _087_
rlabel metal1 9476 11118 9476 11118 0 _088_
rlabel metal2 4830 12580 4830 12580 0 _089_
rlabel metal1 13340 14042 13340 14042 0 _090_
rlabel metal1 12834 13498 12834 13498 0 _091_
rlabel metal1 11730 12716 11730 12716 0 _092_
rlabel metal1 10856 13838 10856 13838 0 _093_
rlabel metal1 10534 11628 10534 11628 0 _094_
rlabel metal1 9752 14994 9752 14994 0 _095_
rlabel metal1 12788 14450 12788 14450 0 _096_
rlabel metal1 12006 13498 12006 13498 0 _097_
rlabel metal1 12052 14926 12052 14926 0 _098_
rlabel metal1 10488 13498 10488 13498 0 _099_
rlabel metal1 11500 12274 11500 12274 0 _100_
rlabel metal2 10534 14756 10534 14756 0 _101_
rlabel metal2 9338 9384 9338 9384 0 _102_
rlabel metal1 7820 10574 7820 10574 0 _103_
rlabel metal1 6118 7514 6118 7514 0 _104_
rlabel metal1 5750 10540 5750 10540 0 _105_
rlabel metal1 6440 7922 6440 7922 0 _106_
rlabel metal1 9384 8534 9384 8534 0 _107_
rlabel metal1 6670 10642 6670 10642 0 _108_
rlabel metal1 7958 8398 7958 8398 0 _109_
rlabel metal1 5704 9554 5704 9554 0 _110_
rlabel metal2 7682 8262 7682 8262 0 _111_
rlabel metal1 4416 16150 4416 16150 0 _112_
rlabel metal1 3496 16626 3496 16626 0 _113_
rlabel metal1 3818 16116 3818 16116 0 _114_
rlabel metal1 3726 12274 3726 12274 0 _115_
rlabel metal1 6118 16626 6118 16626 0 _116_
rlabel metal1 4554 15606 4554 15606 0 _117_
rlabel metal2 2438 15708 2438 15708 0 _118_
rlabel metal1 4048 15538 4048 15538 0 _119_
rlabel metal1 3634 11254 3634 11254 0 _120_
rlabel metal1 6072 15130 6072 15130 0 _121_
rlabel metal1 2346 13872 2346 13872 0 _122_
rlabel metal1 2392 14382 2392 14382 0 _123_
rlabel metal1 5152 13906 5152 13906 0 _124_
rlabel metal2 3358 13124 3358 13124 0 _125_
rlabel metal1 1886 14892 1886 14892 0 _126_
rlabel metal1 4738 13430 4738 13430 0 _127_
rlabel metal1 2438 5338 2438 5338 0 _128_
rlabel metal2 2438 6596 2438 6596 0 _129_
rlabel metal2 4278 3876 4278 3876 0 _130_
rlabel metal1 2208 2958 2208 2958 0 _131_
rlabel metal2 2070 6596 2070 6596 0 _132_
rlabel metal1 4462 4250 4462 4250 0 _133_
rlabel metal1 5934 2618 5934 2618 0 _134_
rlabel metal1 9154 2924 9154 2924 0 _135_
rlabel metal1 6026 3128 6026 3128 0 _136_
rlabel metal1 8970 3502 8970 3502 0 _137_
rlabel metal1 5290 4250 5290 4250 0 _138_
rlabel metal1 8372 3706 8372 3706 0 _139_
rlabel metal1 6762 3910 6762 3910 0 _140_
rlabel metal1 6854 3570 6854 3570 0 _141_
rlabel metal1 5980 6358 5980 6358 0 _142_
rlabel metal1 6762 6290 6762 6290 0 _143_
rlabel metal1 5842 6698 5842 6698 0 _144_
rlabel metal1 6532 6426 6532 6426 0 _145_
rlabel metal1 2645 7242 2645 7242 0 _146_
rlabel metal2 8602 7684 8602 7684 0 _147_
rlabel metal1 3910 7922 3910 7922 0 _148_
rlabel metal1 8878 8058 8878 8058 0 _149_
rlabel metal1 4646 8534 4646 8534 0 _150_
rlabel metal2 4278 8228 4278 8228 0 _151_
rlabel metal1 4692 8874 4692 8874 0 _152_
rlabel metal1 5106 9452 5106 9452 0 _153_
rlabel metal1 8188 15130 8188 15130 0 _154_
rlabel metal2 7498 16388 7498 16388 0 _155_
rlabel metal2 8510 15368 8510 15368 0 _156_
rlabel metal1 7130 15674 7130 15674 0 _157_
rlabel metal1 11730 10540 11730 10540 0 _158_
rlabel metal1 10994 15674 10994 15674 0 _159_
rlabel metal1 12052 11118 12052 11118 0 _160_
rlabel metal1 10718 14586 10718 14586 0 _161_
rlabel metal2 13754 1095 13754 1095 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 14766 3026 14766 3026 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 13938 2448 13938 2448 0 ccff_head
rlabel metal2 14398 3213 14398 3213 0 ccff_tail
rlabel metal3 866 10404 866 10404 0 chanx_left_in[0]
rlabel metal3 820 11220 820 11220 0 chanx_left_in[1]
rlabel metal3 820 12036 820 12036 0 chanx_left_in[2]
rlabel metal3 820 12852 820 12852 0 chanx_left_in[3]
rlabel metal3 1050 13668 1050 13668 0 chanx_left_in[4]
rlabel metal3 820 14484 820 14484 0 chanx_left_in[5]
rlabel metal3 866 15300 866 15300 0 chanx_left_in[6]
rlabel metal3 820 16116 820 16116 0 chanx_left_in[7]
rlabel metal3 820 16932 820 16932 0 chanx_left_in[8]
rlabel metal3 820 3060 820 3060 0 chanx_left_out[0]
rlabel metal3 820 3876 820 3876 0 chanx_left_out[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_out[2]
rlabel metal3 1096 5508 1096 5508 0 chanx_left_out[3]
rlabel metal3 820 6324 820 6324 0 chanx_left_out[4]
rlabel metal3 820 7140 820 7140 0 chanx_left_out[5]
rlabel metal3 820 7956 820 7956 0 chanx_left_out[6]
rlabel metal3 820 8772 820 8772 0 chanx_left_out[7]
rlabel metal3 1096 9588 1096 9588 0 chanx_left_out[8]
rlabel metal2 2162 1027 2162 1027 0 chany_bottom_in[0]
rlabel metal2 3450 1588 3450 1588 0 chany_bottom_in[1]
rlabel metal2 4738 1588 4738 1588 0 chany_bottom_in[2]
rlabel metal2 6026 1554 6026 1554 0 chany_bottom_in[3]
rlabel metal2 7314 1027 7314 1027 0 chany_bottom_in[4]
rlabel metal2 8602 1588 8602 1588 0 chany_bottom_in[5]
rlabel metal2 9890 1588 9890 1588 0 chany_bottom_in[6]
rlabel metal2 11178 1588 11178 1588 0 chany_bottom_in[7]
rlabel metal2 12466 1588 12466 1588 0 chany_bottom_in[8]
rlabel metal2 14398 11373 14398 11373 0 chany_bottom_out[0]
rlabel metal1 14628 12410 14628 12410 0 chany_bottom_out[1]
rlabel metal2 14398 13005 14398 13005 0 chany_bottom_out[2]
rlabel metal1 14444 13838 14444 13838 0 chany_bottom_out[3]
rlabel metal2 14398 14637 14398 14637 0 chany_bottom_out[4]
rlabel metal1 14628 15674 14628 15674 0 chany_bottom_out[5]
rlabel metal2 14398 16269 14398 16269 0 chany_bottom_out[6]
rlabel via2 14398 16949 14398 16949 0 chany_bottom_out[7]
rlabel metal1 14122 17306 14122 17306 0 chany_bottom_out[8]
rlabel metal1 1702 17204 1702 17204 0 chany_top_in[0]
rlabel metal1 2530 17204 2530 17204 0 chany_top_in[1]
rlabel metal1 3864 17170 3864 17170 0 chany_top_in[2]
rlabel metal1 5336 17170 5336 17170 0 chany_top_in[3]
rlabel metal1 6716 17170 6716 17170 0 chany_top_in[4]
rlabel metal1 8142 17170 8142 17170 0 chany_top_in[5]
rlabel metal1 9384 17170 9384 17170 0 chany_top_in[6]
rlabel metal1 10856 17170 10856 17170 0 chany_top_in[7]
rlabel metal1 12236 17170 12236 17170 0 chany_top_in[8]
rlabel via2 14398 3893 14398 3893 0 chany_top_out[0]
rlabel metal2 14398 4845 14398 4845 0 chany_top_out[1]
rlabel metal1 14490 5610 14490 5610 0 chany_top_out[2]
rlabel metal2 14398 6477 14398 6477 0 chany_top_out[3]
rlabel via2 14398 7157 14398 7157 0 chany_top_out[4]
rlabel metal1 14444 8330 14444 8330 0 chany_top_out[5]
rlabel metal1 14628 9146 14628 9146 0 chany_top_out[6]
rlabel metal1 13800 9894 13800 9894 0 chany_top_out[7]
rlabel via2 14398 10421 14398 10421 0 chany_top_out[8]
rlabel metal1 7866 5304 7866 5304 0 clknet_0_prog_clk
rlabel metal1 5290 7854 5290 7854 0 clknet_2_0__leaf_prog_clk
rlabel metal1 12926 8500 12926 8500 0 clknet_2_1__leaf_prog_clk
rlabel metal1 2944 13362 2944 13362 0 clknet_2_2__leaf_prog_clk
rlabel metal1 9568 14450 9568 14450 0 clknet_2_3__leaf_prog_clk
rlabel metal3 912 17748 912 17748 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 2438 17136 2438 17136 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 10212 8942 10212 8942 0 mem_bottom_track_1.DFF_0_.D
rlabel metal1 8321 11118 8321 11118 0 mem_bottom_track_1.DFF_0_.Q
rlabel metal1 7038 12410 7038 12410 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal1 8280 13362 8280 13362 0 mem_bottom_track_1.DFF_2_.Q
rlabel metal1 13018 14926 13018 14926 0 mem_bottom_track_17.DFF_0_.D
rlabel viali 2710 12206 2710 12206 0 mem_bottom_track_17.DFF_0_.Q
rlabel metal2 3634 15300 3634 15300 0 mem_bottom_track_17.DFF_1_.Q
rlabel metal2 4186 14620 4186 14620 0 mem_bottom_track_17.DFF_2_.Q
rlabel metal1 9936 12614 9936 12614 0 mem_bottom_track_9.DFF_0_.Q
rlabel metal2 12098 14178 12098 14178 0 mem_bottom_track_9.DFF_1_.Q
rlabel metal1 4646 14042 4646 14042 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 2346 12886 2346 12886 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 5428 7378 5428 7378 0 mem_left_track_11.DFF_0_.D
rlabel metal1 8050 7854 8050 7854 0 mem_left_track_11.DFF_0_.Q
rlabel metal2 1886 9078 1886 9078 0 mem_left_track_11.DFF_1_.Q
rlabel metal1 3542 9520 3542 9520 0 mem_left_track_13.DFF_0_.Q
rlabel metal1 3956 10166 3956 10166 0 mem_left_track_13.DFF_1_.Q
rlabel metal1 7038 15470 7038 15470 0 mem_left_track_15.DFF_0_.Q
rlabel metal1 8878 14382 8878 14382 0 mem_left_track_15.DFF_1_.Q
rlabel metal1 9844 15130 9844 15130 0 mem_left_track_17.DFF_0_.Q
rlabel metal1 2162 6324 2162 6324 0 mem_left_track_3.DFF_0_.Q
rlabel metal2 2162 4284 2162 4284 0 mem_left_track_3.DFF_1_.Q
rlabel metal1 4554 3468 4554 3468 0 mem_left_track_5.DFF_0_.Q
rlabel metal2 5796 2414 5796 2414 0 mem_left_track_5.DFF_1_.Q
rlabel metal1 6762 4590 6762 4590 0 mem_left_track_7.DFF_0_.Q
rlabel metal1 5106 4454 5106 4454 0 mem_left_track_7.DFF_1_.Q
rlabel metal1 6026 6222 6026 6222 0 mem_left_track_9.DFF_0_.Q
rlabel metal1 1978 11764 1978 11764 0 mem_top_track_0.DFF_0_.Q
rlabel metal1 9729 4114 9729 4114 0 mem_top_track_0.DFF_1_.Q
rlabel metal1 9614 4692 9614 4692 0 mem_top_track_0.DFF_2_.Q
rlabel metal1 13478 7854 13478 7854 0 mem_top_track_16.DFF_0_.D
rlabel metal1 10074 8840 10074 8840 0 mem_top_track_16.DFF_0_.Q
rlabel metal1 6900 11118 6900 11118 0 mem_top_track_16.DFF_1_.Q
rlabel metal1 11270 9588 11270 9588 0 mem_top_track_8.DFF_0_.Q
rlabel metal1 11362 8466 11362 8466 0 mem_top_track_8.DFF_1_.Q
rlabel metal1 4784 12818 4784 12818 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 5612 14790 5612 14790 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 10028 2890 10028 2890 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 5658 11084 5658 11084 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 2116 14246 2116 14246 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 5658 13294 5658 13294 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 5428 12614 5428 12614 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7406 11730 7406 11730 0 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 6302 13158 6302 13158 0 mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 8464 12138 8464 12138 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7820 13702 7820 13702 0 mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 13938 11900 13938 11900 0 mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 6348 16014 6348 16014 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal2 6578 15861 6578 15861 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal2 3450 8908 3450 8908 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 3818 12172 3818 12172 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 1978 15538 1978 15538 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 5750 16218 5750 16218 0 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 4692 15436 4692 15436 0 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4508 15946 4508 15946 0 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 4186 16014 4186 16014 0 mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 13271 16082 13271 16082 0 mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 10764 14994 10764 14994 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 9246 14994 9246 14994 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 11224 2890 11224 2890 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 2070 11560 2070 11560 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 1978 13838 1978 13838 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal2 10718 14705 10718 14705 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal1 10488 14858 10488 14858 0 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 11730 12614 11730 12614 0 mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 10994 13906 10994 13906 0 mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 12190 13838 12190 13838 0 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 12650 14212 12650 14212 0 mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 13432 14518 13432 14518 0 mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 5014 14110 5014 14110 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 1886 14994 1886 14994 0 mux_left_track_1.INVTX1_2_.out
rlabel metal2 4554 13600 4554 13600 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 2070 14688 2070 14688 0 mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 1794 13260 1794 13260 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9108 7922 9108 7922 0 mux_left_track_11.INVTX1_1_.out
rlabel metal1 7544 7786 7544 7786 0 mux_left_track_11.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 1794 6732 1794 6732 0 mux_left_track_11.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 6762 8466 6762 8466 0 mux_left_track_13.INVTX1_1_.out
rlabel metal2 4738 9248 4738 9248 0 mux_left_track_13.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5014 8364 5014 8364 0 mux_left_track_13.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9798 16660 9798 16660 0 mux_left_track_15.INVTX1_1_.out
rlabel metal1 7268 16218 7268 16218 0 mux_left_track_15.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 1794 9588 1794 9588 0 mux_left_track_15.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10672 16082 10672 16082 0 mux_left_track_17.INVTX1_1_.out
rlabel metal2 11086 15674 11086 15674 0 mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 12190 10880 12190 10880 0 mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 3818 5134 3818 5134 0 mux_left_track_3.INVTX1_0_.out
rlabel metal1 4692 2618 4692 2618 0 mux_left_track_3.INVTX1_1_.out
rlabel metal2 1840 7956 1840 7956 0 mux_left_track_3.INVTX1_2_.out
rlabel metal1 4140 3978 4140 3978 0 mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2530 5814 2530 5814 0 mux_left_track_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 3312 4046 3312 4046 0 mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9936 3706 9936 3706 0 mux_left_track_5.INVTX1_0_.out
rlabel metal1 10074 2958 10074 2958 0 mux_left_track_5.INVTX1_1_.out
rlabel metal1 8832 3162 8832 3162 0 mux_left_track_5.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 1794 2958 1794 2958 0 mux_left_track_5.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6808 5882 6808 5882 0 mux_left_track_7.INVTX1_0_.out
rlabel metal1 11316 3706 11316 3706 0 mux_left_track_7.INVTX1_1_.out
rlabel metal2 7222 4420 7222 4420 0 mux_left_track_7.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 5842 5100 5842 5100 0 mux_left_track_7.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6854 6834 6854 6834 0 mux_left_track_9.INVTX1_1_.out
rlabel metal1 6532 6698 6532 6698 0 mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 2162 5882 2162 5882 0 mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 12788 16422 12788 16422 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 8280 6222 8280 6222 0 mux_top_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6302 6902 6302 6902 0 mux_top_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 3910 9486 3910 9486 0 mux_top_track_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 8786 6426 8786 6426 0 mux_top_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7820 5610 7820 5610 0 mux_top_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 14122 4794 14122 4794 0 mux_top_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 7268 8398 7268 8398 0 mux_top_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6118 9690 6118 9690 0 mux_top_track_16.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 7820 8602 7820 8602 0 mux_top_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8050 10438 8050 10438 0 mux_top_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 9890 9078 9890 9078 0 mux_top_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 13846 12920 13846 12920 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 10580 6426 10580 6426 0 mux_top_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 10074 8126 10074 8126 0 mux_top_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 11408 10166 11408 10166 0 mux_top_track_8.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 12673 7446 12673 7446 0 mux_top_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13110 8568 13110 8568 0 mux_top_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 13340 8398 13340 8398 0 mux_top_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 12834 2856 12834 2856 0 net1
rlabel metal1 1840 16082 1840 16082 0 net10
rlabel metal1 7176 11254 7176 11254 0 net100
rlabel metal1 7033 8874 7033 8874 0 net101
rlabel metal2 7222 9554 7222 9554 0 net102
rlabel metal1 10248 12206 10248 12206 0 net103
rlabel metal1 2488 4590 2488 4590 0 net104
rlabel via1 3077 15062 3077 15062 0 net105
rlabel metal2 9890 7174 9890 7174 0 net106
rlabel metal1 11081 6766 11081 6766 0 net107
rlabel metal1 11316 13498 11316 13498 0 net108
rlabel metal1 7912 4250 7912 4250 0 net109
rlabel metal1 2415 16422 2415 16422 0 net11
rlabel via1 2534 13294 2534 13294 0 net110
rlabel via1 5386 15062 5386 15062 0 net111
rlabel metal1 8694 4038 8694 4038 0 net112
rlabel metal1 8648 16558 8648 16558 0 net12
rlabel metal1 2392 5202 2392 5202 0 net13
rlabel metal2 4002 2176 4002 2176 0 net14
rlabel metal1 5198 2550 5198 2550 0 net15
rlabel metal1 4738 2346 4738 2346 0 net16
rlabel metal2 7590 2689 7590 2689 0 net17
rlabel metal1 10120 8466 10120 8466 0 net18
rlabel metal1 12466 9112 12466 9112 0 net19
rlabel metal1 10350 3026 10350 3026 0 net2
rlabel metal1 11408 2618 11408 2618 0 net20
rlabel metal2 12558 3060 12558 3060 0 net21
rlabel metal1 3910 12818 3910 12818 0 net22
rlabel metal2 13386 14178 13386 14178 0 net23
rlabel metal2 13754 14620 13754 14620 0 net24
rlabel metal1 4646 14382 4646 14382 0 net25
rlabel metal1 6532 15470 6532 15470 0 net26
rlabel metal1 9108 16082 9108 16082 0 net27
rlabel metal1 9614 17000 9614 17000 0 net28
rlabel metal2 10810 16762 10810 16762 0 net29
rlabel metal2 13754 2822 13754 2822 0 net3
rlabel metal1 11822 16592 11822 16592 0 net30
rlabel metal1 1794 16592 1794 16592 0 net31
rlabel metal2 2162 16218 2162 16218 0 net32
rlabel metal1 13248 16558 13248 16558 0 net33
rlabel metal1 13754 16592 13754 16592 0 net34
rlabel metal2 13938 7242 13938 7242 0 net35
rlabel metal1 1748 3502 1748 3502 0 net36
rlabel metal1 2254 3094 2254 3094 0 net37
rlabel metal1 1748 3162 1748 3162 0 net38
rlabel metal1 1794 5576 1794 5576 0 net39
rlabel metal1 1840 10642 1840 10642 0 net4
rlabel metal1 1932 5882 1932 5882 0 net40
rlabel metal1 1748 6970 1748 6970 0 net41
rlabel metal1 1932 7786 1932 7786 0 net42
rlabel metal1 1748 8942 1748 8942 0 net43
rlabel metal1 3358 10030 3358 10030 0 net44
rlabel metal1 14122 11730 14122 11730 0 net45
rlabel metal2 14214 12410 14214 12410 0 net46
rlabel metal1 14076 13294 14076 13294 0 net47
rlabel metal1 14030 13974 14030 13974 0 net48
rlabel metal2 14214 14790 14214 14790 0 net49
rlabel metal1 1656 11118 1656 11118 0 net5
rlabel metal1 13317 15470 13317 15470 0 net50
rlabel metal2 13938 16388 13938 16388 0 net51
rlabel metal2 14122 16830 14122 16830 0 net52
rlabel metal1 14122 16218 14122 16218 0 net53
rlabel metal2 14214 4284 14214 4284 0 net54
rlabel metal1 13317 5202 13317 5202 0 net55
rlabel metal2 13570 5202 13570 5202 0 net56
rlabel metal1 14260 5882 14260 5882 0 net57
rlabel metal1 14122 7378 14122 7378 0 net58
rlabel metal2 14122 7684 14122 7684 0 net59
rlabel metal1 1518 11730 1518 11730 0 net6
rlabel metal2 10718 8755 10718 8755 0 net60
rlabel metal1 13662 9146 13662 9146 0 net61
rlabel metal1 14214 10540 14214 10540 0 net62
rlabel metal2 10626 5168 10626 5168 0 net63
rlabel metal1 12236 8942 12236 8942 0 net64
rlabel metal1 8188 13838 8188 13838 0 net65
rlabel metal1 12834 13906 12834 13906 0 net66
rlabel metal2 7130 10778 7130 10778 0 net67
rlabel metal1 3680 16558 3680 16558 0 net68
rlabel metal1 2438 14518 2438 14518 0 net69
rlabel metal1 2254 12206 2254 12206 0 net7
rlabel metal1 2438 6834 2438 6834 0 net70
rlabel metal1 5290 2414 5290 2414 0 net71
rlabel metal2 5566 5406 5566 5406 0 net72
rlabel metal1 5658 6222 5658 6222 0 net73
rlabel metal1 2852 7854 2852 7854 0 net74
rlabel metal1 4692 7922 4692 7922 0 net75
rlabel metal1 8510 15402 8510 15402 0 net76
rlabel metal1 11592 10642 11592 10642 0 net77
rlabel metal2 5382 5440 5382 5440 0 net78
rlabel via1 6665 15062 6665 15062 0 net79
rlabel metal1 1564 14382 1564 14382 0 net8
rlabel metal1 8689 15062 8689 15062 0 net80
rlabel metal1 4646 9690 4646 9690 0 net81
rlabel metal1 5857 4522 5857 4522 0 net82
rlabel via1 8781 12818 8781 12818 0 net83
rlabel metal2 9062 5202 9062 5202 0 net84
rlabel metal2 5290 7650 5290 7650 0 net85
rlabel via1 2525 3434 2525 3434 0 net86
rlabel metal2 12834 8262 12834 8262 0 net87
rlabel metal1 7007 14314 7007 14314 0 net88
rlabel metal1 2428 8942 2428 8942 0 net89
rlabel metal1 1656 13906 1656 13906 0 net9
rlabel metal2 10074 9826 10074 9826 0 net90
rlabel metal1 4753 13974 4753 13974 0 net91
rlabel metal1 4232 6426 4232 6426 0 net92
rlabel metal1 5239 3434 5239 3434 0 net93
rlabel via1 3178 10030 3178 10030 0 net94
rlabel metal1 4170 3094 4170 3094 0 net95
rlabel metal1 10483 11118 10483 11118 0 net96
rlabel metal1 7498 14246 7498 14246 0 net97
rlabel via1 2994 8466 2994 8466 0 net98
rlabel via1 7309 12818 7309 12818 0 net99
rlabel metal2 4094 2363 4094 2363 0 prog_clk
rlabel metal1 13524 16558 13524 16558 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 13110 17204 13110 17204 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 16000 20000
<< end >>
