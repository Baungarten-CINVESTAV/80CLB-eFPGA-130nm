magic
tech sky130A
magscale 1 2
timestamp 1707853339
<< viali >>
rect 6653 9673 6687 9707
rect 7941 9673 7975 9707
rect 8585 9673 8619 9707
rect 10425 9673 10459 9707
rect 4353 9605 4387 9639
rect 10149 9605 10183 9639
rect 1685 9537 1719 9571
rect 1777 9537 1811 9571
rect 2145 9537 2179 9571
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 3249 9537 3283 9571
rect 3617 9537 3651 9571
rect 4997 9537 5031 9571
rect 5273 9537 5307 9571
rect 5641 9537 5675 9571
rect 5917 9537 5951 9571
rect 6377 9537 6411 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 7481 9537 7515 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 7849 9537 7883 9571
rect 8769 9537 8803 9571
rect 9505 9537 9539 9571
rect 9781 9537 9815 9571
rect 4445 9469 4479 9503
rect 5825 9469 5859 9503
rect 6193 9469 6227 9503
rect 8125 9469 8159 9503
rect 1501 9401 1535 9435
rect 3893 9401 3927 9435
rect 9597 9401 9631 9435
rect 2421 9333 2455 9367
rect 3433 9333 3467 9367
rect 4813 9333 4847 9367
rect 5089 9333 5123 9367
rect 5549 9333 5583 9367
rect 6561 9333 6595 9367
rect 7021 9333 7055 9367
rect 7297 9333 7331 9367
rect 9321 9333 9355 9367
rect 2237 9129 2271 9163
rect 6101 9129 6135 9163
rect 6837 9129 6871 9163
rect 7205 9129 7239 9163
rect 7481 9061 7515 9095
rect 10425 9061 10459 9095
rect 4997 8993 5031 9027
rect 5917 8993 5951 9027
rect 6469 8993 6503 9027
rect 6653 8993 6687 9027
rect 2697 8925 2731 8959
rect 3065 8925 3099 8959
rect 4629 8925 4663 8959
rect 5733 8925 5767 8959
rect 7389 8925 7423 8959
rect 7665 8925 7699 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 1777 8857 1811 8891
rect 2329 8857 2363 8891
rect 3893 8857 3927 8891
rect 3985 8857 4019 8891
rect 4537 8857 4571 8891
rect 1501 8789 1535 8823
rect 2881 8789 2915 8823
rect 3617 8789 3651 8823
rect 4813 8789 4847 8823
rect 5549 8789 5583 8823
rect 9965 8789 9999 8823
rect 1777 8585 1811 8619
rect 4721 8585 4755 8619
rect 6193 8585 6227 8619
rect 6377 8585 6411 8619
rect 9229 8585 9263 8619
rect 5080 8517 5114 8551
rect 7972 8517 8006 8551
rect 1593 8449 1627 8483
rect 1869 8449 1903 8483
rect 2125 8449 2159 8483
rect 3341 8449 3375 8483
rect 3597 8449 3631 8483
rect 4813 8449 4847 8483
rect 6561 8449 6595 8483
rect 8493 8449 8527 8483
rect 9413 8449 9447 8483
rect 10149 8449 10183 8483
rect 8217 8381 8251 8415
rect 3249 8313 3283 8347
rect 6837 8245 6871 8279
rect 8401 8245 8435 8279
rect 10425 8245 10459 8279
rect 1869 8041 1903 8075
rect 3249 8041 3283 8075
rect 5733 8041 5767 8075
rect 5825 8041 5859 8075
rect 10149 8041 10183 8075
rect 3433 7973 3467 8007
rect 7849 7973 7883 8007
rect 9965 7973 9999 8007
rect 1685 7905 1719 7939
rect 2605 7905 2639 7939
rect 2789 7905 2823 7939
rect 4629 7905 4663 7939
rect 5089 7905 5123 7939
rect 5273 7905 5307 7939
rect 8217 7905 8251 7939
rect 1593 7837 1627 7871
rect 2513 7837 2547 7871
rect 3617 7837 3651 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 7665 7837 7699 7871
rect 8033 7837 8067 7871
rect 10057 7837 10091 7871
rect 10333 7837 10367 7871
rect 3801 7769 3835 7803
rect 4169 7769 4203 7803
rect 4905 7769 4939 7803
rect 6561 7701 6595 7735
rect 7573 7701 7607 7735
rect 8677 7701 8711 7735
rect 8953 7701 8987 7735
rect 2973 7497 3007 7531
rect 6745 7497 6779 7531
rect 7757 7497 7791 7531
rect 8309 7497 8343 7531
rect 2614 7361 2648 7395
rect 2881 7361 2915 7395
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 8953 7361 8987 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 3433 7293 3467 7327
rect 3709 7293 3743 7327
rect 3893 7293 3927 7327
rect 8125 7293 8159 7327
rect 8769 7293 8803 7327
rect 9045 7293 9079 7327
rect 9229 7293 9263 7327
rect 1501 7157 1535 7191
rect 4353 7157 4387 7191
rect 5733 7157 5767 7191
rect 6469 7157 6503 7191
rect 9413 7157 9447 7191
rect 10425 7157 10459 7191
rect 9413 6953 9447 6987
rect 5457 6885 5491 6919
rect 8125 6885 8159 6919
rect 8493 6885 8527 6919
rect 2789 6817 2823 6851
rect 2973 6817 3007 6851
rect 3617 6817 3651 6851
rect 4077 6817 4111 6851
rect 4445 6817 4479 6851
rect 8953 6817 8987 6851
rect 9137 6817 9171 6851
rect 9689 6817 9723 6851
rect 4629 6749 4663 6783
rect 5089 6749 5123 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 8677 6749 8711 6783
rect 9873 6749 9907 6783
rect 2544 6681 2578 6715
rect 3065 6681 3099 6715
rect 4353 6681 4387 6715
rect 6184 6681 6218 6715
rect 1409 6613 1443 6647
rect 4721 6613 4755 6647
rect 4905 6613 4939 6647
rect 7297 6613 7331 6647
rect 8309 6613 8343 6647
rect 10333 6613 10367 6647
rect 2697 6409 2731 6443
rect 2789 6409 2823 6443
rect 4353 6409 4387 6443
rect 5549 6409 5583 6443
rect 10057 6409 10091 6443
rect 10425 6409 10459 6443
rect 1777 6341 1811 6375
rect 7604 6341 7638 6375
rect 8677 6341 8711 6375
rect 1409 6273 1443 6307
rect 4997 6273 5031 6307
rect 7849 6273 7883 6307
rect 9597 6273 9631 6307
rect 10241 6273 10275 6307
rect 2053 6205 2087 6239
rect 3341 6205 3375 6239
rect 4077 6205 4111 6239
rect 4261 6205 4295 6239
rect 4813 6205 4847 6239
rect 5089 6205 5123 6239
rect 6009 6205 6043 6239
rect 6193 6205 6227 6239
rect 8585 6205 8619 6239
rect 9229 6205 9263 6239
rect 9413 6205 9447 6239
rect 3617 6069 3651 6103
rect 6469 6069 6503 6103
rect 7941 6069 7975 6103
rect 3249 5865 3283 5899
rect 3617 5865 3651 5899
rect 5181 5865 5215 5899
rect 8677 5865 8711 5899
rect 4169 5797 4203 5831
rect 8493 5797 8527 5831
rect 4813 5729 4847 5763
rect 6929 5729 6963 5763
rect 7113 5729 7147 5763
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 3893 5661 3927 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 7380 5661 7414 5695
rect 8585 5661 8619 5695
rect 9137 5677 9171 5711
rect 9413 5637 9447 5671
rect 9689 5661 9723 5695
rect 2728 5593 2762 5627
rect 9781 5593 9815 5627
rect 10149 5593 10183 5627
rect 10517 5593 10551 5627
rect 1593 5525 1627 5559
rect 4077 5525 4111 5559
rect 8953 5525 8987 5559
rect 9597 5525 9631 5559
rect 2881 5321 2915 5355
rect 6101 5321 6135 5355
rect 8217 5321 8251 5355
rect 8953 5321 8987 5355
rect 9965 5321 9999 5355
rect 1593 5253 1627 5287
rect 4353 5253 4387 5287
rect 1501 5185 1535 5219
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 2329 5185 2363 5219
rect 4445 5185 4479 5219
rect 5181 5185 5215 5219
rect 5641 5185 5675 5219
rect 5733 5185 5767 5219
rect 6193 5185 6227 5219
rect 7205 5185 7239 5219
rect 9689 5185 9723 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 2421 5117 2455 5151
rect 4629 5117 4663 5151
rect 5273 5117 5307 5151
rect 5825 5117 5859 5151
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 7573 5117 7607 5151
rect 7757 5117 7791 5151
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 4997 5049 5031 5083
rect 9873 5049 9907 5083
rect 5457 4981 5491 5015
rect 6929 4981 6963 5015
rect 7389 4981 7423 5015
rect 10425 4981 10459 5015
rect 1501 4777 1535 4811
rect 2329 4777 2363 4811
rect 3617 4777 3651 4811
rect 3985 4777 4019 4811
rect 4905 4777 4939 4811
rect 5089 4777 5123 4811
rect 5917 4777 5951 4811
rect 7297 4777 7331 4811
rect 8125 4777 8159 4811
rect 3249 4709 3283 4743
rect 5365 4709 5399 4743
rect 8401 4709 8435 4743
rect 1777 4573 1811 4607
rect 2145 4573 2179 4607
rect 2605 4573 2639 4607
rect 2789 4573 2823 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 6193 4573 6227 4607
rect 6653 4573 6687 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 7113 4573 7147 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 8217 4573 8251 4607
rect 6009 4437 6043 4471
rect 1685 4233 1719 4267
rect 3617 4233 3651 4267
rect 5089 4233 5123 4267
rect 5733 4233 5767 4267
rect 1777 4097 1811 4131
rect 1869 4097 1903 4131
rect 2605 4097 2639 4131
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 4077 4097 4111 4131
rect 4445 4097 4479 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 5549 4097 5583 4131
rect 10241 4097 10275 4131
rect 2329 4029 2363 4063
rect 2513 4029 2547 4063
rect 2789 4029 2823 4063
rect 4261 4029 4295 4063
rect 3157 3961 3191 3995
rect 10425 3893 10459 3927
rect 1501 3689 1535 3723
rect 3249 3689 3283 3723
rect 4169 3689 4203 3723
rect 2697 3621 2731 3655
rect 2513 3485 2547 3519
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 10241 3485 10275 3519
rect 1777 3417 1811 3451
rect 1961 3417 1995 3451
rect 2329 3417 2363 3451
rect 3801 3349 3835 3383
rect 10425 3349 10459 3383
rect 1685 3145 1719 3179
rect 2237 3145 2271 3179
rect 2513 3145 2547 3179
rect 2973 3145 3007 3179
rect 3157 3145 3191 3179
rect 3801 3145 3835 3179
rect 10425 3145 10459 3179
rect 1501 3009 1535 3043
rect 1961 3009 1995 3043
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4353 3009 4387 3043
rect 9873 3009 9907 3043
rect 10241 3009 10275 3043
rect 2605 2873 2639 2907
rect 4169 2873 4203 2907
rect 10057 2873 10091 2907
rect 1777 2805 1811 2839
rect 4077 2805 4111 2839
rect 2421 2601 2455 2635
rect 3801 2601 3835 2635
rect 4537 2601 4571 2635
rect 5641 2601 5675 2635
rect 6837 2601 6871 2635
rect 8033 2601 8067 2635
rect 9229 2601 9263 2635
rect 10425 2601 10459 2635
rect 3525 2533 3559 2567
rect 4813 2533 4847 2567
rect 1777 2397 1811 2431
rect 2145 2397 2179 2431
rect 2513 2397 2547 2431
rect 2605 2397 2639 2431
rect 3065 2397 3099 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 5457 2397 5491 2431
rect 6653 2397 6687 2431
rect 7849 2397 7883 2431
rect 9045 2397 9079 2431
rect 9873 2397 9907 2431
rect 10241 2397 10275 2431
rect 1409 2329 1443 2363
rect 2053 2329 2087 2363
rect 2789 2261 2823 2295
rect 3249 2261 3283 2295
rect 4445 2261 4479 2295
rect 10057 2261 10091 2295
<< metal1 >>
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 9858 10112 9864 10124
rect 5776 10084 9864 10112
rect 5776 10072 5782 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 7926 9976 7932 9988
rect 4304 9948 7932 9976
rect 4304 9936 4310 9948
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 6914 9908 6920 9920
rect 4396 9880 6920 9908
rect 4396 9868 4402 9880
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 750 9664 756 9716
rect 808 9704 814 9716
rect 808 9676 2774 9704
rect 808 9664 814 9676
rect 934 9596 940 9648
rect 992 9636 998 9648
rect 2746 9636 2774 9676
rect 4614 9664 4620 9716
rect 4672 9664 4678 9716
rect 6178 9664 6184 9716
rect 6236 9664 6242 9716
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 6328 9676 6653 9704
rect 6328 9664 6334 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 7926 9664 7932 9716
rect 7984 9664 7990 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8573 9707 8631 9713
rect 8573 9704 8585 9707
rect 8076 9676 8585 9704
rect 8076 9664 8082 9676
rect 8573 9673 8585 9676
rect 8619 9673 8631 9707
rect 8573 9667 8631 9673
rect 8662 9664 8668 9716
rect 8720 9664 8726 9716
rect 9766 9664 9772 9716
rect 9824 9664 9830 9716
rect 10413 9707 10471 9713
rect 10413 9673 10425 9707
rect 10459 9704 10471 9707
rect 10502 9704 10508 9716
rect 10459 9676 10508 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 992 9608 1808 9636
rect 2746 9608 3648 9636
rect 992 9596 998 9608
rect 1780 9577 1808 9608
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1596 9540 1685 9568
rect 1394 9392 1400 9444
rect 1452 9432 1458 9444
rect 1489 9435 1547 9441
rect 1489 9432 1501 9435
rect 1452 9404 1501 9432
rect 1452 9392 1458 9404
rect 1489 9401 1501 9404
rect 1535 9401 1547 9435
rect 1596 9432 1624 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2130 9528 2136 9580
rect 2188 9528 2194 9580
rect 2682 9528 2688 9580
rect 2740 9528 2746 9580
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3510 9568 3516 9580
rect 3283 9540 3516 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3620 9577 3648 9608
rect 4338 9596 4344 9648
rect 4396 9596 4402 9648
rect 4632 9636 4660 9664
rect 4632 9608 5304 9636
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5276 9577 5304 9608
rect 5350 9596 5356 9648
rect 5408 9636 5414 9648
rect 6196 9636 6224 9664
rect 5408 9608 6040 9636
rect 6196 9608 6868 9636
rect 5408 9596 5414 9608
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 6012 9568 6040 9608
rect 6012 9540 6316 9568
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 3234 9432 3240 9444
rect 1596 9404 3240 9432
rect 1489 9395 1547 9401
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 3881 9435 3939 9441
rect 3881 9401 3893 9435
rect 3927 9401 3939 9435
rect 4448 9432 4476 9463
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 4672 9472 5825 9500
rect 4672 9460 4678 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 6178 9460 6184 9512
rect 6236 9460 6242 9512
rect 6288 9500 6316 9540
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6840 9577 6868 9608
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 7208 9568 7236 9664
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7208 9540 7481 9568
rect 6917 9531 6975 9537
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 6932 9500 6960 9531
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 7834 9528 7840 9580
rect 7892 9528 7898 9580
rect 8680 9568 8708 9664
rect 9784 9636 9812 9664
rect 9508 9608 9812 9636
rect 9508 9577 9536 9608
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 9916 9608 10149 9636
rect 9916 9596 9922 9608
rect 10137 9605 10149 9608
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8680 9540 8769 9568
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 6288 9472 6960 9500
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 9784 9500 9812 9531
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10520 9500 10548 9528
rect 9784 9472 10548 9500
rect 8113 9463 8171 9469
rect 8128 9432 8156 9463
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 4448 9404 8156 9432
rect 8220 9404 9597 9432
rect 3881 9395 3939 9401
rect 1210 9324 1216 9376
rect 1268 9364 1274 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 1268 9336 2421 9364
rect 1268 9324 1274 9336
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 2648 9336 3433 9364
rect 2648 9324 2654 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3896 9364 3924 9395
rect 4338 9364 4344 9376
rect 3896 9336 4344 9364
rect 3421 9327 3479 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4580 9336 4813 9364
rect 4580 9324 4586 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 5074 9324 5080 9376
rect 5132 9324 5138 9376
rect 5534 9324 5540 9376
rect 5592 9324 5598 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6788 9336 7021 9364
rect 6788 9324 6794 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7374 9364 7380 9376
rect 7331 9336 7380 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8220 9364 8248 9404
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 8168 9336 8248 9364
rect 8168 9324 8174 9336
rect 9306 9324 9312 9376
rect 9364 9324 9370 9376
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2774 9160 2780 9172
rect 2271 9132 2780 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 4430 9160 4436 9172
rect 3568 9132 4436 9160
rect 3568 9120 3574 9132
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5960 9132 6101 9160
rect 5960 9120 5966 9132
rect 6089 9129 6101 9132
rect 6135 9160 6147 9163
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6135 9132 6837 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 6825 9123 6883 9129
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6972 9132 7205 9160
rect 6972 9120 6978 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 2682 9052 2688 9104
rect 2740 9052 2746 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 4126 9064 7481 9092
rect 2700 9024 2728 9052
rect 4126 9024 4154 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 7469 9055 7527 9061
rect 10410 9052 10416 9104
rect 10468 9052 10474 9104
rect 11054 9052 11060 9104
rect 11112 9052 11118 9104
rect 2700 8996 4154 9024
rect 4522 8984 4528 9036
rect 4580 8984 4586 9036
rect 4982 8984 4988 9036
rect 5040 8984 5046 9036
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5592 8996 5917 9024
rect 5592 8984 5598 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6236 8996 6469 9024
rect 6236 8984 6242 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 6604 8996 6653 9024
rect 6604 8984 6610 8996
rect 6641 8993 6653 8996
rect 6687 8993 6699 9027
rect 11072 9024 11100 9052
rect 6641 8987 6699 8993
rect 10152 8996 11100 9024
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2096 8928 2697 8956
rect 2096 8916 2102 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3694 8956 3700 8968
rect 3108 8928 3700 8956
rect 3108 8916 3114 8928
rect 3694 8916 3700 8928
rect 3752 8916 3758 8968
rect 4540 8956 4568 8984
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4540 8928 4629 8956
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 5368 8956 5396 8984
rect 4617 8919 4675 8925
rect 4816 8928 5396 8956
rect 1762 8848 1768 8900
rect 1820 8848 1826 8900
rect 2317 8891 2375 8897
rect 2317 8857 2329 8891
rect 2363 8888 2375 8891
rect 2406 8888 2412 8900
rect 2363 8860 2412 8888
rect 2363 8857 2375 8860
rect 2317 8851 2375 8857
rect 2406 8848 2412 8860
rect 2464 8848 2470 8900
rect 3878 8848 3884 8900
rect 3936 8848 3942 8900
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8857 4031 8891
rect 3973 8851 4031 8857
rect 1486 8780 1492 8832
rect 1544 8780 1550 8832
rect 2866 8780 2872 8832
rect 2924 8780 2930 8832
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3605 8823 3663 8829
rect 3605 8820 3617 8823
rect 3292 8792 3617 8820
rect 3292 8780 3298 8792
rect 3605 8789 3617 8792
rect 3651 8789 3663 8823
rect 3988 8820 4016 8851
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 4396 8860 4537 8888
rect 4396 8848 4402 8860
rect 4525 8857 4537 8860
rect 4571 8888 4583 8891
rect 4816 8888 4844 8928
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 10152 8965 10180 8996
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6886 8928 7389 8956
rect 4571 8860 4844 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 6886 8888 6914 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 10137 8959 10195 8965
rect 7699 8928 8708 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 4948 8860 6914 8888
rect 4948 8848 4954 8860
rect 8680 8832 8708 8928
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 4246 8820 4252 8832
rect 3988 8792 4252 8820
rect 3605 8783 3663 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 5166 8820 5172 8832
rect 4847 8792 5172 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 8720 8792 9965 8820
rect 8720 8780 8726 8792
rect 9953 8789 9965 8792
rect 9999 8789 10011 8823
rect 9953 8783 10011 8789
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 4709 8619 4767 8625
rect 1811 8588 4660 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2866 8548 2872 8560
rect 1872 8520 2872 8548
rect 1872 8489 1900 8520
rect 2866 8508 2872 8520
rect 2924 8548 2930 8560
rect 4632 8548 4660 8588
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 4982 8616 4988 8628
rect 4755 8588 4988 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 5684 8588 6193 8616
rect 5684 8576 5690 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6181 8579 6239 8585
rect 4890 8548 4896 8560
rect 2924 8520 4154 8548
rect 4632 8520 4896 8548
rect 2924 8508 2930 8520
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 1596 8412 1624 8443
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2113 8483 2171 8489
rect 2113 8480 2125 8483
rect 2004 8452 2125 8480
rect 2004 8440 2010 8452
rect 2113 8449 2125 8452
rect 2159 8449 2171 8483
rect 2113 8443 2171 8449
rect 3050 8440 3056 8492
rect 3108 8440 3114 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3344 8489 3372 8520
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3585 8483 3643 8489
rect 3585 8480 3597 8483
rect 3329 8443 3387 8449
rect 3436 8452 3597 8480
rect 1596 8384 1900 8412
rect 1872 8276 1900 8384
rect 3068 8344 3096 8440
rect 3252 8412 3280 8440
rect 3436 8412 3464 8452
rect 3585 8449 3597 8452
rect 3631 8449 3643 8483
rect 4126 8480 4154 8520
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 5068 8551 5126 8557
rect 5068 8517 5080 8551
rect 5114 8548 5126 8551
rect 5534 8548 5540 8560
rect 5114 8520 5540 8548
rect 5114 8517 5126 8520
rect 5068 8511 5126 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4126 8452 4813 8480
rect 3585 8443 3643 8449
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 6196 8480 6224 8579
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 8662 8576 8668 8628
rect 8720 8576 8726 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 9306 8576 9312 8628
rect 9364 8576 9370 8628
rect 7960 8551 8018 8557
rect 7960 8517 7972 8551
rect 8006 8548 8018 8551
rect 8110 8548 8116 8560
rect 8006 8520 8116 8548
rect 8006 8517 8018 8520
rect 7960 8511 8018 8517
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6196 8452 6561 8480
rect 4801 8443 4859 8449
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8680 8480 8708 8576
rect 8527 8452 8708 8480
rect 9324 8480 9352 8576
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9324 8452 9413 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 3252 8384 3464 8412
rect 8202 8372 8208 8424
rect 8260 8372 8266 8424
rect 3237 8347 3295 8353
rect 3237 8344 3249 8347
rect 2792 8316 3249 8344
rect 2792 8276 2820 8316
rect 3237 8313 3249 8316
rect 3283 8313 3295 8347
rect 3237 8307 3295 8313
rect 1872 8248 2820 8276
rect 6822 8236 6828 8288
rect 6880 8236 6886 8288
rect 8386 8236 8392 8288
rect 8444 8236 8450 8288
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 10502 8276 10508 8288
rect 10459 8248 10508 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 1857 8075 1915 8081
rect 1857 8041 1869 8075
rect 1903 8072 1915 8075
rect 1946 8072 1952 8084
rect 1903 8044 1952 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3878 8072 3884 8084
rect 3292 8044 3884 8072
rect 3292 8032 3298 8044
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 5074 8072 5080 8084
rect 4540 8044 5080 8072
rect 3421 8007 3479 8013
rect 3421 8004 3433 8007
rect 2792 7976 3433 8004
rect 2792 7945 2820 7976
rect 3421 7973 3433 7976
rect 3467 7973 3479 8007
rect 3421 7967 3479 7973
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2593 7939 2651 7945
rect 2593 7936 2605 7939
rect 1719 7908 2605 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2593 7905 2605 7908
rect 2639 7905 2651 7939
rect 2593 7899 2651 7905
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1452 7840 1593 7868
rect 1452 7828 1458 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2038 7868 2044 7880
rect 1627 7840 2044 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2498 7828 2504 7880
rect 2556 7828 2562 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 3970 7868 3976 7880
rect 3651 7840 3976 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4540 7877 4568 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5776 8044 5825 8072
rect 5776 8032 5782 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 10226 8032 10232 8084
rect 10284 8032 10290 8084
rect 7650 7964 7656 8016
rect 7708 7964 7714 8016
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 10244 8004 10272 8032
rect 9999 7976 10272 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4663 7908 5089 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 5224 7908 5273 7936
rect 5224 7896 5230 7908
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 7668 7936 7696 7964
rect 5261 7899 5319 7905
rect 7392 7908 7696 7936
rect 7852 7936 7880 7967
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 7852 7908 8217 7936
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4264 7840 4537 7868
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 3789 7803 3847 7809
rect 3789 7800 3801 7803
rect 1360 7772 3801 7800
rect 1360 7760 1366 7772
rect 3789 7769 3801 7772
rect 3835 7769 3847 7803
rect 3789 7763 3847 7769
rect 4154 7760 4160 7812
rect 4212 7760 4218 7812
rect 4264 7744 4292 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4982 7868 4988 7880
rect 4847 7840 4988 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 6288 7800 6316 7831
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7392 7877 7420 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6880 7840 7205 7868
rect 6880 7828 6886 7840
rect 7193 7837 7205 7840
rect 7239 7868 7251 7871
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7239 7840 7389 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7377 7831 7435 7837
rect 7576 7840 7665 7868
rect 4939 7772 6316 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 7576 7741 7604 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8404 7868 8432 7896
rect 8067 7840 8432 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10336 7744 10364 7831
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 8662 7692 8668 7744
rect 8720 7692 8726 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2590 7528 2596 7540
rect 2004 7500 2596 7528
rect 2004 7488 2010 7500
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3234 7528 3240 7540
rect 3007 7500 3240 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 4154 7488 4160 7540
rect 4212 7488 4218 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6512 7500 6745 7528
rect 6512 7488 6518 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 6733 7491 6791 7497
rect 6886 7500 7757 7528
rect 4172 7460 4200 7488
rect 6886 7460 6914 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8662 7528 8668 7540
rect 8343 7500 8668 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 8036 7460 8064 7488
rect 4172 7432 6914 7460
rect 7944 7432 8064 7460
rect 2590 7352 2596 7404
rect 2648 7401 2654 7404
rect 2648 7355 2660 7401
rect 2648 7352 2654 7355
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 4062 7392 4068 7404
rect 3651 7364 4068 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3016 7296 3433 7324
rect 3016 7284 3022 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3786 7324 3792 7336
rect 3743 7296 3792 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 3878 7284 3884 7336
rect 3936 7284 3942 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6564 7324 6592 7355
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 7944 7401 7972 7432
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8680 7392 8708 7488
rect 8941 7395 8999 7401
rect 8680 7364 8892 7392
rect 8021 7355 8079 7361
rect 7374 7324 7380 7336
rect 5592 7296 7380 7324
rect 5592 7284 5598 7296
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 8036 7324 8064 7355
rect 7708 7296 8064 7324
rect 8113 7327 8171 7333
rect 7708 7284 7714 7296
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8159 7296 8769 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8864 7324 8892 7364
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 8987 7364 9873 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8864 7296 9045 7324
rect 8757 7287 8815 7293
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9968 7324 9996 7355
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 10318 7324 10324 7336
rect 9968 7296 10324 7324
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 2498 7188 2504 7200
rect 1535 7160 2504 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 5718 7148 5724 7200
rect 5776 7148 5782 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5868 7160 6469 7188
rect 5868 7148 5874 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 9398 7148 9404 7200
rect 9456 7148 9462 7200
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 2866 6944 2872 6996
rect 2924 6944 2930 6996
rect 7558 6984 7564 6996
rect 4172 6956 7564 6984
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 2884 6848 2912 6944
rect 2823 6820 2912 6848
rect 2961 6851 3019 6857
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3142 6848 3148 6860
rect 3007 6820 3148 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3605 6851 3663 6857
rect 3605 6817 3617 6851
rect 3651 6848 3663 6851
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3651 6820 4077 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 4065 6817 4077 6820
rect 4111 6848 4123 6851
rect 4172 6848 4200 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 9398 6984 9404 6996
rect 8128 6956 9168 6984
rect 9359 6956 9404 6984
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 4396 6888 4476 6916
rect 4396 6876 4402 6888
rect 4448 6857 4476 6888
rect 5442 6876 5448 6928
rect 5500 6876 5506 6928
rect 8128 6925 8156 6956
rect 8113 6919 8171 6925
rect 8113 6885 8125 6919
rect 8159 6885 8171 6919
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 8113 6879 8171 6885
rect 8266 6888 8493 6916
rect 4111 6820 4200 6848
rect 4433 6851 4491 6857
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 8266 6848 8294 6888
rect 8481 6885 8493 6888
rect 8527 6885 8539 6919
rect 8481 6879 8539 6885
rect 8846 6848 8852 6860
rect 4433 6811 4491 6817
rect 7944 6820 8294 6848
rect 8404 6820 8852 6848
rect 4614 6740 4620 6792
rect 4672 6740 4678 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5534 6780 5540 6792
rect 5123 6752 5540 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 7944 6789 7972 6820
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 7929 6783 7987 6789
rect 5951 6752 6914 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6886 6724 6914 6752
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8404 6780 8432 6820
rect 8680 6789 8708 6820
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 9140 6857 9168 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6817 9183 6851
rect 9416 6848 9444 6944
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9416 6820 9689 6848
rect 9125 6811 9183 6817
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 8251 6752 8432 6780
rect 8665 6783 8723 6789
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8665 6749 8677 6783
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 2532 6715 2590 6721
rect 2532 6681 2544 6715
rect 2578 6712 2590 6715
rect 2774 6712 2780 6724
rect 2578 6684 2780 6712
rect 2578 6681 2590 6684
rect 2532 6675 2590 6681
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 3050 6672 3056 6724
rect 3108 6672 3114 6724
rect 4062 6672 4068 6724
rect 4120 6672 4126 6724
rect 4341 6715 4399 6721
rect 4341 6681 4353 6715
rect 4387 6712 4399 6715
rect 4430 6712 4436 6724
rect 4387 6684 4436 6712
rect 4387 6681 4399 6684
rect 4341 6675 4399 6681
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 6172 6715 6230 6721
rect 6172 6681 6184 6715
rect 6218 6712 6230 6715
rect 6546 6712 6552 6724
rect 6218 6684 6552 6712
rect 6218 6681 6230 6684
rect 6172 6675 6230 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 6886 6684 6920 6724
rect 6914 6672 6920 6684
rect 6972 6712 6978 6724
rect 8128 6712 8156 6740
rect 6972 6684 8156 6712
rect 6972 6672 6978 6684
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 1670 6644 1676 6656
rect 1443 6616 1676 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 4080 6644 4108 6672
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4080 6616 4721 6644
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4890 6604 4896 6656
rect 4948 6604 4954 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 8220 6644 8248 6743
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 7331 6616 8248 6644
rect 8297 6647 8355 6653
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 9214 6644 9220 6656
rect 8343 6616 9220 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 10042 6604 10048 6656
rect 10100 6644 10106 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10100 6616 10333 6644
rect 10100 6604 10106 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2648 6412 2697 6440
rect 2648 6400 2654 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 4338 6400 4344 6452
rect 4396 6400 4402 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 5500 6412 5549 6440
rect 5500 6400 5506 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 10042 6400 10048 6452
rect 10100 6400 10106 6452
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 1765 6375 1823 6381
rect 1765 6341 1777 6375
rect 1811 6372 1823 6375
rect 4890 6372 4896 6384
rect 1811 6344 4896 6372
rect 1811 6341 1823 6344
rect 1765 6335 1823 6341
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4985 6307 5043 6313
rect 3844 6276 4936 6304
rect 3844 6264 3850 6276
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1728 6208 2053 6236
rect 1728 6196 1734 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 3326 6196 3332 6248
rect 3384 6196 3390 6248
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 4028 6208 4077 6236
rect 4028 6196 4034 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4246 6196 4252 6248
rect 4304 6196 4310 6248
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4908 6236 4936 6276
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5460 6304 5488 6400
rect 7592 6375 7650 6381
rect 7592 6341 7604 6375
rect 7638 6372 7650 6375
rect 8665 6375 8723 6381
rect 8665 6372 8677 6375
rect 7638 6344 8677 6372
rect 7638 6341 7650 6344
rect 7592 6335 7650 6341
rect 8665 6341 8677 6344
rect 8711 6341 8723 6375
rect 8665 6335 8723 6341
rect 5031 6276 5488 6304
rect 7837 6307 7895 6313
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8110 6304 8116 6316
rect 7883 6276 8116 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9180 6276 9597 6304
rect 9180 6264 9186 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10192 6276 10241 6304
rect 10192 6264 10198 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4908 6208 5089 6236
rect 4801 6199 4859 6205
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 4816 6168 4844 6199
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5592 6208 6009 6236
rect 5592 6196 5598 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6178 6196 6184 6248
rect 6236 6196 6242 6248
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8846 6236 8852 6248
rect 8619 6208 8852 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 8996 6208 9229 6236
rect 8996 6196 9002 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 3292 6140 4844 6168
rect 3292 6128 3298 6140
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3200 6072 3617 6100
rect 3200 6060 3206 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 6454 6060 6460 6112
rect 6512 6060 6518 6112
rect 7926 6060 7932 6112
rect 7984 6060 7990 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3878 5896 3884 5908
rect 3651 5868 3884 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5626 5896 5632 5908
rect 5215 5868 5632 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 9122 5896 9128 5908
rect 8711 5868 9128 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 4157 5831 4215 5837
rect 4157 5828 4169 5831
rect 3068 5800 4169 5828
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2924 5664 2973 5692
rect 2924 5652 2930 5664
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 2716 5627 2774 5633
rect 2716 5593 2728 5627
rect 2762 5624 2774 5627
rect 3068 5624 3096 5800
rect 4157 5797 4169 5800
rect 4203 5797 4215 5831
rect 4157 5791 4215 5797
rect 8481 5831 8539 5837
rect 8481 5797 8493 5831
rect 8527 5828 8539 5831
rect 8527 5800 8616 5828
rect 8527 5797 8539 5800
rect 8481 5791 8539 5797
rect 3326 5760 3332 5772
rect 3160 5732 3332 5760
rect 3160 5701 3188 5732
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 3896 5732 4813 5760
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3786 5692 3792 5704
rect 3467 5664 3792 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 2762 5596 3096 5624
rect 2762 5593 2774 5596
rect 2716 5587 2774 5593
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1544 5528 1593 5556
rect 1544 5516 1550 5528
rect 1581 5525 1593 5528
rect 1627 5556 1639 5559
rect 3160 5556 3188 5655
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 3896 5701 3924 5732
rect 4801 5729 4813 5732
rect 4847 5760 4859 5763
rect 5166 5760 5172 5772
rect 4847 5732 5172 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5166 5720 5172 5732
rect 5224 5760 5230 5772
rect 6454 5760 6460 5772
rect 5224 5732 6460 5760
rect 5224 5720 5230 5732
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 6972 5732 7113 5760
rect 6972 5720 6978 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7101 5723 7159 5729
rect 8588 5760 8616 5800
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 9214 5828 9220 5840
rect 8904 5800 9220 5828
rect 8904 5788 8910 5800
rect 9214 5788 9220 5800
rect 9272 5828 9278 5840
rect 9272 5800 9720 5828
rect 9272 5788 9278 5800
rect 8938 5760 8944 5772
rect 8588 5732 8944 5760
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5000 5624 5028 5655
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5718 5692 5724 5704
rect 5316 5664 5724 5692
rect 5316 5652 5322 5664
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 7368 5695 7426 5701
rect 7368 5661 7380 5695
rect 7414 5692 7426 5695
rect 7926 5692 7932 5704
rect 7414 5664 7932 5692
rect 7414 5661 7426 5664
rect 7368 5655 7426 5661
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8588 5701 8616 5732
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 4080 5596 5028 5624
rect 8956 5624 8984 5720
rect 9125 5711 9183 5717
rect 9125 5677 9137 5711
rect 9171 5708 9183 5711
rect 9171 5704 9260 5708
rect 9171 5680 9220 5704
rect 9171 5677 9183 5680
rect 9125 5671 9183 5677
rect 9214 5652 9220 5680
rect 9272 5652 9278 5704
rect 9692 5701 9720 5800
rect 9677 5695 9735 5701
rect 9401 5671 9459 5677
rect 9401 5668 9413 5671
rect 9324 5640 9413 5668
rect 8956 5596 9076 5624
rect 3234 5556 3240 5568
rect 1627 5528 3240 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 4080 5565 4108 5596
rect 4065 5559 4123 5565
rect 4065 5525 4077 5559
rect 4111 5525 4123 5559
rect 4065 5519 4123 5525
rect 8938 5516 8944 5568
rect 8996 5516 9002 5568
rect 9048 5556 9076 5596
rect 9324 5556 9352 5640
rect 9401 5637 9413 5640
rect 9447 5637 9459 5671
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 9401 5631 9459 5637
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9548 5596 9781 5624
rect 9548 5584 9554 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 9950 5584 9956 5636
rect 10008 5624 10014 5636
rect 10137 5627 10195 5633
rect 10137 5624 10149 5627
rect 10008 5596 10149 5624
rect 10008 5584 10014 5596
rect 10137 5593 10149 5596
rect 10183 5593 10195 5627
rect 10137 5587 10195 5593
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 9048 5528 9352 5556
rect 9582 5516 9588 5568
rect 9640 5516 9646 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 2498 5312 2504 5364
rect 2556 5312 2562 5364
rect 2866 5312 2872 5364
rect 2924 5312 2930 5364
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 4062 5352 4068 5364
rect 3384 5324 4068 5352
rect 3384 5312 3390 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 6089 5355 6147 5361
rect 6089 5321 6101 5355
rect 6135 5352 6147 5355
rect 6178 5352 6184 5364
rect 6135 5324 6184 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6270 5312 6276 5364
rect 6328 5312 6334 5364
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8251 5324 8953 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 8941 5321 8953 5324
rect 8987 5352 8999 5355
rect 9398 5352 9404 5364
rect 8987 5324 9404 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9490 5312 9496 5364
rect 9548 5312 9554 5364
rect 9582 5312 9588 5364
rect 9640 5312 9646 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9916 5324 9965 5352
rect 9916 5312 9922 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 10226 5312 10232 5364
rect 10284 5312 10290 5364
rect 1581 5287 1639 5293
rect 1581 5253 1593 5287
rect 1627 5284 1639 5287
rect 1627 5256 2268 5284
rect 1627 5253 1639 5256
rect 1581 5247 1639 5253
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 1670 5216 1676 5228
rect 1535 5188 1676 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1780 5148 1808 5179
rect 992 5120 1808 5148
rect 992 5108 998 5120
rect 2148 5012 2176 5179
rect 2240 5080 2268 5256
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2516 5216 2544 5312
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 5258 5284 5264 5296
rect 4387 5256 5264 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 6288 5284 6316 5312
rect 9508 5284 9536 5312
rect 5736 5256 6316 5284
rect 7760 5256 9536 5284
rect 9600 5284 9628 5312
rect 10244 5284 10272 5312
rect 9600 5256 10180 5284
rect 10244 5256 10364 5284
rect 2363 5188 2544 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 2740 5188 4445 5216
rect 2740 5176 2746 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 5736 5225 5764 5256
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5675 5188 5733 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6822 5216 6828 5228
rect 6227 5188 6828 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6822 5176 6828 5188
rect 6880 5216 6886 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6880 5188 7205 5216
rect 6880 5176 6886 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2958 5148 2964 5160
rect 2455 5120 2964 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5074 5148 5080 5160
rect 4663 5120 5080 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5534 5148 5540 5160
rect 5307 5120 5540 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 5859 5120 6469 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 7760 5157 7788 5256
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 10152 5225 10180 5256
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9272 5188 9689 5216
rect 9272 5176 9278 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 6604 5120 6653 5148
rect 6604 5108 6610 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 6641 5111 6699 5117
rect 6748 5120 7573 5148
rect 3050 5080 3056 5092
rect 2240 5052 3056 5080
rect 3050 5040 3056 5052
rect 3108 5040 3114 5092
rect 4982 5040 4988 5092
rect 5040 5080 5046 5092
rect 6748 5080 6776 5120
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 8312 5080 8340 5111
rect 8478 5108 8484 5160
rect 8536 5108 8542 5160
rect 5040 5052 6776 5080
rect 6932 5052 8340 5080
rect 9861 5083 9919 5089
rect 5040 5040 5046 5052
rect 6932 5024 6960 5052
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 10336 5080 10364 5256
rect 9907 5052 10364 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 4062 5012 4068 5024
rect 2148 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5442 4972 5448 5024
rect 5500 4972 5506 5024
rect 6914 4972 6920 5024
rect 6972 4972 6978 5024
rect 7377 5015 7435 5021
rect 7377 4981 7389 5015
rect 7423 5012 7435 5015
rect 9950 5012 9956 5024
rect 7423 4984 9956 5012
rect 7423 4981 7435 4984
rect 7377 4975 7435 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1026 4768 1032 4820
rect 1084 4808 1090 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1084 4780 1501 4808
rect 1084 4768 1090 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 3326 4808 3332 4820
rect 2363 4780 3332 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3786 4808 3792 4820
rect 3651 4780 3792 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 3973 4811 4031 4817
rect 3973 4777 3985 4811
rect 4019 4808 4031 4811
rect 4430 4808 4436 4820
rect 4019 4780 4436 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 4982 4808 4988 4820
rect 4939 4780 4988 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5074 4768 5080 4820
rect 5132 4768 5138 4820
rect 5442 4808 5448 4820
rect 5184 4780 5448 4808
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 3878 4740 3884 4752
rect 3283 4712 3884 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 3878 4700 3884 4712
rect 3936 4740 3942 4752
rect 4246 4740 4252 4752
rect 3936 4712 4252 4740
rect 3936 4700 3942 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 5184 4672 5212 4780
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4808 5963 4811
rect 6546 4808 6552 4820
rect 5951 4780 6552 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6972 4780 7297 4808
rect 6972 4768 6978 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 7650 4768 7656 4820
rect 7708 4768 7714 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8478 4808 8484 4820
rect 8159 4780 8484 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 10226 4768 10232 4820
rect 10284 4768 10290 4820
rect 5353 4743 5411 4749
rect 5353 4709 5365 4743
rect 5399 4709 5411 4743
rect 5353 4703 5411 4709
rect 1780 4644 5212 4672
rect 1780 4613 1808 4644
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2498 4604 2504 4616
rect 2179 4576 2504 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2682 4604 2688 4616
rect 2639 4576 2688 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3234 4604 3240 4616
rect 2823 4576 3240 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3384 4576 3433 4604
rect 3384 4564 3390 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5368 4604 5396 4703
rect 7668 4672 7696 4768
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 10244 4740 10272 4768
rect 8435 4712 10272 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 8938 4672 8944 4684
rect 5552 4644 7880 4672
rect 5552 4613 5580 4644
rect 6196 4613 6224 4644
rect 7852 4613 7880 4644
rect 7944 4644 8944 4672
rect 7944 4613 7972 4644
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5307 4576 5396 4604
rect 5460 4576 5549 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 3344 4536 3372 4564
rect 5460 4548 5488 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6181 4607 6239 4613
rect 5767 4576 6040 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 3108 4508 3372 4536
rect 3108 4496 3114 4508
rect 5442 4496 5448 4548
rect 5500 4496 5506 4548
rect 6012 4477 6040 4576
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 6917 4607 6975 4613
rect 6917 4604 6929 4607
rect 6779 4576 6929 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6917 4573 6929 4576
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7147 4576 7757 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 6546 4496 6552 4548
rect 6604 4536 6610 4548
rect 6656 4536 6684 4567
rect 8220 4536 8248 4567
rect 6604 4508 8248 4536
rect 6604 4496 6610 4508
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4437 6055 4471
rect 5997 4431 6055 4437
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 2682 4264 2688 4276
rect 1719 4236 2688 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 3050 4224 3056 4276
rect 3108 4224 3114 4276
rect 3605 4267 3663 4273
rect 3605 4233 3617 4267
rect 3651 4264 3663 4267
rect 3878 4264 3884 4276
rect 3651 4236 3884 4264
rect 3651 4233 3663 4236
rect 3605 4227 3663 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4488 4236 5089 4264
rect 4488 4224 4494 4236
rect 5077 4233 5089 4236
rect 5123 4233 5135 4267
rect 5077 4227 5135 4233
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 1946 4196 1952 4208
rect 1780 4168 1952 4196
rect 1780 4137 1808 4168
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 3068 4196 3096 4224
rect 5184 4196 5212 4224
rect 3068 4168 3372 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 1903 4100 2605 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2593 4097 2605 4100
rect 2639 4128 2651 4131
rect 3234 4128 3240 4140
rect 2639 4100 3240 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3344 4137 3372 4168
rect 4540 4168 5212 4196
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3970 4128 3976 4140
rect 3467 4100 3976 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4540 4137 4568 4168
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4111 4100 4445 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 5169 4131 5227 4137
rect 4571 4100 4605 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5442 4128 5448 4140
rect 5215 4100 5448 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5534 4088 5540 4140
rect 5592 4088 5598 4140
rect 5736 4128 5764 4227
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 5736 4100 10241 4128
rect 10229 4097 10241 4100
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2363 4032 2452 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2424 3924 2452 4032
rect 2498 4020 2504 4072
rect 2556 4020 2562 4072
rect 2774 4020 2780 4072
rect 2832 4020 2838 4072
rect 4246 4020 4252 4072
rect 4304 4020 4310 4072
rect 5552 4060 5580 4088
rect 6730 4060 6736 4072
rect 5552 4032 6736 4060
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 3142 3952 3148 4004
rect 3200 3952 3206 4004
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 4522 3992 4528 4004
rect 4028 3964 4528 3992
rect 4028 3952 4034 3964
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 2590 3924 2596 3936
rect 2424 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 10410 3884 10416 3936
rect 10468 3884 10474 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 934 3680 940 3732
rect 992 3720 998 3732
rect 1489 3723 1547 3729
rect 1489 3720 1501 3723
rect 992 3692 1501 3720
rect 992 3680 998 3692
rect 1489 3689 1501 3692
rect 1535 3689 1547 3723
rect 1489 3683 1547 3689
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 3786 3680 3792 3732
rect 3844 3680 3850 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 4246 3720 4252 3732
rect 4203 3692 4252 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 2685 3655 2743 3661
rect 2685 3621 2697 3655
rect 2731 3652 2743 3655
rect 3804 3652 3832 3680
rect 2731 3624 3832 3652
rect 2731 3621 2743 3624
rect 2685 3615 2743 3621
rect 4430 3584 4436 3596
rect 1596 3556 4436 3584
rect 1596 3448 1624 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 1728 3488 2513 3516
rect 1728 3476 1734 3488
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2866 3476 2872 3528
rect 2924 3476 2930 3528
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3344 3488 3985 3516
rect 1765 3451 1823 3457
rect 1765 3448 1777 3451
rect 1596 3420 1777 3448
rect 1765 3417 1777 3420
rect 1811 3417 1823 3451
rect 1765 3411 1823 3417
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3417 2007 3451
rect 1949 3411 2007 3417
rect 2317 3451 2375 3457
rect 2317 3417 2329 3451
rect 2363 3448 2375 3451
rect 3142 3448 3148 3460
rect 2363 3420 3148 3448
rect 2363 3417 2375 3420
rect 2317 3411 2375 3417
rect 1026 3340 1032 3392
rect 1084 3380 1090 3392
rect 1964 3380 1992 3411
rect 3142 3408 3148 3420
rect 3200 3408 3206 3460
rect 1084 3352 1992 3380
rect 1084 3340 1090 3352
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 3344 3380 3372 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 3418 3408 3424 3460
rect 3476 3408 3482 3460
rect 4080 3448 4108 3479
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 3896 3420 4108 3448
rect 2280 3352 3372 3380
rect 3436 3380 3464 3408
rect 3896 3392 3924 3420
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3436 3352 3801 3380
rect 2280 3340 2286 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 10410 3340 10416 3392
rect 10468 3340 10474 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3145 1731 3179
rect 1673 3139 1731 3145
rect 1688 3108 1716 3139
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2774 3176 2780 3188
rect 2547 3148 2780 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2924 3148 2973 3176
rect 2924 3136 2930 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3142 3136 3148 3188
rect 3200 3136 3206 3188
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 10226 3176 10232 3188
rect 3835 3148 10232 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10376 3148 10425 3176
rect 10376 3136 10382 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 1688 3080 2360 3108
rect 1486 3000 1492 3052
rect 1544 3000 1550 3052
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2332 3049 2360 3080
rect 2590 3068 2596 3120
rect 2648 3068 2654 3120
rect 4522 3108 4528 3120
rect 2792 3080 4528 3108
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2056 2972 2084 3003
rect 1964 2944 2084 2972
rect 1964 2916 1992 2944
rect 1946 2864 1952 2916
rect 2004 2864 2010 2916
rect 2608 2913 2636 3068
rect 2792 3049 2820 3080
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 1762 2796 1768 2848
rect 1820 2796 1826 2848
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3068 2836 3096 3003
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3292 3012 3341 3040
rect 3292 3000 3298 3012
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3620 2904 3648 3003
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 8076 3012 9873 3040
rect 8076 3000 8082 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10226 3000 10232 3052
rect 10284 3000 10290 3052
rect 3970 2932 3976 2984
rect 4028 2932 4034 2984
rect 4080 2972 4108 3000
rect 4080 2944 4200 2972
rect 3988 2904 4016 2932
rect 4172 2913 4200 2944
rect 10134 2932 10140 2984
rect 10192 2932 10198 2984
rect 3620 2876 4016 2904
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2904 10103 2907
rect 10152 2904 10180 2932
rect 10091 2876 10180 2904
rect 10091 2873 10103 2876
rect 10045 2867 10103 2873
rect 3694 2836 3700 2848
rect 2924 2808 3700 2836
rect 2924 2796 2930 2808
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 9858 2836 9864 2848
rect 4111 2808 9864 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2498 2632 2504 2644
rect 2455 2604 2504 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 3234 2632 3240 2644
rect 2648 2604 3240 2632
rect 2648 2592 2654 2604
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3786 2592 3792 2644
rect 3844 2592 3850 2644
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 4522 2592 4528 2644
rect 4580 2592 4586 2644
rect 5258 2592 5264 2644
rect 5316 2592 5322 2644
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 6546 2632 6552 2644
rect 5675 2604 6552 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 6822 2592 6828 2644
rect 6880 2592 6886 2644
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 9214 2592 9220 2644
rect 9272 2592 9278 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10459 2604 10916 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 3513 2567 3571 2573
rect 1912 2536 3464 2564
rect 1912 2524 1918 2536
rect 566 2456 572 2508
rect 624 2496 630 2508
rect 624 2468 3372 2496
rect 624 2456 630 2468
rect 1762 2388 1768 2440
rect 1820 2388 1826 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 2004 2400 2145 2428
rect 2004 2388 2010 2400
rect 2133 2397 2145 2400
rect 2179 2428 2191 2431
rect 2406 2428 2412 2440
rect 2179 2400 2412 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2498 2388 2504 2440
rect 2556 2388 2562 2440
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2866 2428 2872 2440
rect 2639 2400 2872 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 3344 2437 3372 2468
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3436 2428 3464 2536
rect 3513 2533 3525 2567
rect 3559 2564 3571 2567
rect 3878 2564 3884 2576
rect 3559 2536 3884 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4448 2564 4476 2592
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4448 2536 4813 2564
rect 4801 2533 4813 2536
rect 4847 2533 4859 2567
rect 4801 2527 4859 2533
rect 5276 2496 5304 2592
rect 10888 2576 10916 2604
rect 10870 2524 10876 2576
rect 10928 2524 10934 2576
rect 4724 2468 5304 2496
rect 4724 2440 4752 2468
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3436 2400 3985 2428
rect 3329 2391 3387 2397
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4246 2388 4252 2440
rect 4304 2388 4310 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 4982 2388 4988 2440
rect 5040 2388 5046 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 992 2332 1409 2360
rect 992 2320 998 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2041 2363 2099 2369
rect 2041 2329 2053 2363
rect 2087 2360 2099 2363
rect 2682 2360 2688 2372
rect 2087 2332 2688 2360
rect 2087 2329 2099 2332
rect 2041 2323 2099 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 10244 2360 10272 2391
rect 2792 2332 10272 2360
rect 2792 2301 2820 2332
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3970 2292 3976 2304
rect 3283 2264 3976 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 5534 2292 5540 2304
rect 4479 2264 5540 2292
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 10042 2252 10048 2304
rect 10100 2252 10106 2304
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 2406 2048 2412 2100
rect 2464 2088 2470 2100
rect 4706 2088 4712 2100
rect 2464 2060 4712 2088
rect 2464 2048 2470 2060
rect 4706 2048 4712 2060
rect 4764 2048 4770 2100
rect 2130 1980 2136 2032
rect 2188 2020 2194 2032
rect 4982 2020 4988 2032
rect 2188 1992 4988 2020
rect 2188 1980 2194 1992
rect 4982 1980 4988 1992
rect 5040 1980 5046 2032
<< via1 >>
rect 5724 10072 5776 10124
rect 9864 10072 9916 10124
rect 4252 9936 4304 9988
rect 7932 9936 7984 9988
rect 4344 9868 4396 9920
rect 6920 9868 6972 9920
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 756 9664 808 9716
rect 940 9596 992 9648
rect 4620 9664 4672 9716
rect 6184 9664 6236 9716
rect 6276 9664 6328 9716
rect 7196 9664 7248 9716
rect 7932 9707 7984 9716
rect 7932 9673 7941 9707
rect 7941 9673 7975 9707
rect 7975 9673 7984 9707
rect 7932 9664 7984 9673
rect 8024 9664 8076 9716
rect 8668 9664 8720 9716
rect 9772 9664 9824 9716
rect 10508 9664 10560 9716
rect 1400 9392 1452 9444
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3516 9528 3568 9580
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5356 9596 5408 9648
rect 5724 9528 5776 9580
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 3240 9392 3292 9444
rect 4620 9460 4672 9512
rect 6184 9503 6236 9512
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 9864 9596 9916 9648
rect 10508 9528 10560 9580
rect 1216 9324 1268 9376
rect 2596 9324 2648 9376
rect 4344 9324 4396 9376
rect 4528 9324 4580 9376
rect 5080 9367 5132 9376
rect 5080 9333 5089 9367
rect 5089 9333 5123 9367
rect 5123 9333 5132 9367
rect 5080 9324 5132 9333
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 6736 9324 6788 9376
rect 7380 9324 7432 9376
rect 8116 9324 8168 9376
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 2780 9120 2832 9172
rect 3516 9120 3568 9172
rect 4436 9120 4488 9172
rect 5908 9120 5960 9172
rect 6920 9120 6972 9172
rect 2688 9052 2740 9104
rect 10416 9095 10468 9104
rect 10416 9061 10425 9095
rect 10425 9061 10459 9095
rect 10459 9061 10468 9095
rect 10416 9052 10468 9061
rect 11060 9052 11112 9104
rect 4528 8984 4580 9036
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5356 8984 5408 9036
rect 5540 8984 5592 9036
rect 6184 8984 6236 9036
rect 6552 8984 6604 9036
rect 2044 8916 2096 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3700 8916 3752 8968
rect 1768 8891 1820 8900
rect 1768 8857 1777 8891
rect 1777 8857 1811 8891
rect 1811 8857 1820 8891
rect 1768 8848 1820 8857
rect 2412 8848 2464 8900
rect 3884 8891 3936 8900
rect 3884 8857 3893 8891
rect 3893 8857 3927 8891
rect 3927 8857 3936 8891
rect 3884 8848 3936 8857
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 3240 8780 3292 8832
rect 4344 8848 4396 8900
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 4896 8848 4948 8900
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 4252 8780 4304 8832
rect 5172 8780 5224 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 8668 8780 8720 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 2872 8508 2924 8560
rect 4988 8576 5040 8628
rect 5632 8576 5684 8628
rect 1952 8440 2004 8492
rect 3056 8440 3108 8492
rect 3240 8440 3292 8492
rect 4896 8508 4948 8560
rect 5540 8508 5592 8560
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 8668 8576 8720 8628
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 9312 8576 9364 8628
rect 8116 8508 8168 8560
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 6828 8279 6880 8288
rect 6828 8245 6837 8279
rect 6837 8245 6871 8279
rect 6871 8245 6880 8279
rect 6828 8236 6880 8245
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 10508 8236 10560 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 1952 8032 2004 8084
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 3884 8032 3936 8084
rect 1400 7828 1452 7880
rect 2044 7828 2096 7880
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3976 7828 4028 7880
rect 5080 8032 5132 8084
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10232 8032 10284 8084
rect 7656 7964 7708 8016
rect 5172 7896 5224 7948
rect 1308 7760 1360 7812
rect 4160 7803 4212 7812
rect 4160 7769 4169 7803
rect 4169 7769 4203 7803
rect 4203 7769 4212 7803
rect 4160 7760 4212 7769
rect 4988 7828 5040 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6828 7828 6880 7880
rect 8392 7896 8444 7948
rect 4252 7692 4304 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 10324 7692 10376 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 1952 7488 2004 7540
rect 2596 7488 2648 7540
rect 3240 7488 3292 7540
rect 4160 7488 4212 7540
rect 6460 7488 6512 7540
rect 8024 7488 8076 7540
rect 8668 7488 8720 7540
rect 2596 7395 2648 7404
rect 2596 7361 2614 7395
rect 2614 7361 2648 7395
rect 2596 7352 2648 7361
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 4068 7352 4120 7404
rect 4160 7352 4212 7404
rect 2964 7284 3016 7336
rect 3792 7284 3844 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 5540 7284 5592 7336
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 7380 7284 7432 7336
rect 7656 7284 7708 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10324 7284 10376 7336
rect 2504 7148 2556 7200
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 5816 7148 5868 7200
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 2872 6944 2924 6996
rect 3148 6808 3200 6860
rect 7564 6944 7616 6996
rect 9404 6987 9456 6996
rect 4344 6876 4396 6928
rect 5448 6919 5500 6928
rect 5448 6885 5457 6919
rect 5457 6885 5491 6919
rect 5491 6885 5500 6919
rect 5448 6876 5500 6885
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 5540 6740 5592 6792
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 8116 6740 8168 6792
rect 8852 6808 8904 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 2780 6672 2832 6724
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 3056 6672 3108 6681
rect 4068 6672 4120 6724
rect 4436 6672 4488 6724
rect 6552 6672 6604 6724
rect 6920 6672 6972 6724
rect 1676 6604 1728 6656
rect 4896 6647 4948 6656
rect 4896 6613 4905 6647
rect 4905 6613 4939 6647
rect 4939 6613 4948 6647
rect 4896 6604 4948 6613
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 9220 6604 9272 6656
rect 10048 6604 10100 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 2596 6400 2648 6452
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 5448 6400 5500 6452
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 4896 6332 4948 6384
rect 940 6264 992 6316
rect 3792 6264 3844 6316
rect 1676 6196 1728 6248
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 3976 6196 4028 6248
rect 4252 6239 4304 6248
rect 4252 6205 4261 6239
rect 4261 6205 4295 6239
rect 4295 6205 4304 6239
rect 4252 6196 4304 6205
rect 8116 6264 8168 6316
rect 9128 6264 9180 6316
rect 10140 6264 10192 6316
rect 3240 6128 3292 6180
rect 5540 6196 5592 6248
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 8852 6196 8904 6248
rect 8944 6196 8996 6248
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 3148 6060 3200 6112
rect 6460 6103 6512 6112
rect 6460 6069 6469 6103
rect 6469 6069 6503 6103
rect 6503 6069 6512 6103
rect 6460 6060 6512 6069
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3884 5856 3936 5908
rect 5632 5856 5684 5908
rect 9128 5856 9180 5908
rect 2872 5652 2924 5704
rect 3332 5720 3384 5772
rect 1492 5516 1544 5568
rect 3792 5652 3844 5704
rect 5172 5720 5224 5772
rect 6460 5720 6512 5772
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 8852 5788 8904 5840
rect 9220 5788 9272 5840
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5724 5652 5776 5704
rect 7932 5652 7984 5704
rect 8944 5720 8996 5772
rect 9220 5652 9272 5704
rect 3240 5516 3292 5568
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9496 5584 9548 5636
rect 9956 5584 10008 5636
rect 10508 5627 10560 5636
rect 10508 5593 10517 5627
rect 10517 5593 10551 5627
rect 10551 5593 10560 5627
rect 10508 5584 10560 5593
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 2504 5312 2556 5364
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 3332 5312 3384 5364
rect 4068 5312 4120 5364
rect 6184 5312 6236 5364
rect 6276 5312 6328 5364
rect 9404 5312 9456 5364
rect 9496 5312 9548 5364
rect 9588 5312 9640 5364
rect 9864 5312 9916 5364
rect 10232 5312 10284 5364
rect 1676 5176 1728 5228
rect 940 5108 992 5160
rect 5264 5244 5316 5296
rect 2688 5176 2740 5228
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 6828 5176 6880 5228
rect 2964 5108 3016 5160
rect 5080 5108 5132 5160
rect 5540 5108 5592 5160
rect 6552 5108 6604 5160
rect 9220 5176 9272 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 3056 5040 3108 5092
rect 4988 5083 5040 5092
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 4988 5040 5040 5049
rect 4068 4972 4120 5024
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 9956 4972 10008 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 1032 4768 1084 4820
rect 3332 4768 3384 4820
rect 3792 4768 3844 4820
rect 4436 4768 4488 4820
rect 4988 4768 5040 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 3884 4700 3936 4752
rect 4252 4700 4304 4752
rect 5448 4768 5500 4820
rect 6552 4768 6604 4820
rect 6920 4768 6972 4820
rect 7656 4768 7708 4820
rect 8484 4768 8536 4820
rect 10232 4768 10284 4820
rect 2504 4564 2556 4616
rect 2688 4564 2740 4616
rect 3240 4564 3292 4616
rect 3332 4564 3384 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 8944 4632 8996 4684
rect 3056 4496 3108 4548
rect 5448 4496 5500 4548
rect 6552 4496 6604 4548
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 2688 4224 2740 4276
rect 3056 4224 3108 4276
rect 3884 4224 3936 4276
rect 4436 4224 4488 4276
rect 5172 4224 5224 4276
rect 1952 4156 2004 4208
rect 3240 4088 3292 4140
rect 3976 4088 4028 4140
rect 5448 4088 5500 4140
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 4252 4063 4304 4072
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 6736 4020 6788 4072
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 3976 3952 4028 4004
rect 4528 3952 4580 4004
rect 2596 3884 2648 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 940 3680 992 3732
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 3792 3680 3844 3732
rect 4252 3680 4304 3732
rect 4436 3544 4488 3596
rect 1676 3476 1728 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 1032 3340 1084 3392
rect 3148 3408 3200 3460
rect 2228 3340 2280 3392
rect 3424 3408 3476 3460
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 3884 3340 3936 3392
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 2780 3136 2832 3188
rect 2872 3136 2924 3188
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 10232 3136 10284 3188
rect 10324 3136 10376 3188
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2596 3068 2648 3120
rect 1952 2864 2004 2916
rect 4528 3068 4580 3120
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2872 2796 2924 2848
rect 3240 3000 3292 3052
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4068 3000 4120 3052
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 8024 3000 8076 3052
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 3976 2932 4028 2984
rect 10140 2932 10192 2984
rect 3700 2796 3752 2848
rect 9864 2796 9916 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 2504 2592 2556 2644
rect 2596 2592 2648 2644
rect 3240 2592 3292 2644
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4436 2592 4488 2644
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 5264 2592 5316 2644
rect 6552 2592 6604 2644
rect 6828 2635 6880 2644
rect 6828 2601 6837 2635
rect 6837 2601 6871 2635
rect 6871 2601 6880 2635
rect 6828 2592 6880 2601
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 1860 2524 1912 2576
rect 572 2456 624 2508
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 1952 2388 2004 2440
rect 2412 2388 2464 2440
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 2872 2388 2924 2440
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3884 2524 3936 2576
rect 10876 2524 10928 2576
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 940 2320 992 2372
rect 2688 2320 2740 2372
rect 3976 2252 4028 2304
rect 5540 2252 5592 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 2412 2048 2464 2100
rect 4712 2048 4764 2100
rect 2136 1980 2188 2032
rect 4988 1980 5040 2032
<< metal2 >>
rect 754 11200 810 12000
rect 2042 11200 2098 12000
rect 2870 11248 2926 11257
rect 768 9722 796 11200
rect 756 9716 808 9722
rect 756 9658 808 9664
rect 940 9648 992 9654
rect 938 9616 940 9625
rect 992 9616 994 9625
rect 938 9551 994 9560
rect 1400 9444 1452 9450
rect 1400 9386 1452 9392
rect 1216 9376 1268 9382
rect 1216 9318 1268 9324
rect 1228 8809 1256 9318
rect 1214 8800 1270 8809
rect 1214 8735 1270 8744
rect 1412 7886 1440 9386
rect 2056 8974 2084 11200
rect 3330 11200 3386 12000
rect 4618 11200 4674 12000
rect 5906 11200 5962 12000
rect 6012 11206 6224 11234
rect 2870 11183 2926 11192
rect 2778 10432 2834 10441
rect 2778 10367 2834 10376
rect 2134 9616 2190 9625
rect 2134 9551 2136 9560
rect 2188 9551 2190 9560
rect 2688 9580 2740 9586
rect 2136 9522 2188 9528
rect 2688 9522 2740 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2410 9072 2466 9081
rect 2410 9007 2466 9016
rect 2044 8968 2096 8974
rect 1766 8936 1822 8945
rect 2044 8910 2096 8916
rect 2424 8906 2452 9007
rect 1766 8871 1768 8880
rect 1820 8871 1822 8880
rect 2412 8900 2464 8906
rect 1768 8842 1820 8848
rect 2412 8842 2464 8848
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8265 1532 8774
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1964 8090 1992 8434
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1320 7177 1348 7754
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1306 7168 1362 7177
rect 1306 7103 1362 7112
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 938 6352 994 6361
rect 938 6287 940 6296
rect 992 6287 994 6296
rect 940 6258 992 6264
rect 1688 6254 1716 6598
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1492 5568 1544 5574
rect 1030 5536 1086 5545
rect 1492 5510 1544 5516
rect 1030 5471 1086 5480
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 1044 4826 1072 5471
rect 1032 4820 1084 4826
rect 1032 4762 1084 4768
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 938 3904 994 3913
rect 938 3839 994 3848
rect 952 3738 980 3839
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 1032 3392 1084 3398
rect 1032 3334 1084 3340
rect 1044 3097 1072 3334
rect 1030 3088 1086 3097
rect 1504 3058 1532 5510
rect 1688 5234 1716 6190
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 3534 1716 5170
rect 1964 4214 1992 7482
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1964 3058 1992 4150
rect 1030 3023 1086 3032
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 572 2508 624 2514
rect 572 2450 624 2456
rect 584 800 612 2450
rect 1780 2446 1808 2790
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2281 980 2314
rect 938 2272 994 2281
rect 938 2207 994 2216
rect 1872 1306 1900 2518
rect 1964 2446 1992 2858
rect 2056 2530 2084 7822
rect 2516 7206 2544 7822
rect 2608 7546 2636 9318
rect 2700 9110 2728 9522
rect 2792 9178 2820 10367
rect 2884 9586 2912 11183
rect 3344 10146 3372 11200
rect 3252 10118 3372 10146
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 3252 9450 3280 10118
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3528 9178 3556 9522
rect 3698 9480 3754 9489
rect 3698 9415 3754 9424
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 3712 8974 3740 9415
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8650 2912 8774
rect 2792 8622 2912 8650
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2516 5370 2544 7142
rect 2608 6458 2636 7346
rect 2792 6882 2820 8622
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2884 7410 2912 8502
rect 3068 8498 3096 8910
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8498 3280 8774
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3896 8090 3924 8842
rect 4264 8838 4292 9930
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 9654 4384 9862
rect 4632 9722 4660 11200
rect 5920 11098 5948 11200
rect 6012 11098 6040 11206
rect 5920 11070 6040 11098
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4620 9512 4672 9518
rect 4448 9460 4620 9466
rect 4448 9454 4672 9460
rect 4448 9438 4660 9454
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 8906 4384 9318
rect 4448 9178 4476 9438
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4540 9042 4568 9318
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 5000 9042 5028 9522
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4908 8566 4936 8842
rect 5000 8634 5028 8978
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3252 7546 3280 8026
rect 5000 7886 5028 8570
rect 5092 8090 5120 9318
rect 5368 9042 5396 9590
rect 5736 9586 5764 10066
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6196 9722 6224 11206
rect 7194 11200 7250 12000
rect 8482 11200 8538 12000
rect 9770 11200 9826 12000
rect 11058 11200 11114 12000
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 9042 5580 9318
rect 5736 9058 5764 9522
rect 5920 9178 5948 9522
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5644 9030 5764 9058
rect 6196 9042 6224 9454
rect 6184 9036 6236 9042
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7954 5212 8774
rect 5552 8566 5580 8774
rect 5644 8634 5672 9030
rect 6184 8978 6236 8984
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5736 8090 5764 8910
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 7002 2912 7346
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2700 6854 2820 6882
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6338 2728 6854
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2792 6458 2820 6666
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2700 6310 2820 6338
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2516 4622 2544 5306
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2700 4622 2728 5170
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4282 2728 4558
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2792 4162 2820 6310
rect 2884 5710 2912 6938
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5370 2912 5646
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2976 5166 3004 7278
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3068 5098 3096 6666
rect 3160 6118 3188 6802
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3804 6322 3832 7278
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3056 5092 3108 5098
rect 3056 5034 3108 5040
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3068 4282 3096 4490
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2792 4134 3096 4162
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3194 2268 3334
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2516 2650 2544 4014
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3126 2636 3878
rect 2792 3194 2820 4014
rect 3068 3618 3096 4134
rect 3160 4010 3188 6054
rect 3252 5914 3280 6122
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3344 5778 3372 6190
rect 3896 5914 3924 7278
rect 3988 6338 4016 7822
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4172 7546 4200 7754
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4080 6730 4108 7346
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3988 6310 4108 6338
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 4706 3280 5510
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3344 4826 3372 5306
rect 3804 4826 3832 5646
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3884 4752 3936 4758
rect 3252 4678 3372 4706
rect 3884 4694 3936 4700
rect 3344 4622 3372 4678
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3252 4264 3280 4558
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3252 4236 3372 4264
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3252 3738 3280 4082
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3068 3590 3280 3618
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2884 3194 2912 3470
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2596 3120 2648 3126
rect 3068 3074 3096 3470
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3160 3194 3188 3402
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2596 3062 2648 3068
rect 2792 3046 3096 3074
rect 3252 3058 3280 3590
rect 3344 3482 3372 4236
rect 3804 3738 3832 4558
rect 3896 4282 3924 4694
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 4146 4016 6190
rect 4080 5370 4108 6310
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3344 3466 3464 3482
rect 3344 3460 3476 3466
rect 3344 3454 3424 3460
rect 3424 3402 3476 3408
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3896 3058 3924 3334
rect 3240 3052 3292 3058
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2608 2530 2636 2586
rect 2056 2502 2176 2530
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2148 2038 2176 2502
rect 2516 2502 2636 2530
rect 2516 2446 2544 2502
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2504 2440 2556 2446
rect 2792 2394 2820 3046
rect 3240 2994 3292 3000
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2446 2912 2790
rect 3252 2650 3280 2994
rect 3700 2848 3752 2854
rect 3752 2796 3832 2802
rect 3700 2790 3832 2796
rect 3712 2774 3832 2790
rect 3804 2650 3832 2774
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3896 2582 3924 2994
rect 3988 2990 4016 3946
rect 4080 3058 4108 4966
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 2504 2382 2556 2388
rect 2424 2106 2452 2382
rect 2700 2378 2820 2394
rect 2872 2440 2924 2446
rect 3056 2440 3108 2446
rect 2872 2382 2924 2388
rect 2976 2400 3056 2428
rect 2688 2372 2820 2378
rect 2740 2366 2820 2372
rect 2688 2314 2740 2320
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 2136 2032 2188 2038
rect 2136 1974 2188 1980
rect 1780 1278 1900 1306
rect 1780 800 1808 1278
rect 2976 800 3004 2400
rect 3056 2382 3108 2388
rect 3988 2310 4016 2926
rect 4172 2774 4200 7346
rect 4264 6338 4292 7686
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 6934 4384 7142
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 4356 6458 4384 6870
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4264 6310 4384 6338
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 4758 4292 6190
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4078 4292 4558
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4264 3738 4292 4014
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4356 3058 4384 6310
rect 4448 4826 4476 6666
rect 4632 6202 4660 6734
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6390 4936 6598
rect 5460 6458 5488 6870
rect 5552 6798 5580 7278
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4540 6174 4660 6202
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 4282 4476 4558
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4540 4010 4568 6174
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5234 5212 5714
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5276 5302 5304 5646
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 5000 4826 5028 5034
rect 5092 4826 5120 5102
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5184 4282 5212 5170
rect 5552 5166 5580 6190
rect 5644 5914 5672 6734
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5710 5764 7142
rect 5828 6798 5856 7142
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6196 5370 6224 6190
rect 6288 5370 6316 9658
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 8634 6408 9522
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6564 9042 6592 9318
rect 6748 9081 6776 9318
rect 6932 9178 6960 9862
rect 7208 9722 7236 11200
rect 8496 10282 8524 11200
rect 8496 10254 8708 10282
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7944 9722 7972 9930
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8680 9722 8708 10254
rect 9784 9722 9812 11200
rect 10506 10432 10562 10441
rect 10506 10367 10562 10376
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 7654 9616 7710 9625
rect 7564 9580 7616 9586
rect 7654 9551 7656 9560
rect 7564 9522 7616 9528
rect 7708 9551 7710 9560
rect 7840 9580 7892 9586
rect 7656 9522 7708 9528
rect 7840 9522 7892 9528
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6734 9072 6790 9081
rect 6552 9036 6604 9042
rect 6734 9007 6790 9016
rect 6552 8978 6604 8984
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7886 6868 8230
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6472 7546 6500 7822
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6564 6730 6592 7686
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6472 5778 6500 6054
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4826 5488 4966
rect 6564 4826 6592 5102
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5184 4154 5212 4218
rect 5184 4126 5304 4154
rect 5460 4146 5488 4490
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4080 2746 4200 2774
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 4080 1465 4108 2746
rect 4448 2650 4476 3538
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4540 2650 4568 3062
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 5276 2650 5304 4126
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 4264 1306 4292 2382
rect 4724 2106 4752 2382
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 5000 2038 5028 2382
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 5460 1306 5488 2382
rect 5552 2310 5580 4082
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 6564 2650 6592 4490
rect 6656 4154 6684 7346
rect 7392 7342 7420 9318
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7576 7002 7604 9522
rect 7852 9489 7880 9522
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7668 7342 7696 7958
rect 8036 7546 8064 9658
rect 9876 9654 9904 10066
rect 10520 9722 10548 10367
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10506 9616 10562 9625
rect 10506 9551 10508 9560
rect 10560 9551 10562 9560
rect 10508 9522 10560 9528
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8128 8566 8156 9318
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8680 8634 8708 8774
rect 9232 8634 9260 8871
rect 9324 8634 9352 9318
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 11072 9110 11100 11200
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10232 8968 10284 8974
rect 10428 8945 10456 9046
rect 10232 8910 10284 8916
rect 10414 8936 10470 8945
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 7732 8248 8366
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7954 8432 8230
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 10152 8090 10180 8434
rect 10244 8090 10272 8910
rect 10414 8871 10470 8880
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10520 7993 10548 8230
rect 10506 7984 10562 7993
rect 8392 7948 8444 7954
rect 10506 7919 10562 7928
rect 8392 7890 8444 7896
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 8128 7704 8248 7732
rect 8668 7744 8720 7750
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 5778 6960 6666
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6656 4126 6776 4154
rect 6748 4078 6776 4126
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6840 2650 6868 5170
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4826 6960 4966
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7668 4826 7696 7278
rect 8128 6798 8156 7704
rect 8668 7686 8720 7692
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8680 7546 8708 7686
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8956 6866 8984 7686
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6322 8156 6734
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8864 6254 8892 6802
rect 9232 6662 9260 7278
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 7002 9444 7142
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5710 7972 6054
rect 8864 5846 8892 6190
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8956 5778 8984 6190
rect 9140 5914 9168 6258
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 9232 5710 9260 5782
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8496 4826 8524 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8956 4690 8984 5510
rect 9416 5370 9444 6190
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5370 9536 5578
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5370 9628 5510
rect 9876 5370 9904 6734
rect 10060 6662 10088 7822
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6458 10088 6598
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 8036 2650 8064 2994
rect 9232 2650 9260 5170
rect 9968 5030 9996 5578
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 10152 2990 10180 6258
rect 10244 5370 10272 7346
rect 10336 7342 10364 7686
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 4826 10272 5170
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3194 10272 3470
rect 10336 3194 10364 7278
rect 10416 7200 10468 7206
rect 10414 7168 10416 7177
rect 10468 7168 10470 7177
rect 10414 7103 10470 7112
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10428 6361 10456 6394
rect 10414 6352 10470 6361
rect 10414 6287 10470 6296
rect 10506 5672 10562 5681
rect 10506 5607 10508 5616
rect 10560 5607 10562 5616
rect 10508 5578 10560 5584
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4729 10456 4966
rect 10414 4720 10470 4729
rect 10414 4655 10470 4664
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10416 3936 10468 3942
rect 10414 3904 10416 3913
rect 10468 3904 10470 3913
rect 10414 3839 10470 3848
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10428 3097 10456 3334
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10414 3088 10470 3097
rect 10232 3052 10284 3058
rect 10414 3023 10470 3032
rect 10232 2994 10284 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9876 2446 9904 2790
rect 10244 2774 10272 2994
rect 10152 2746 10272 2774
rect 6644 2440 6696 2446
rect 7840 2440 7892 2446
rect 6644 2382 6696 2388
rect 7760 2400 7840 2428
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6656 1306 6684 2382
rect 4172 1278 4292 1306
rect 5368 1278 5488 1306
rect 6564 1278 6684 1306
rect 4172 800 4200 1278
rect 5368 800 5396 1278
rect 6564 800 6592 1278
rect 7760 800 7788 2400
rect 9036 2440 9088 2446
rect 7840 2382 7892 2388
rect 8956 2400 9036 2428
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8956 800 8984 2400
rect 9036 2382 9088 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10060 1465 10088 2246
rect 10046 1456 10102 1465
rect 10046 1391 10102 1400
rect 10152 800 10180 2746
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10888 2417 10916 2518
rect 10874 2408 10930 2417
rect 10874 2343 10930 2352
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
<< via2 >>
rect 938 9596 940 9616
rect 940 9596 992 9616
rect 992 9596 994 9616
rect 938 9560 994 9596
rect 1214 8744 1270 8800
rect 2870 11192 2926 11248
rect 2778 10376 2834 10432
rect 2134 9580 2190 9616
rect 2134 9560 2136 9580
rect 2136 9560 2188 9580
rect 2188 9560 2190 9580
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 2410 9016 2466 9072
rect 1766 8900 1822 8936
rect 1766 8880 1768 8900
rect 1768 8880 1820 8900
rect 1820 8880 1822 8900
rect 1490 8200 1546 8256
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 1306 7112 1362 7168
rect 938 6316 994 6352
rect 938 6296 940 6316
rect 940 6296 992 6316
rect 992 6296 994 6316
rect 1030 5480 1086 5536
rect 938 4664 994 4720
rect 938 3848 994 3904
rect 1030 3032 1086 3088
rect 938 2216 994 2272
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 3698 9424 3754 9480
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 10506 10376 10562 10432
rect 7654 9580 7710 9616
rect 7654 9560 7656 9580
rect 7656 9560 7708 9580
rect 7708 9560 7710 9580
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 6734 9016 6790 9072
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 4066 1400 4122 1456
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7838 9424 7894 9480
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10506 9580 10562 9616
rect 10506 9560 10508 9580
rect 10508 9560 10560 9580
rect 10560 9560 10562 9580
rect 9218 8880 9274 8936
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10414 8880 10470 8936
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10506 7928 10562 7984
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10414 7148 10416 7168
rect 10416 7148 10468 7168
rect 10468 7148 10470 7168
rect 10414 7112 10470 7148
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10414 6296 10470 6352
rect 10506 5636 10562 5672
rect 10506 5616 10508 5636
rect 10508 5616 10560 5636
rect 10560 5616 10562 5636
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10414 4664 10470 4720
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10414 3884 10416 3904
rect 10416 3884 10468 3904
rect 10468 3884 10470 3904
rect 10414 3848 10470 3884
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 10414 3032 10470 3088
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10046 1400 10102 1456
rect 10874 2352 10930 2408
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
<< metal3 >>
rect 0 11250 800 11280
rect 2865 11250 2931 11253
rect 0 11248 2931 11250
rect 0 11192 2870 11248
rect 2926 11192 2931 11248
rect 0 11190 2931 11192
rect 0 11160 800 11190
rect 2865 11187 2931 11190
rect 0 10434 800 10464
rect 2773 10434 2839 10437
rect 0 10432 2839 10434
rect 0 10376 2778 10432
rect 2834 10376 2839 10432
rect 0 10374 2839 10376
rect 0 10344 800 10374
rect 2773 10371 2839 10374
rect 10501 10434 10567 10437
rect 11200 10434 12000 10464
rect 10501 10432 12000 10434
rect 10501 10376 10506 10432
rect 10562 10376 12000 10432
rect 10501 10374 12000 10376
rect 10501 10371 10567 10374
rect 11200 10344 12000 10374
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 0 9618 800 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 2129 9618 2195 9621
rect 7649 9618 7715 9621
rect 2129 9616 7715 9618
rect 2129 9560 2134 9616
rect 2190 9560 7654 9616
rect 7710 9560 7715 9616
rect 2129 9558 7715 9560
rect 2129 9555 2195 9558
rect 7649 9555 7715 9558
rect 10501 9618 10567 9621
rect 11200 9618 12000 9648
rect 10501 9616 12000 9618
rect 10501 9560 10506 9616
rect 10562 9560 12000 9616
rect 10501 9558 12000 9560
rect 10501 9555 10567 9558
rect 11200 9528 12000 9558
rect 3693 9482 3759 9485
rect 7833 9482 7899 9485
rect 3693 9480 7899 9482
rect 3693 9424 3698 9480
rect 3754 9424 7838 9480
rect 7894 9424 7899 9480
rect 3693 9422 7899 9424
rect 3693 9419 3759 9422
rect 7833 9419 7899 9422
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 2405 9074 2471 9077
rect 6729 9074 6795 9077
rect 2405 9072 6795 9074
rect 2405 9016 2410 9072
rect 2466 9016 6734 9072
rect 6790 9016 6795 9072
rect 2405 9014 6795 9016
rect 2405 9011 2471 9014
rect 6729 9011 6795 9014
rect 1761 8938 1827 8941
rect 9213 8938 9279 8941
rect 1761 8936 9279 8938
rect 1761 8880 1766 8936
rect 1822 8880 9218 8936
rect 9274 8880 9279 8936
rect 1761 8878 9279 8880
rect 1761 8875 1827 8878
rect 9213 8875 9279 8878
rect 10409 8938 10475 8941
rect 10409 8936 11162 8938
rect 10409 8880 10414 8936
rect 10470 8880 11162 8936
rect 10409 8878 11162 8880
rect 10409 8875 10475 8878
rect 11102 8836 11162 8878
rect 11102 8832 11346 8836
rect 0 8802 800 8832
rect 1209 8802 1275 8805
rect 0 8800 1275 8802
rect 0 8744 1214 8800
rect 1270 8744 1275 8800
rect 11102 8776 12000 8832
rect 0 8742 1275 8744
rect 0 8712 800 8742
rect 1209 8739 1275 8742
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 11200 8712 12000 8776
rect 10698 8671 11014 8672
rect 1485 8258 1551 8261
rect 798 8256 1551 8258
rect 798 8200 1490 8256
rect 1546 8200 1551 8256
rect 798 8198 1551 8200
rect 798 8016 858 8198
rect 1485 8195 1551 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7926 858 8016
rect 10501 7986 10567 7989
rect 11200 7986 12000 8016
rect 10501 7984 12000 7986
rect 10501 7928 10506 7984
rect 10562 7928 12000 7984
rect 10501 7926 12000 7928
rect 0 7896 800 7926
rect 10501 7923 10567 7926
rect 11200 7896 12000 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 0 7170 800 7200
rect 1301 7170 1367 7173
rect 0 7168 1367 7170
rect 0 7112 1306 7168
rect 1362 7112 1367 7168
rect 0 7110 1367 7112
rect 0 7080 800 7110
rect 1301 7107 1367 7110
rect 10409 7170 10475 7173
rect 11200 7170 12000 7200
rect 10409 7168 12000 7170
rect 10409 7112 10414 7168
rect 10470 7112 12000 7168
rect 10409 7110 12000 7112
rect 10409 7107 10475 7110
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 11200 7080 12000 7110
rect 9479 7039 9795 7040
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 10409 6354 10475 6357
rect 11200 6354 12000 6384
rect 10409 6352 12000 6354
rect 10409 6296 10414 6352
rect 10470 6296 12000 6352
rect 10409 6294 12000 6296
rect 10409 6291 10475 6294
rect 11200 6264 12000 6294
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 10501 5674 10567 5677
rect 10501 5672 11162 5674
rect 10501 5616 10506 5672
rect 10562 5616 11162 5672
rect 10501 5614 11162 5616
rect 10501 5611 10567 5614
rect 11102 5572 11162 5614
rect 11102 5568 11346 5572
rect 0 5538 800 5568
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 11102 5512 12000 5568
rect 0 5478 1091 5480
rect 0 5448 800 5478
rect 1025 5475 1091 5478
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 11200 5448 12000 5512
rect 10698 5407 11014 5408
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 10409 4722 10475 4725
rect 11200 4722 12000 4752
rect 10409 4720 12000 4722
rect 10409 4664 10414 4720
rect 10470 4664 12000 4720
rect 10409 4662 12000 4664
rect 10409 4659 10475 4662
rect 11200 4632 12000 4662
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 10409 3906 10475 3909
rect 11200 3906 12000 3936
rect 10409 3904 12000 3906
rect 10409 3848 10414 3904
rect 10470 3848 12000 3904
rect 10409 3846 12000 3848
rect 10409 3843 10475 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 11200 3816 12000 3846
rect 9479 3775 9795 3776
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 0 3090 800 3120
rect 1025 3090 1091 3093
rect 0 3088 1091 3090
rect 0 3032 1030 3088
rect 1086 3032 1091 3088
rect 0 3030 1091 3032
rect 0 3000 800 3030
rect 1025 3027 1091 3030
rect 10409 3090 10475 3093
rect 11200 3090 12000 3120
rect 10409 3088 12000 3090
rect 10409 3032 10414 3088
rect 10470 3032 12000 3088
rect 10409 3030 12000 3032
rect 10409 3027 10475 3030
rect 11200 3000 12000 3030
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 10869 2410 10935 2413
rect 10869 2408 11162 2410
rect 10869 2352 10874 2408
rect 10930 2352 11162 2408
rect 10869 2350 11162 2352
rect 10869 2347 10935 2350
rect 11102 2308 11162 2350
rect 11102 2304 11346 2308
rect 0 2274 800 2304
rect 933 2274 999 2277
rect 0 2272 999 2274
rect 0 2216 938 2272
rect 994 2216 999 2272
rect 11102 2248 12000 2304
rect 0 2214 999 2216
rect 0 2184 800 2214
rect 933 2211 999 2214
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 11200 2184 12000 2248
rect 10698 2143 11014 2144
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 10041 1458 10107 1461
rect 11200 1458 12000 1488
rect 10041 1456 12000 1458
rect 10041 1400 10046 1456
rect 10102 1400 12000 1456
rect 10041 1398 12000 1400
rect 10041 1395 10107 1398
rect 11200 1368 12000 1398
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform -1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform -1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform -1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform 1 0 1472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1688980957
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1688980957
transform -1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform -1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform -1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform -1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform -1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1688980957
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1688980957
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform -1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform -1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform -1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1688980957
transform -1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1688980957
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1688980957
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1688980957
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1688980957
transform -1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1688980957
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1688980957
transform -1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1688980957
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1688980957
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1688980957
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1688980957
transform -1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _119_
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 1688980957
transform -1 0 2852 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 1688980957
transform -1 0 3036 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _123_
timestamp 1688980957
transform -1 0 7912 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _125_
timestamp 1688980957
transform -1 0 2944 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _126_
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _127_
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform -1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1688980957
transform -1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform -1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1688980957
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1688980957
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1688980957
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform -1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform -1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _150__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _150_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _151_
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _152_
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _153_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _154_
timestamp 1688980957
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _155_
timestamp 1688980957
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _156_
timestamp 1688980957
transform 1 0 4232 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _157_
timestamp 1688980957
transform 1 0 6900 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _158_
timestamp 1688980957
transform -1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _159_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _160_
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _161_
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _162_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _163_
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _163__44
timestamp 1688980957
transform 1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _164_
timestamp 1688980957
transform 1 0 2576 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _165_
timestamp 1688980957
transform -1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _166_
timestamp 1688980957
transform -1 0 2576 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _167_
timestamp 1688980957
transform 1 0 2576 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _168_
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _169_
timestamp 1688980957
transform -1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _170_
timestamp 1688980957
transform -1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _171_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _172_
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _173_
timestamp 1688980957
transform -1 0 4324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _174__45
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _174_
timestamp 1688980957
transform -1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _175_
timestamp 1688980957
transform 1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _176_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _177_
timestamp 1688980957
transform -1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _178__46
timestamp 1688980957
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _178_
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _179_
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _180_
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _181_
timestamp 1688980957
transform -1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_32
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_25
timestamp 1688980957
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_36 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_98
timestamp 1688980957
transform 1 0 10120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_18
timestamp 1688980957
transform 1 0 2760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_35
timestamp 1688980957
transform 1 0 4324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_47
timestamp 1688980957
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_59
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_71
timestamp 1688980957
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_38
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_45
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_14
timestamp 1688980957
transform 1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_24
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_32
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_42
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_49
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_56
timestamp 1688980957
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1688980957
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_92
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_21
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_88
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_26
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_46
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_68
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_101
timestamp 1688980957
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_63
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_71
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_97
timestamp 1688980957
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_24
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_35
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_67
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_74
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_88
timestamp 1688980957
transform 1 0 9200 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_94
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_60
timestamp 1688980957
transform 1 0 6624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_91
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_49
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_46
timestamp 1688980957
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_66
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 7268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 10212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 2852 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output30 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1688980957
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 3404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1688980957
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal3 s 11200 9528 12000 9648 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 11200 10344 12000 10464 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 3 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 4 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 5 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 6 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 7 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 8 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 9 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 10 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 11 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 12 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 13 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 14 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 15 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 16 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 17 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 18 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 19 nsew signal tristate
flabel metal2 s 754 11200 810 12000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 20 nsew signal input
flabel metal2 s 2042 11200 2098 12000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 21 nsew signal input
flabel metal2 s 3330 11200 3386 12000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 22 nsew signal input
flabel metal2 s 4618 11200 4674 12000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 23 nsew signal input
flabel metal2 s 5906 11200 5962 12000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 24 nsew signal input
flabel metal2 s 7194 11200 7250 12000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 25 nsew signal input
flabel metal2 s 8482 11200 8538 12000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 26 nsew signal input
flabel metal2 s 9770 11200 9826 12000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 27 nsew signal input
flabel metal2 s 11058 11200 11114 12000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 28 nsew signal input
flabel metal3 s 11200 1368 12000 1488 0 FreeSans 480 0 0 0 chany_top_out[0]
port 29 nsew signal tristate
flabel metal3 s 11200 2184 12000 2304 0 FreeSans 480 0 0 0 chany_top_out[1]
port 30 nsew signal tristate
flabel metal3 s 11200 3000 12000 3120 0 FreeSans 480 0 0 0 chany_top_out[2]
port 31 nsew signal tristate
flabel metal3 s 11200 3816 12000 3936 0 FreeSans 480 0 0 0 chany_top_out[3]
port 32 nsew signal tristate
flabel metal3 s 11200 4632 12000 4752 0 FreeSans 480 0 0 0 chany_top_out[4]
port 33 nsew signal tristate
flabel metal3 s 11200 5448 12000 5568 0 FreeSans 480 0 0 0 chany_top_out[5]
port 34 nsew signal tristate
flabel metal3 s 11200 6264 12000 6384 0 FreeSans 480 0 0 0 chany_top_out[6]
port 35 nsew signal tristate
flabel metal3 s 11200 7080 12000 7200 0 FreeSans 480 0 0 0 chany_top_out[7]
port 36 nsew signal tristate
flabel metal3 s 11200 7896 12000 8016 0 FreeSans 480 0 0 0 chany_top_out[8]
port 37 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 38 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 39 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 40 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 41 nsew signal input
flabel metal3 s 11200 8712 12000 8832 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
port 42 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 3266 3638 3266 3638 0 _000_
rlabel metal1 4094 5576 4094 5576 0 _001_
rlabel metal1 3726 4794 3726 4794 0 _002_
rlabel metal1 7958 4624 7958 4624 0 _003_
rlabel metal1 5888 4590 5888 4590 0 _004_
rlabel metal1 10166 5236 10166 5236 0 _005_
rlabel metal1 7636 7854 7636 7854 0 _006_
rlabel metal1 5336 4590 5336 4590 0 _007_
rlabel metal1 8395 6902 8395 6902 0 _008_
rlabel metal1 4600 8942 4600 8942 0 _009_
rlabel metal2 6394 9078 6394 9078 0 _010_
rlabel metal2 3358 5066 3358 5066 0 _011_
rlabel metal1 4646 8568 4646 8568 0 _012_
rlabel metal2 2254 3264 2254 3264 0 _013_
rlabel metal1 2346 3060 2346 3060 0 _014_
rlabel metal1 2806 3060 2806 3060 0 _015_
rlabel metal1 8648 6970 8648 6970 0 _016_
rlabel metal2 5106 4964 5106 4964 0 _017_
rlabel metal1 9936 5338 9936 5338 0 _018_
rlabel metal1 6256 4794 6256 4794 0 _019_
rlabel metal1 8050 7922 8050 7922 0 _020_
rlabel metal1 8326 4794 8326 4794 0 _021_
rlabel metal1 4784 4250 4784 4250 0 _022_
rlabel metal1 7452 4590 7452 4590 0 _023_
rlabel metal1 8464 7310 8464 7310 0 _024_
rlabel metal1 7774 5202 7774 5202 0 _025_
rlabel metal1 8786 6630 8786 6630 0 _026_
rlabel metal1 8924 5882 8924 5882 0 _027_
rlabel metal2 4462 5746 4462 5746 0 _028_
rlabel metal1 3772 5882 3772 5882 0 _029_
rlabel metal2 2806 3604 2806 3604 0 _030_
rlabel metal1 5428 5882 5428 5882 0 _031_
rlabel metal1 2622 2992 2622 2992 0 _032_
rlabel metal1 3634 3366 3634 3366 0 _033_
rlabel metal1 1932 5270 1932 5270 0 _034_
rlabel metal2 3266 6018 3266 6018 0 _035_
rlabel metal1 3726 4114 3726 4114 0 _036_
rlabel metal1 5428 5134 5428 5134 0 _037_
rlabel metal1 2392 2346 2392 2346 0 _038_
rlabel metal1 4278 4114 4278 4114 0 _039_
rlabel metal2 4370 9758 4370 9758 0 _040_
rlabel metal1 2806 7956 2806 7956 0 _041_
rlabel metal1 4002 8840 4002 8840 0 _042_
rlabel metal2 2990 6222 2990 6222 0 _043_
rlabel metal1 6624 9010 6624 9010 0 _044_
rlabel metal1 5244 7922 5244 7922 0 _045_
rlabel metal1 5750 9010 5750 9010 0 _046_
rlabel metal1 6302 7820 6302 7820 0 _047_
rlabel metal1 9798 9520 9798 9520 0 ccff_head
rlabel metal1 10488 9690 10488 9690 0 ccff_tail
rlabel metal2 598 1622 598 1622 0 chany_bottom_in[0]
rlabel metal2 1794 1027 1794 1027 0 chany_bottom_in[1]
rlabel metal2 2990 1588 2990 1588 0 chany_bottom_in[2]
rlabel metal2 4186 1027 4186 1027 0 chany_bottom_in[3]
rlabel metal2 5382 1027 5382 1027 0 chany_bottom_in[4]
rlabel metal2 6578 1027 6578 1027 0 chany_bottom_in[5]
rlabel metal2 7774 1588 7774 1588 0 chany_bottom_in[6]
rlabel metal2 8970 1588 8970 1588 0 chany_bottom_in[7]
rlabel metal2 10166 1761 10166 1761 0 chany_bottom_in[8]
rlabel metal3 820 2244 820 2244 0 chany_bottom_out[0]
rlabel metal3 866 3060 866 3060 0 chany_bottom_out[1]
rlabel metal3 820 3876 820 3876 0 chany_bottom_out[2]
rlabel metal3 820 4692 820 4692 0 chany_bottom_out[3]
rlabel metal3 866 5508 866 5508 0 chany_bottom_out[4]
rlabel metal3 820 6324 820 6324 0 chany_bottom_out[5]
rlabel metal3 1004 7140 1004 7140 0 chany_bottom_out[6]
rlabel metal3 751 7956 751 7956 0 chany_bottom_out[7]
rlabel metal3 958 8772 958 8772 0 chany_bottom_out[8]
rlabel metal2 782 10448 782 10448 0 chany_top_in[0]
rlabel metal1 2392 8942 2392 8942 0 chany_top_in[1]
rlabel metal1 1656 9554 1656 9554 0 chany_top_in[2]
rlabel metal1 5290 9588 5290 9588 0 chany_top_in[3]
rlabel metal1 6854 9588 6854 9588 0 chany_top_in[4]
rlabel metal1 7360 9554 7360 9554 0 chany_top_in[5]
rlabel metal1 8740 9554 8740 9554 0 chany_top_in[6]
rlabel metal1 9522 9588 9522 9588 0 chany_top_in[7]
rlabel metal1 10166 8976 10166 8976 0 chany_top_in[8]
rlabel metal2 10074 1853 10074 1853 0 chany_top_out[0]
rlabel metal1 10672 2618 10672 2618 0 chany_top_out[1]
rlabel metal2 10442 3213 10442 3213 0 chany_top_out[2]
rlabel via2 10442 3893 10442 3893 0 chany_top_out[3]
rlabel metal2 10442 4845 10442 4845 0 chany_top_out[4]
rlabel via2 10534 5627 10534 5627 0 chany_top_out[5]
rlabel metal2 10442 6375 10442 6375 0 chany_top_out[6]
rlabel via2 10442 7157 10442 7157 0 chany_top_out[7]
rlabel metal1 10488 8262 10488 8262 0 chany_top_out[8]
rlabel metal1 5520 5678 5520 5678 0 clknet_0_prog_clk
rlabel metal1 1886 8500 1886 8500 0 clknet_1_0__leaf_prog_clk
rlabel metal2 8188 7718 8188 7718 0 clknet_1_1__leaf_prog_clk
rlabel metal3 820 9588 820 9588 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal2 2806 9775 2806 9775 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal2 2898 10387 2898 10387 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal1 5336 4114 5336 4114 0 mem_left_ipin_0.DFF_0_.Q
rlabel metal1 8740 6222 8740 6222 0 mem_left_ipin_0.DFF_1_.Q
rlabel metal1 8602 5712 8602 5712 0 mem_left_ipin_0.DFF_2_.Q
rlabel metal1 2300 2414 2300 2414 0 mem_right_ipin_0.DFF_0_.Q
rlabel metal1 1564 5542 1564 5542 0 mem_right_ipin_0.DFF_1_.Q
rlabel metal1 1610 5202 1610 5202 0 mem_right_ipin_0.DFF_2_.Q
rlabel metal1 2438 5202 2438 5202 0 mem_right_ipin_1.DFF_0_.Q
rlabel metal1 1610 8432 1610 8432 0 mem_right_ipin_1.DFF_1_.Q
rlabel metal2 5014 9282 5014 9282 0 mem_right_ipin_2.DFF_0_.Q
rlabel metal1 4232 3706 4232 3706 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 2668 4590 2668 4590 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 6854 4590 6854 4590 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal1 6164 5134 6164 5134 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 9430 7378 9430 7378 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 8234 7854 8234 7854 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 5888 5066 5888 5066 0 mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7130 4794 7130 4794 0 mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 8510 7514 8510 7514 0 mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 9200 5338 9200 5338 0 mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 9430 7072 9430 7072 0 mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 10212 6630 10212 6630 0 mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 2944 3162 2944 3162 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal1 2484 2618 2484 2618 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal1 6164 5338 6164 5338 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal2 5842 6970 5842 6970 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 3772 4250 3772 4250 0 mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2254 4114 2254 4114 0 mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 5520 6426 5520 6426 0 mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 3404 6086 3404 6086 0 mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 4462 6868 4462 6868 0 mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 3864 6834 3864 6834 0 mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 4094 6664 4094 6664 0 mux_right_ipin_1.INVTX1_0_.out
rlabel metal1 2162 7922 2162 7922 0 mux_right_ipin_1.INVTX1_1_.out
rlabel metal1 3588 8058 3588 8058 0 mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3910 9384 3910 9384 0 mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6624 7514 6624 7514 0 mux_right_ipin_2.INVTX1_0_.out
rlabel metal1 4876 7922 4876 7922 0 mux_right_ipin_2.INVTX1_1_.out
rlabel metal2 5750 8500 5750 8500 0 mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6026 9146 6026 9146 0 mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8065 8534 8065 8534 0 net1
rlabel metal1 9982 7344 9982 7344 0 net10
rlabel metal1 1794 4148 1794 4148 0 net11
rlabel metal2 2714 6596 2714 6596 0 net12
rlabel metal2 2116 2516 2116 2516 0 net13
rlabel metal1 4416 7854 4416 7854 0 net14
rlabel metal1 5750 5236 5750 5236 0 net15
rlabel metal1 6578 7344 6578 7344 0 net16
rlabel metal1 7958 7412 7958 7412 0 net17
rlabel metal1 9384 8466 9384 8466 0 net18
rlabel metal1 8602 8466 8602 8466 0 net19
rlabel metal2 3910 2788 3910 2788 0 net2
rlabel metal1 5704 9554 5704 9554 0 net20
rlabel metal2 1794 2618 1794 2618 0 net21
rlabel metal2 3174 3298 3174 3298 0 net22
rlabel metal1 1610 3502 1610 3502 0 net23
rlabel metal1 2162 5100 2162 5100 0 net24
rlabel metal1 1794 4624 1794 4624 0 net25
rlabel metal2 4922 6494 4922 6494 0 net26
rlabel metal1 4186 7480 4186 7480 0 net27
rlabel via2 1794 8891 1794 8891 0 net28
rlabel metal1 2714 9044 2714 9044 0 net29
rlabel metal1 2760 2414 2760 2414 0 net3
rlabel metal1 6992 2822 6992 2822 0 net30
rlabel metal1 2806 2312 2806 2312 0 net31
rlabel metal2 10258 3332 10258 3332 0 net32
rlabel metal1 5750 4182 5750 4182 0 net33
rlabel metal1 9338 4726 9338 4726 0 net34
rlabel metal1 8694 4998 8694 4998 0 net35
rlabel metal1 10120 2890 10120 2890 0 net36
rlabel metal1 10120 5066 10120 5066 0 net37
rlabel metal2 10166 8262 10166 8262 0 net38
rlabel via2 2162 9571 2162 9571 0 net39
rlabel metal1 3634 2278 3634 2278 0 net4
rlabel metal1 2392 8874 2392 8874 0 net40
rlabel metal2 3542 9350 3542 9350 0 net41
rlabel metal1 10120 7990 10120 7990 0 net42
rlabel metal2 8970 7276 8970 7276 0 net43
rlabel metal2 3818 6800 3818 6800 0 net44
rlabel metal1 4462 9452 4462 9452 0 net45
rlabel metal1 6348 9010 6348 9010 0 net46
rlabel metal1 5331 8534 5331 8534 0 net47
rlabel metal1 1932 8058 1932 8058 0 net48
rlabel metal1 3532 8466 3532 8466 0 net49
rlabel metal2 5566 3196 5566 3196 0 net5
rlabel metal1 8157 6358 8157 6358 0 net50
rlabel metal1 2668 6426 2668 6426 0 net51
rlabel metal1 3082 5712 3082 5712 0 net52
rlabel metal1 7677 5678 7677 5678 0 net53
rlabel metal2 2806 6562 2806 6562 0 net54
rlabel metal1 6389 6698 6389 6698 0 net55
rlabel metal1 6118 2618 6118 2618 0 net6
rlabel metal1 6532 5202 6532 5202 0 net7
rlabel metal1 8970 3026 8970 3026 0 net8
rlabel metal1 9476 5202 9476 5202 0 net9
rlabel metal3 2384 1428 2384 1428 0 prog_clk
rlabel metal2 10442 8993 10442 8993 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
