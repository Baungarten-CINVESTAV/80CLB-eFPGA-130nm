magic
tech sky130A
magscale 1 2
timestamp 1707850947
<< viali >>
rect 4169 9673 4203 9707
rect 8217 9673 8251 9707
rect 2421 9605 2455 9639
rect 3433 9605 3467 9639
rect 5457 9605 5491 9639
rect 6837 9605 6871 9639
rect 7481 9605 7515 9639
rect 9505 9605 9539 9639
rect 10517 9605 10551 9639
rect 1501 9537 1535 9571
rect 2053 9537 2087 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 4077 9537 4111 9571
rect 5089 9537 5123 9571
rect 6009 9537 6043 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 7757 9537 7791 9571
rect 8125 9537 8159 9571
rect 8769 9537 8803 9571
rect 9137 9537 9171 9571
rect 9781 9537 9815 9571
rect 10149 9537 10183 9571
rect 1685 9401 1719 9435
rect 8585 9401 8619 9435
rect 9597 9401 9631 9435
rect 2697 9333 2731 9367
rect 6193 9333 6227 9367
rect 7573 9333 7607 9367
rect 1777 9129 1811 9163
rect 4261 9129 4295 9163
rect 5273 9129 5307 9163
rect 10241 9129 10275 9163
rect 2053 9061 2087 9095
rect 9873 9061 9907 9095
rect 1409 8925 1443 8959
rect 1961 8925 1995 8959
rect 2237 8925 2271 8959
rect 4445 8925 4479 8959
rect 5457 8925 5491 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 6736 8857 6770 8891
rect 9321 8857 9355 8891
rect 9597 8857 9631 8891
rect 10149 8857 10183 8891
rect 1593 8789 1627 8823
rect 6101 8789 6135 8823
rect 7849 8789 7883 8823
rect 8677 8789 8711 8823
rect 8953 8789 8987 8823
rect 7389 8585 7423 8619
rect 7665 8585 7699 8619
rect 8677 8585 8711 8619
rect 9873 8585 9907 8619
rect 10241 8585 10275 8619
rect 1593 8449 1627 8483
rect 7297 8449 7331 8483
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8769 8449 8803 8483
rect 10057 8449 10091 8483
rect 10149 8449 10183 8483
rect 6561 8381 6595 8415
rect 8217 8381 8251 8415
rect 8953 8381 8987 8415
rect 9505 8381 9539 8415
rect 1409 8245 1443 8279
rect 7113 8245 7147 8279
rect 9413 8245 9447 8279
rect 2513 8041 2547 8075
rect 9413 8041 9447 8075
rect 1593 7973 1627 8007
rect 8493 7973 8527 8007
rect 6101 7905 6135 7939
rect 8953 7905 8987 7939
rect 9137 7905 9171 7939
rect 9689 7905 9723 7939
rect 1777 7837 1811 7871
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 6368 7837 6402 7871
rect 7757 7837 7791 7871
rect 8677 7837 8711 7871
rect 9873 7837 9907 7871
rect 2053 7701 2087 7735
rect 7481 7701 7515 7735
rect 8401 7701 8435 7735
rect 10333 7701 10367 7735
rect 2789 7497 2823 7531
rect 7113 7497 7147 7531
rect 9873 7497 9907 7531
rect 9965 7497 9999 7531
rect 10241 7497 10275 7531
rect 5089 7429 5123 7463
rect 8024 7429 8058 7463
rect 1409 7361 1443 7395
rect 1961 7361 1995 7395
rect 2973 7361 3007 7395
rect 3249 7361 3283 7395
rect 3341 7361 3375 7395
rect 4997 7361 5031 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 10149 7361 10183 7395
rect 10425 7361 10459 7395
rect 2145 7293 2179 7327
rect 4077 7293 4111 7327
rect 6377 7293 6411 7327
rect 7757 7293 7791 7327
rect 9229 7293 9263 7327
rect 9413 7293 9447 7327
rect 1593 7225 1627 7259
rect 3433 7225 3467 7259
rect 1777 7157 1811 7191
rect 2697 7157 2731 7191
rect 3065 7157 3099 7191
rect 5733 7157 5767 7191
rect 6101 7157 6135 7191
rect 7021 7157 7055 7191
rect 7573 7157 7607 7191
rect 9137 7157 9171 7191
rect 2881 6953 2915 6987
rect 8585 6953 8619 6987
rect 10057 6953 10091 6987
rect 3801 6885 3835 6919
rect 9321 6885 9355 6919
rect 4077 6817 4111 6851
rect 6101 6817 6135 6851
rect 7665 6817 7699 6851
rect 8125 6817 8159 6851
rect 8401 6817 8435 6851
rect 8953 6817 8987 6851
rect 1501 6749 1535 6783
rect 1768 6749 1802 6783
rect 3157 6749 3191 6783
rect 3433 6749 3467 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 5089 6749 5123 6783
rect 5181 6749 5215 6783
rect 5365 6749 5399 6783
rect 5917 6749 5951 6783
rect 6653 6749 6687 6783
rect 7481 6749 7515 6783
rect 8309 6749 8343 6783
rect 8769 6749 8803 6783
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 9965 6749 9999 6783
rect 10425 6749 10459 6783
rect 6745 6681 6779 6715
rect 2973 6613 3007 6647
rect 3525 6613 3559 6647
rect 4721 6613 4755 6647
rect 4905 6613 4939 6647
rect 5825 6613 5859 6647
rect 6561 6613 6595 6647
rect 9689 6613 9723 6647
rect 10241 6613 10275 6647
rect 2053 6409 2087 6443
rect 4353 6409 4387 6443
rect 7113 6409 7147 6443
rect 9045 6409 9079 6443
rect 10333 6409 10367 6443
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 2493 6273 2527 6307
rect 4445 6273 4479 6307
rect 6377 6273 6411 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 9229 6273 9263 6307
rect 9597 6273 9631 6307
rect 9965 6273 9999 6307
rect 10517 6273 10551 6307
rect 3709 6205 3743 6239
rect 3893 6205 3927 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8309 6205 8343 6239
rect 8493 6205 8527 6239
rect 9689 6205 9723 6239
rect 1593 6137 1627 6171
rect 3617 6137 3651 6171
rect 6837 6137 6871 6171
rect 1777 6069 1811 6103
rect 5733 6069 5767 6103
rect 6469 6069 6503 6103
rect 8217 6069 8251 6103
rect 8677 6069 8711 6103
rect 9413 6069 9447 6103
rect 10057 6069 10091 6103
rect 3157 5865 3191 5899
rect 3525 5865 3559 5899
rect 4445 5865 4479 5899
rect 6561 5865 6595 5899
rect 7757 5865 7791 5899
rect 2881 5797 2915 5831
rect 7481 5797 7515 5831
rect 8677 5797 8711 5831
rect 9321 5797 9355 5831
rect 3801 5729 3835 5763
rect 7205 5729 7239 5763
rect 8033 5729 8067 5763
rect 8953 5729 8987 5763
rect 9689 5729 9723 5763
rect 9873 5729 9907 5763
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2237 5661 2271 5695
rect 2329 5661 2363 5695
rect 2605 5661 2639 5695
rect 3065 5661 3099 5695
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 4537 5661 4571 5695
rect 7113 5661 7147 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 8217 5661 8251 5695
rect 9137 5661 9171 5695
rect 2697 5593 2731 5627
rect 5273 5593 5307 5627
rect 1501 5525 1535 5559
rect 1777 5525 1811 5559
rect 2053 5525 2087 5559
rect 2421 5525 2455 5559
rect 5181 5525 5215 5559
rect 10333 5525 10367 5559
rect 1593 5321 1627 5355
rect 1869 5321 1903 5355
rect 2789 5321 2823 5355
rect 3525 5321 3559 5355
rect 5181 5321 5215 5355
rect 7665 5321 7699 5355
rect 9505 5321 9539 5355
rect 10241 5321 10275 5355
rect 4068 5253 4102 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 2329 5185 2363 5219
rect 3065 5185 3099 5219
rect 3801 5185 3835 5219
rect 5549 5185 5583 5219
rect 7573 5185 7607 5219
rect 8033 5185 8067 5219
rect 8125 5185 8159 5219
rect 8392 5185 8426 5219
rect 9597 5185 9631 5219
rect 10333 5185 10367 5219
rect 2145 5117 2179 5151
rect 2881 5117 2915 5151
rect 5733 5117 5767 5151
rect 6377 5117 6411 5151
rect 6561 5117 6595 5151
rect 7113 5117 7147 5151
rect 9781 5117 9815 5151
rect 10517 5049 10551 5083
rect 5917 4981 5951 5015
rect 6745 4981 6779 5015
rect 7849 4981 7883 5015
rect 1869 4777 1903 4811
rect 5457 4777 5491 4811
rect 7205 4777 7239 4811
rect 9597 4777 9631 4811
rect 9965 4777 9999 4811
rect 2881 4709 2915 4743
rect 3341 4709 3375 4743
rect 6561 4709 6595 4743
rect 8769 4709 8803 4743
rect 9689 4709 9723 4743
rect 2237 4641 2271 4675
rect 2973 4641 3007 4675
rect 3985 4641 4019 4675
rect 5825 4641 5859 4675
rect 6009 4641 6043 4675
rect 7389 4641 7423 4675
rect 1409 4573 1443 4607
rect 1685 4573 1719 4607
rect 2145 4573 2179 4607
rect 2421 4573 2455 4607
rect 3157 4573 3191 4607
rect 4252 4573 4286 4607
rect 5641 4573 5675 4607
rect 6469 4573 6503 4607
rect 6745 4573 6779 4607
rect 7021 4573 7055 4607
rect 7113 4573 7147 4607
rect 8953 4573 8987 4607
rect 9873 4573 9907 4607
rect 10149 4573 10183 4607
rect 10517 4573 10551 4607
rect 1501 4505 1535 4539
rect 7656 4505 7690 4539
rect 1961 4437 1995 4471
rect 5365 4437 5399 4471
rect 6837 4437 6871 4471
rect 10333 4437 10367 4471
rect 1593 4233 1627 4267
rect 2053 4233 2087 4267
rect 2421 4233 2455 4267
rect 5825 4233 5859 4267
rect 8677 4233 8711 4267
rect 9597 4165 9631 4199
rect 1501 4097 1535 4131
rect 1961 4097 1995 4131
rect 2237 4097 2271 4131
rect 2329 4097 2363 4131
rect 2781 4097 2815 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3617 4097 3651 4131
rect 3709 4097 3743 4131
rect 4169 4097 4203 4131
rect 4261 4097 4295 4131
rect 5365 4097 5399 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 7205 4097 7239 4131
rect 8953 4097 8987 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 10057 4097 10091 4131
rect 10333 4097 10367 4131
rect 2973 4029 3007 4063
rect 4445 4029 4479 4063
rect 5181 4029 5215 4063
rect 6377 4029 6411 4063
rect 7389 4029 7423 4063
rect 8125 4029 8159 4063
rect 2605 3961 2639 3995
rect 3433 3961 3467 3995
rect 9045 3961 9079 3995
rect 1777 3893 1811 3927
rect 3157 3893 3191 3927
rect 3893 3893 3927 3927
rect 3985 3893 4019 3927
rect 4905 3893 4939 3927
rect 7021 3893 7055 3927
rect 7849 3893 7883 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 10149 3893 10183 3927
rect 10517 3893 10551 3927
rect 2145 3689 2179 3723
rect 3893 3689 3927 3723
rect 8401 3689 8435 3723
rect 4997 3621 5031 3655
rect 6745 3621 6779 3655
rect 2697 3553 2731 3587
rect 2881 3553 2915 3587
rect 4445 3553 4479 3587
rect 5181 3553 5215 3587
rect 6193 3553 6227 3587
rect 7021 3553 7055 3587
rect 9045 3553 9079 3587
rect 10149 3553 10183 3587
rect 1869 3485 1903 3519
rect 2329 3485 2363 3519
rect 2421 3485 2455 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 8493 3485 8527 3519
rect 4537 3417 4571 3451
rect 6285 3417 6319 3451
rect 7288 3417 7322 3451
rect 9137 3417 9171 3451
rect 9689 3417 9723 3451
rect 9873 3417 9907 3451
rect 9965 3417 9999 3451
rect 2513 3349 2547 3383
rect 3341 3349 3375 3383
rect 3617 3349 3651 3383
rect 4169 3349 4203 3383
rect 5825 3349 5859 3383
rect 8585 3349 8619 3383
rect 3893 3145 3927 3179
rect 6009 3145 6043 3179
rect 8493 3145 8527 3179
rect 9321 3145 9355 3179
rect 1501 3077 1535 3111
rect 2053 3077 2087 3111
rect 2605 3077 2639 3111
rect 4896 3077 4930 3111
rect 6644 3077 6678 3111
rect 9229 3077 9263 3111
rect 4629 3009 4663 3043
rect 6377 3009 6411 3043
rect 8585 3009 8619 3043
rect 8769 3009 8803 3043
rect 9505 3009 9539 3043
rect 9781 3009 9815 3043
rect 10149 3009 10183 3043
rect 7941 2941 7975 2975
rect 7757 2873 7791 2907
rect 1593 2805 1627 2839
rect 2145 2805 2179 2839
rect 9597 2805 9631 2839
rect 10425 2805 10459 2839
rect 1593 2601 1627 2635
rect 3433 2601 3467 2635
rect 4997 2601 5031 2635
rect 5917 2601 5951 2635
rect 7573 2601 7607 2635
rect 5641 2533 5675 2567
rect 2973 2465 3007 2499
rect 3157 2465 3191 2499
rect 4353 2465 4387 2499
rect 4537 2465 4571 2499
rect 1777 2397 1811 2431
rect 2513 2397 2547 2431
rect 3893 2397 3927 2431
rect 5825 2397 5859 2431
rect 6101 2397 6135 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 10241 2397 10275 2431
rect 1961 2329 1995 2363
rect 2881 2329 2915 2363
rect 5181 2329 5215 2363
rect 6469 2329 6503 2363
rect 8493 2329 8527 2363
rect 9045 2329 9079 2363
rect 9781 2329 9815 2363
rect 2237 2261 2271 2295
rect 3985 2261 4019 2295
rect 5273 2261 5307 2295
rect 6561 2261 6595 2295
rect 7113 2261 7147 2295
rect 8033 2261 8067 2295
rect 9137 2261 9171 2295
rect 9873 2261 9907 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 4157 9707 4215 9713
rect 4157 9704 4169 9707
rect 3936 9676 4169 9704
rect 3936 9664 3942 9676
rect 4157 9673 4169 9676
rect 4203 9673 4215 9707
rect 4157 9667 4215 9673
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7984 9676 8217 9704
rect 7984 9664 7990 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 2409 9639 2467 9645
rect 2409 9636 2421 9639
rect 1912 9608 2421 9636
rect 1912 9596 1918 9608
rect 2409 9605 2421 9608
rect 2455 9605 2467 9639
rect 2409 9599 2467 9605
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 2924 9608 3433 9636
rect 2924 9596 2930 9608
rect 3421 9605 3433 9608
rect 3467 9605 3479 9639
rect 3421 9599 3479 9605
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 4948 9608 5457 9636
rect 4948 9596 4954 9608
rect 5445 9605 5457 9608
rect 5491 9605 5503 9639
rect 5445 9599 5503 9605
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6236 9608 6837 9636
rect 6236 9596 6242 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7469 9639 7527 9645
rect 7469 9636 7481 9639
rect 6972 9608 7481 9636
rect 6972 9596 6978 9608
rect 7469 9605 7481 9608
rect 7515 9605 7527 9639
rect 7469 9599 7527 9605
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8996 9608 9505 9636
rect 8996 9596 9002 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10505 9639 10563 9645
rect 10505 9636 10517 9639
rect 10008 9608 10517 9636
rect 10008 9596 10014 9608
rect 10505 9605 10517 9608
rect 10551 9605 10563 9639
rect 10505 9599 10563 9605
rect 1486 9528 1492 9580
rect 1544 9528 1550 9580
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 1728 9540 2053 9568
rect 1728 9528 1734 9540
rect 2041 9537 2053 9540
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2774 9568 2780 9580
rect 2547 9540 2780 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 4062 9528 4068 9580
rect 4120 9528 4126 9580
rect 5074 9528 5080 9580
rect 5132 9528 5138 9580
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9568 7159 9571
rect 7374 9568 7380 9580
rect 7147 9540 7380 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 842 9392 848 9444
rect 900 9432 906 9444
rect 1673 9435 1731 9441
rect 1673 9432 1685 9435
rect 900 9404 1685 9432
rect 900 9392 906 9404
rect 1673 9401 1685 9404
rect 1719 9401 1731 9435
rect 6012 9432 6040 9531
rect 6472 9500 6500 9531
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7834 9568 7840 9580
rect 7791 9540 7840 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8159 9540 8708 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8680 9500 8708 9540
rect 8754 9528 8760 9580
rect 8812 9528 8818 9580
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9769 9571 9827 9577
rect 9171 9540 9628 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9030 9500 9036 9512
rect 6472 9472 8616 9500
rect 8680 9472 9036 9500
rect 8588 9441 8616 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9600 9441 9628 9540
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 8573 9435 8631 9441
rect 6012 9404 8248 9432
rect 1673 9395 1731 9401
rect 8220 9376 8248 9404
rect 8573 9401 8585 9435
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 9585 9435 9643 9441
rect 9585 9401 9597 9435
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 2682 9324 2688 9376
rect 2740 9324 2746 9376
rect 6178 9324 6184 9376
rect 6236 9324 6242 9376
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 7926 9364 7932 9376
rect 7607 9336 7932 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9784 9364 9812 9531
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 9272 9336 9812 9364
rect 9272 9324 9278 9336
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1765 9163 1823 9169
rect 1765 9160 1777 9163
rect 1544 9132 1777 9160
rect 1544 9120 1550 9132
rect 1765 9129 1777 9132
rect 1811 9129 1823 9163
rect 1765 9123 1823 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4120 9132 4261 9160
rect 4120 9120 4126 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 5132 9132 5273 9160
rect 5132 9120 5138 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6236 9132 7512 9160
rect 6236 9120 6242 9132
rect 2041 9095 2099 9101
rect 2041 9061 2053 9095
rect 2087 9092 2099 9095
rect 7484 9092 7512 9132
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9364 9132 10241 9160
rect 9364 9120 9370 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 11054 9120 11060 9172
rect 11112 9120 11118 9172
rect 9214 9092 9220 9104
rect 2087 9064 6316 9092
rect 7484 9064 9220 9092
rect 2087 9061 2099 9064
rect 2041 9055 2099 9061
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1946 8916 1952 8968
rect 2004 8916 2010 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2958 8956 2964 8968
rect 2271 8928 2964 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 6288 8965 6316 9064
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 9861 9095 9919 9101
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 11072 9092 11100 9120
rect 9907 9064 11100 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 7984 8996 9168 9024
rect 7984 8984 7990 8996
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 5445 8959 5503 8965
rect 4479 8928 5396 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5368 8832 5396 8928
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 5460 8888 5488 8919
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6656 8928 7512 8956
rect 6656 8888 6684 8928
rect 5460 8860 6684 8888
rect 6724 8891 6782 8897
rect 6724 8857 6736 8891
rect 6770 8888 6782 8891
rect 7282 8888 7288 8900
rect 6770 8860 7288 8888
rect 6770 8857 6782 8860
rect 6724 8851 6782 8857
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 7484 8888 7512 8928
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7616 8928 8033 8956
rect 7616 8916 7622 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 9140 8965 9168 8996
rect 9232 8965 9260 9052
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8168 8928 8217 8956
rect 8168 8916 8174 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 7926 8888 7932 8900
rect 7484 8860 7932 8888
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 9309 8891 9367 8897
rect 9309 8888 9321 8891
rect 8036 8860 9321 8888
rect 8036 8832 8064 8860
rect 9309 8857 9321 8860
rect 9355 8857 9367 8891
rect 9309 8851 9367 8857
rect 9585 8891 9643 8897
rect 9585 8857 9597 8891
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 10137 8891 10195 8897
rect 10137 8857 10149 8891
rect 10183 8888 10195 8891
rect 10318 8888 10324 8900
rect 10183 8860 10324 8888
rect 10183 8857 10195 8860
rect 10137 8851 10195 8857
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1544 8792 1593 8820
rect 1544 8780 1550 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 5350 8780 5356 8832
rect 5408 8780 5414 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 7650 8820 7656 8832
rect 6135 8792 7656 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7834 8780 7840 8832
rect 7892 8780 7898 8832
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8904 8792 8953 8820
rect 8904 8780 8910 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9600 8820 9628 8851
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 9180 8792 9628 8820
rect 9180 8780 9186 8792
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 7377 8619 7435 8625
rect 2740 8576 2774 8616
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7558 8616 7564 8628
rect 7423 8588 7564 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7653 8619 7711 8625
rect 7653 8585 7665 8619
rect 7699 8616 7711 8619
rect 8110 8616 8116 8628
rect 7699 8588 8116 8616
rect 7699 8585 7711 8588
rect 7653 8579 7711 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8662 8576 8668 8628
rect 8720 8576 8726 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9088 8588 9873 8616
rect 9088 8576 9094 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 10192 8588 10241 8616
rect 10192 8576 10198 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 2746 8548 2774 8576
rect 2746 8520 9996 8548
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 7300 8489 7328 8520
rect 9968 8492 9996 8520
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7834 8480 7840 8492
rect 7607 8452 7840 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8412 6607 8415
rect 6822 8412 6828 8424
rect 6595 8384 6828 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 6822 8372 6828 8384
rect 6880 8412 6886 8424
rect 7576 8412 7604 8443
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 6880 8384 7604 8412
rect 8205 8415 8263 8421
rect 6880 8372 6886 8384
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8864 8412 8892 8440
rect 8251 8384 8892 8412
rect 8941 8415 8999 8421
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 7340 8316 8800 8344
rect 7340 8304 7346 8316
rect 1394 8236 1400 8288
rect 1452 8236 1458 8288
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 6972 8248 7113 8276
rect 6972 8236 6978 8248
rect 7101 8245 7113 8248
rect 7147 8245 7159 8279
rect 8772 8276 8800 8316
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 8956 8344 8984 8375
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9088 8384 9505 8412
rect 9088 8372 9094 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10152 8412 10180 8443
rect 9916 8384 10180 8412
rect 9916 8372 9922 8384
rect 10410 8344 10416 8356
rect 8904 8316 8984 8344
rect 9048 8316 10416 8344
rect 8904 8304 8910 8316
rect 9048 8276 9076 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 8772 8248 9076 8276
rect 7101 8239 7159 8245
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2498 8072 2504 8084
rect 2004 8044 2504 8072
rect 2004 8032 2010 8044
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 6454 8072 6460 8084
rect 6104 8044 6460 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 2682 8004 2688 8016
rect 1627 7976 2688 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 2682 7964 2688 7976
rect 2740 7964 2746 8016
rect 6104 7945 6132 8044
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 9398 8032 9404 8084
rect 9456 8032 9462 8084
rect 8481 8007 8539 8013
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 8527 7976 9168 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9030 7936 9036 7948
rect 8987 7908 9036 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 9140 7945 9168 7976
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 9416 7936 9444 8032
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9416 7908 9689 7936
rect 9125 7899 9183 7905
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 1872 7840 2237 7868
rect 1872 7744 1900 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 6356 7871 6414 7877
rect 6356 7837 6368 7871
rect 6402 7868 6414 7871
rect 6914 7868 6920 7880
rect 6402 7840 6920 7868
rect 6402 7837 6414 7840
rect 6356 7831 6414 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7484 7840 7757 7868
rect 7484 7744 7512 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 8662 7828 8668 7880
rect 8720 7828 8726 7880
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10226 7868 10232 7880
rect 9907 7840 10232 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 1854 7692 1860 7744
rect 1912 7692 1918 7744
rect 2038 7692 2044 7744
rect 2096 7692 2102 7744
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 6178 7732 6184 7744
rect 2556 7704 6184 7732
rect 2556 7692 2562 7704
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 7466 7692 7472 7744
rect 7524 7692 7530 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 8168 7704 8401 7732
rect 8168 7692 8174 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 8389 7695 8447 7701
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 9916 7704 10333 7732
rect 9916 7692 9922 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 1394 7488 1400 7540
rect 1452 7488 1458 7540
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2777 7531 2835 7537
rect 2004 7500 2268 7528
rect 2004 7488 2010 7500
rect 1412 7460 1440 7488
rect 1412 7432 1992 7460
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1964 7401 1992 7432
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 2240 7392 2268 7500
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 3050 7528 3056 7540
rect 2823 7500 3056 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7374 7528 7380 7540
rect 7147 7500 7380 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 9122 7528 9128 7540
rect 7484 7500 9128 7528
rect 5077 7463 5135 7469
rect 5077 7429 5089 7463
rect 5123 7460 5135 7463
rect 7484 7460 7512 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 9858 7488 9864 7540
rect 9916 7488 9922 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 5123 7432 7512 7460
rect 8012 7463 8070 7469
rect 5123 7429 5135 7432
rect 5077 7423 5135 7429
rect 8012 7429 8024 7463
rect 8058 7460 8070 7463
rect 8110 7460 8116 7472
rect 8058 7432 8116 7460
rect 8058 7429 8070 7432
rect 8012 7423 8070 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 9968 7460 9996 7491
rect 10226 7488 10232 7540
rect 10284 7488 10290 7540
rect 9968 7432 10456 7460
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2240 7364 2973 7392
rect 1949 7355 2007 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4396 7364 4997 7392
rect 4396 7352 4402 7364
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5592 7364 5917 7392
rect 5592 7352 5598 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6043 7364 6316 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2590 7324 2596 7336
rect 2179 7296 2596 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2746 7296 4016 7324
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2746 7256 2774 7296
rect 1627 7228 2774 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2866 7216 2872 7268
rect 2924 7256 2930 7268
rect 3421 7259 3479 7265
rect 3421 7256 3433 7259
rect 2924 7228 3433 7256
rect 2924 7216 2930 7228
rect 3421 7225 3433 7228
rect 3467 7225 3479 7259
rect 3988 7256 4016 7296
rect 4062 7284 4068 7336
rect 4120 7284 4126 7336
rect 4154 7256 4160 7268
rect 3988 7228 4160 7256
rect 3421 7219 3479 7225
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 2406 7188 2412 7200
rect 1811 7160 2412 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2498 7148 2504 7200
rect 2556 7188 2562 7200
rect 2685 7191 2743 7197
rect 2685 7188 2697 7191
rect 2556 7160 2697 7188
rect 2556 7148 2562 7160
rect 2685 7157 2697 7160
rect 2731 7157 2743 7191
rect 2685 7151 2743 7157
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 4982 7188 4988 7200
rect 3099 7160 4988 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5718 7148 5724 7200
rect 5776 7148 5782 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6089 7191 6147 7197
rect 6089 7188 6101 7191
rect 5868 7160 6101 7188
rect 5868 7148 5874 7160
rect 6089 7157 6101 7160
rect 6135 7157 6147 7191
rect 6288 7188 6316 7364
rect 6454 7352 6460 7404
rect 6512 7352 6518 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7374 7392 7380 7404
rect 7331 7364 7380 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 8294 7392 8300 7404
rect 7524 7364 8300 7392
rect 7524 7352 7530 7364
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9140 7364 10149 7392
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6472 7324 6500 7352
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 6472 7296 7757 7324
rect 6365 7287 6423 7293
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 6380 7256 6408 7287
rect 6380 7228 7788 7256
rect 6822 7188 6828 7200
rect 6288 7160 6828 7188
rect 6089 7151 6147 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 6972 7160 7021 7188
rect 6972 7148 6978 7160
rect 7009 7157 7021 7160
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 7760 7188 7788 7228
rect 9140 7197 9168 7364
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 10226 7392 10232 7404
rect 10183 7364 10232 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10428 7401 10456 7432
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 10042 7324 10048 7336
rect 9447 7296 10048 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 7760 7160 9137 7188
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 2648 6956 2881 6984
rect 2648 6944 2654 6956
rect 2869 6953 2881 6956
rect 2915 6953 2927 6987
rect 2869 6947 2927 6953
rect 8573 6987 8631 6993
rect 8573 6953 8585 6987
rect 8619 6984 8631 6987
rect 8662 6984 8668 6996
rect 8619 6956 8668 6984
rect 8619 6953 8631 6956
rect 8573 6947 8631 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 10042 6944 10048 6996
rect 10100 6944 10106 6996
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 3326 6916 3332 6928
rect 2832 6888 3332 6916
rect 2832 6876 2838 6888
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 3786 6876 3792 6928
rect 3844 6876 3850 6928
rect 9214 6916 9220 6928
rect 3988 6888 4200 6916
rect 3988 6848 4016 6888
rect 2746 6820 4016 6848
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1756 6783 1814 6789
rect 1756 6749 1768 6783
rect 1802 6780 1814 6783
rect 2746 6780 2774 6820
rect 4062 6808 4068 6860
rect 4120 6808 4126 6860
rect 4172 6848 4200 6888
rect 5644 6888 6224 6916
rect 5644 6848 5672 6888
rect 4172 6820 5672 6848
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5776 6820 6101 6848
rect 5776 6808 5782 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6196 6848 6224 6888
rect 8312 6888 9220 6916
rect 6196 6820 6960 6848
rect 6089 6811 6147 6817
rect 6932 6792 6960 6820
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7616 6820 7665 6848
rect 7616 6808 7622 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8312 6848 8340 6888
rect 9214 6876 9220 6888
rect 9272 6916 9278 6928
rect 9309 6919 9367 6925
rect 9309 6916 9321 6919
rect 9272 6888 9321 6916
rect 9272 6876 9278 6888
rect 9309 6885 9321 6888
rect 9355 6885 9367 6919
rect 9309 6879 9367 6885
rect 8159 6820 8340 6848
rect 8389 6851 8447 6857
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8389 6817 8401 6851
rect 8435 6848 8447 6851
rect 8846 6848 8852 6860
rect 8435 6820 8852 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 10594 6848 10600 6860
rect 10428 6820 10600 6848
rect 1802 6752 2774 6780
rect 1802 6749 1814 6752
rect 1756 6743 1814 6749
rect 1504 6712 1532 6743
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3384 6752 3433 6780
rect 3384 6740 3390 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3421 6743 3479 6749
rect 3528 6752 3985 6780
rect 2130 6712 2136 6724
rect 1504 6684 2136 6712
rect 2130 6672 2136 6684
rect 2188 6672 2194 6724
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3528 6712 3556 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 3108 6684 3556 6712
rect 3108 6672 3114 6684
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 4264 6712 4292 6743
rect 5074 6740 5080 6792
rect 5132 6740 5138 6792
rect 5166 6740 5172 6792
rect 5224 6740 5230 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5810 6780 5816 6792
rect 5399 6752 5816 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 3844 6684 4292 6712
rect 5920 6712 5948 6743
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 6236 6752 6653 6780
rect 6236 6740 6242 6752
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 5920 6684 6745 6712
rect 3844 6672 3850 6684
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 2958 6604 2964 6656
rect 3016 6604 3022 6656
rect 3513 6647 3571 6653
rect 3513 6613 3525 6647
rect 3559 6644 3571 6647
rect 4246 6644 4252 6656
rect 3559 6616 4252 6644
rect 3559 6613 3571 6616
rect 3513 6607 3571 6613
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4396 6616 4721 6644
rect 4396 6604 4402 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5626 6644 5632 6656
rect 4939 6616 5632 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 5859 6616 6561 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6549 6613 6561 6616
rect 6595 6644 6607 6647
rect 7484 6644 7512 6743
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8352 6752 8769 6780
rect 8352 6740 8358 6752
rect 8757 6749 8769 6752
rect 8803 6780 8815 6783
rect 9125 6783 9183 6789
rect 8803 6752 9076 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 9048 6712 9076 6752
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9171 6752 9720 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9214 6712 9220 6724
rect 9048 6684 9220 6712
rect 9214 6672 9220 6684
rect 9272 6672 9278 6724
rect 9692 6653 9720 6752
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 10226 6780 10232 6792
rect 9999 6752 10232 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10428 6789 10456 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 6595 6616 7512 6644
rect 9677 6647 9735 6653
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 9677 6613 9689 6647
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 10410 6644 10416 6656
rect 10275 6616 10416 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 1946 6440 1952 6452
rect 1688 6412 1952 6440
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1688 6313 1716 6412
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2087 6412 3556 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 3528 6372 3556 6412
rect 4338 6400 4344 6452
rect 4396 6400 4402 6452
rect 5166 6400 5172 6452
rect 5224 6400 5230 6452
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9858 6440 9864 6452
rect 9079 6412 9864 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 5184 6372 5212 6400
rect 3528 6344 5212 6372
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1544 6276 1685 6304
rect 1544 6264 1550 6276
rect 1673 6273 1685 6276
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1946 6264 1952 6316
rect 2004 6264 2010 6316
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2188 6276 2237 6304
rect 2188 6264 2194 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2481 6307 2539 6313
rect 2372 6302 2452 6304
rect 2481 6302 2493 6307
rect 2372 6276 2493 6302
rect 2372 6264 2378 6276
rect 2424 6274 2493 6276
rect 2481 6273 2493 6274
rect 2527 6273 2539 6307
rect 2481 6267 2539 6273
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4212 6276 4445 6304
rect 4212 6264 4218 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 7009 6307 7067 6313
rect 6411 6276 6776 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 1854 6236 1860 6248
rect 1596 6208 1860 6236
rect 1596 6177 1624 6208
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 3786 6236 3792 6248
rect 3743 6208 3792 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 3970 6236 3976 6248
rect 3927 6208 3976 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6137 1639 6171
rect 1581 6131 1639 6137
rect 1780 6140 2268 6168
rect 1780 6109 1808 6140
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6069 1823 6103
rect 2240 6100 2268 6140
rect 3602 6128 3608 6180
rect 3660 6128 3666 6180
rect 3878 6100 3884 6112
rect 2240 6072 3884 6100
rect 1765 6063 1823 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 5258 6060 5264 6112
rect 5316 6100 5322 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5316 6072 5733 6100
rect 5316 6060 5322 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 6236 6072 6469 6100
rect 6236 6060 6242 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6748 6100 6776 6276
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7116 6304 7144 6403
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10192 6412 10333 6440
rect 10192 6400 10198 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 9600 6344 10456 6372
rect 7055 6276 7144 6304
rect 7285 6307 7343 6313
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 8938 6304 8944 6316
rect 7285 6267 7343 6273
rect 8680 6276 8944 6304
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7300 6236 7328 6267
rect 7466 6236 7472 6248
rect 6972 6208 7472 6236
rect 6972 6196 6978 6208
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7558 6196 7564 6248
rect 7616 6196 7622 6248
rect 7742 6196 7748 6248
rect 7800 6196 7806 6248
rect 8294 6196 8300 6248
rect 8352 6196 8358 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 6825 6171 6883 6177
rect 6825 6137 6837 6171
rect 6871 6168 6883 6171
rect 8496 6168 8524 6199
rect 6871 6140 8524 6168
rect 6871 6137 6883 6140
rect 6825 6131 6883 6137
rect 7374 6100 7380 6112
rect 6748 6072 7380 6100
rect 6457 6063 6515 6069
rect 7374 6060 7380 6072
rect 7432 6100 7438 6112
rect 7834 6100 7840 6112
rect 7432 6072 7840 6100
rect 7432 6060 7438 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8680 6109 8708 6276
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9600 6313 9628 6344
rect 10428 6316 10456 6344
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10318 6304 10324 6316
rect 10008 6276 10324 6304
rect 10008 6264 10014 6276
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10410 6264 10416 6316
rect 10468 6264 10474 6316
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 11054 6304 11060 6316
rect 10551 6276 11060 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 8754 6196 8760 6248
rect 8812 6196 8818 6248
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9456 6208 9689 6236
rect 9456 6196 9462 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 8251 6072 8677 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 8772 6100 8800 6196
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 8772 6072 9413 6100
rect 8665 6063 8723 6069
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 10042 6060 10048 6112
rect 10100 6060 10106 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1486 5856 1492 5908
rect 1544 5856 1550 5908
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 2406 5896 2412 5908
rect 1636 5868 2412 5896
rect 1636 5856 1642 5868
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2590 5856 2596 5908
rect 2648 5856 2654 5908
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 3108 5868 3157 5896
rect 3108 5856 3114 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3513 5899 3571 5905
rect 3145 5859 3203 5865
rect 3252 5868 3464 5896
rect 1504 5828 1532 5856
rect 2498 5828 2504 5840
rect 1504 5800 2504 5828
rect 2498 5788 2504 5800
rect 2556 5788 2562 5840
rect 2608 5760 2636 5856
rect 2774 5788 2780 5840
rect 2832 5788 2838 5840
rect 2869 5831 2927 5837
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 3252 5828 3280 5868
rect 2915 5800 3280 5828
rect 3436 5828 3464 5868
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3970 5896 3976 5908
rect 3559 5868 3976 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4706 5896 4712 5908
rect 4479 5868 4712 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6512 5868 6561 5896
rect 6512 5856 6518 5868
rect 6549 5865 6561 5868
rect 6595 5896 6607 5899
rect 6822 5896 6828 5908
rect 6595 5868 6828 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7742 5856 7748 5908
rect 7800 5856 7806 5908
rect 10042 5856 10048 5908
rect 10100 5856 10106 5908
rect 5092 5828 5120 5856
rect 3436 5800 5120 5828
rect 7469 5831 7527 5837
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 8294 5828 8300 5840
rect 7515 5800 8300 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 8294 5788 8300 5800
rect 8352 5828 8358 5840
rect 8665 5831 8723 5837
rect 8352 5800 8616 5828
rect 8352 5788 8358 5800
rect 1964 5732 2636 5760
rect 2792 5760 2820 5788
rect 3602 5760 3608 5772
rect 2792 5732 3096 5760
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 1964 5701 1992 5732
rect 2332 5701 2360 5732
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2240 5624 2268 5655
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2464 5664 2605 5692
rect 2464 5652 2470 5664
rect 2593 5661 2605 5664
rect 2639 5692 2651 5695
rect 2774 5692 2780 5704
rect 2639 5664 2780 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3068 5701 3096 5732
rect 3344 5732 3608 5760
rect 3344 5701 3372 5732
rect 3602 5720 3608 5732
rect 3660 5760 3666 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3660 5732 3801 5760
rect 3660 5720 3666 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 7193 5763 7251 5769
rect 4120 5732 7144 5760
rect 4120 5720 4126 5732
rect 7116 5701 7144 5732
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 7558 5760 7564 5772
rect 7239 5732 7564 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 7558 5720 7564 5732
rect 7616 5760 7622 5772
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7616 5732 8033 5760
rect 7616 5720 7622 5732
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8588 5760 8616 5800
rect 8665 5797 8677 5831
rect 8711 5828 8723 5831
rect 9309 5831 9367 5837
rect 9309 5828 9321 5831
rect 8711 5800 9321 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 9309 5797 9321 5800
rect 9355 5797 9367 5831
rect 9309 5791 9367 5797
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8588 5732 8953 5760
rect 8021 5723 8079 5729
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 9324 5760 9352 5791
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9324 5732 9689 5760
rect 8941 5723 8999 5729
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5760 9919 5763
rect 10060 5760 10088 5856
rect 9907 5732 10088 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3329 5695 3387 5701
rect 3099 5664 3280 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 1780 5596 2268 5624
rect 2685 5627 2743 5633
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 1780 5565 1808 5596
rect 2685 5593 2697 5627
rect 2731 5624 2743 5627
rect 3252 5624 3280 5664
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 3375 5664 3433 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3421 5661 3433 5664
rect 3467 5661 3479 5695
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3421 5655 3479 5661
rect 3988 5664 4537 5692
rect 3988 5636 4016 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 3970 5624 3976 5636
rect 2731 5596 3188 5624
rect 3252 5596 3976 5624
rect 2731 5593 2743 5596
rect 2685 5587 2743 5593
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 1765 5519 1823 5525
rect 2038 5516 2044 5568
rect 2096 5516 2102 5568
rect 2406 5516 2412 5568
rect 2464 5516 2470 5568
rect 3160 5556 3188 5596
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 5258 5624 5264 5636
rect 4396 5596 5264 5624
rect 4396 5584 4402 5596
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 7392 5624 7420 5655
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7524 5664 7665 5692
rect 7524 5652 7530 5664
rect 7653 5661 7665 5664
rect 7699 5692 7711 5695
rect 7699 5664 7788 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7760 5636 7788 5664
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 8168 5664 8217 5692
rect 8168 5652 8174 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 7392 5596 7512 5624
rect 4982 5556 4988 5568
rect 3160 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 7484 5556 7512 5596
rect 7742 5584 7748 5636
rect 7800 5584 7806 5636
rect 7944 5556 7972 5652
rect 10226 5556 10232 5568
rect 7484 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10318 5516 10324 5568
rect 10376 5516 10382 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1670 5352 1676 5364
rect 1627 5324 1676 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1857 5355 1915 5361
rect 1857 5352 1869 5355
rect 1820 5324 1869 5352
rect 1820 5312 1826 5324
rect 1857 5321 1869 5324
rect 1903 5321 1915 5355
rect 1857 5315 1915 5321
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 2823 5324 3525 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 3513 5321 3525 5324
rect 3559 5352 3571 5355
rect 3786 5352 3792 5364
rect 3559 5324 3792 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 4028 5324 5181 5352
rect 4028 5312 4034 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 5169 5315 5227 5321
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 8110 5352 8116 5364
rect 7699 5324 8116 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9950 5352 9956 5364
rect 9539 5324 9956 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10318 5352 10324 5364
rect 10275 5324 10324 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10502 5312 10508 5364
rect 10560 5312 10566 5364
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 4056 5287 4114 5293
rect 2096 5256 2774 5284
rect 2096 5244 2102 5256
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2406 5216 2412 5228
rect 2363 5188 2412 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2746 5216 2774 5256
rect 4056 5253 4068 5287
rect 4102 5284 4114 5287
rect 4706 5284 4712 5296
rect 4102 5256 4712 5284
rect 4102 5253 4114 5256
rect 4056 5247 4114 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 7374 5284 7380 5296
rect 6972 5256 7380 5284
rect 6972 5244 6978 5256
rect 7374 5244 7380 5256
rect 7432 5284 7438 5296
rect 7432 5256 8156 5284
rect 7432 5244 7438 5256
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 2746 5188 3065 5216
rect 3053 5185 3065 5188
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3786 5216 3792 5228
rect 3292 5188 3792 5216
rect 3292 5176 3298 5188
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 6178 5216 6184 5228
rect 5583 5188 6184 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7926 5216 7932 5228
rect 7607 5188 7932 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 8128 5225 8156 5256
rect 8220 5256 9260 5284
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2133 5151 2191 5157
rect 2133 5148 2145 5151
rect 1912 5120 2145 5148
rect 1912 5108 1918 5120
rect 2133 5117 2145 5120
rect 2179 5117 2191 5151
rect 2133 5111 2191 5117
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 2915 5120 3096 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3068 5024 3096 5120
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5684 5120 5733 5148
rect 5684 5108 5690 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5721 5111 5779 5117
rect 5920 5120 6377 5148
rect 3050 4972 3056 5024
rect 3108 4972 3114 5024
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 5920 5021 5948 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 6914 5148 6920 5160
rect 6595 5120 6920 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 7116 5080 7144 5111
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8220 5148 8248 5256
rect 8380 5219 8438 5225
rect 8380 5185 8392 5219
rect 8426 5216 8438 5219
rect 8938 5216 8944 5228
rect 8426 5188 8944 5216
rect 8426 5185 8438 5188
rect 8380 5179 8438 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 7892 5120 8248 5148
rect 7892 5108 7898 5120
rect 9122 5108 9128 5160
rect 9180 5108 9186 5160
rect 6512 5052 7144 5080
rect 6512 5040 6518 5052
rect 5905 5015 5963 5021
rect 5905 5012 5917 5015
rect 5776 4984 5917 5012
rect 5776 4972 5782 4984
rect 5905 4981 5917 4984
rect 5951 4981 5963 5015
rect 5905 4975 5963 4981
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6604 4984 6745 5012
rect 6604 4972 6610 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 6733 4975 6791 4981
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 9140 5012 9168 5108
rect 9232 5080 9260 5256
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 9456 5188 9597 5216
rect 9456 5176 9462 5188
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10520 5216 10548 5312
rect 10367 5188 10548 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 9769 5151 9827 5157
rect 9769 5117 9781 5151
rect 9815 5148 9827 5151
rect 9950 5148 9956 5160
rect 9815 5120 9956 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 9232 5052 10517 5080
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 10505 5043 10563 5049
rect 7883 4984 9168 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1670 4768 1676 4820
rect 1728 4768 1734 4820
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 1946 4808 1952 4820
rect 1903 4780 1952 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3234 4808 3240 4820
rect 2832 4780 3240 4808
rect 2832 4768 2838 4780
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 4246 4808 4252 4820
rect 3344 4780 4252 4808
rect 1688 4672 1716 4768
rect 3344 4749 3372 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5534 4808 5540 4820
rect 5491 4780 5540 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 6454 4808 6460 4820
rect 5828 4780 6460 4808
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 3329 4743 3387 4749
rect 3329 4740 3341 4743
rect 2915 4712 3341 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 3329 4709 3341 4712
rect 3375 4709 3387 4743
rect 3329 4703 3387 4709
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 1412 4644 1716 4672
rect 1872 4644 2237 4672
rect 1412 4613 1440 4644
rect 1872 4616 1900 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2225 4635 2283 4641
rect 2332 4644 2973 4672
rect 2332 4616 2360 4644
rect 2961 4641 2973 4644
rect 3007 4672 3019 4675
rect 3050 4672 3056 4684
rect 3007 4644 3056 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 5828 4681 5856 4780
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6972 4780 7205 4808
rect 6972 4768 6978 4780
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 7193 4771 7251 4777
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8076 4780 8892 4808
rect 8076 4768 8082 4780
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 6012 4712 6561 4740
rect 6012 4681 6040 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4709 8815 4743
rect 8864 4740 8892 4780
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 8996 4780 9597 4808
rect 8996 4768 9002 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 9950 4768 9956 4820
rect 10008 4768 10014 4820
rect 10042 4768 10048 4820
rect 10100 4768 10106 4820
rect 9677 4743 9735 4749
rect 9677 4740 9689 4743
rect 8864 4712 9689 4740
rect 8757 4703 8815 4709
rect 9677 4709 9689 4712
rect 9723 4709 9735 4743
rect 9677 4703 9735 4709
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3844 4644 3985 4672
rect 3844 4632 3850 4644
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 5813 4675 5871 4681
rect 3973 4635 4031 4641
rect 5368 4644 5764 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 2130 4564 2136 4616
rect 2188 4564 2194 4616
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2406 4564 2412 4616
rect 2464 4564 2470 4616
rect 3145 4607 3203 4613
rect 3145 4598 3157 4607
rect 2884 4573 3157 4598
rect 3191 4573 3203 4607
rect 2884 4570 3203 4573
rect 1489 4539 1547 4545
rect 1489 4505 1501 4539
rect 1535 4536 1547 4539
rect 2498 4536 2504 4548
rect 1535 4508 2504 4536
rect 1535 4505 1547 4508
rect 1489 4499 1547 4505
rect 2498 4496 2504 4508
rect 2556 4496 2562 4548
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 2884 4468 2912 4570
rect 3145 4567 3203 4570
rect 4240 4607 4298 4613
rect 4240 4573 4252 4607
rect 4286 4604 4298 4607
rect 5166 4604 5172 4616
rect 4286 4576 5172 4604
rect 4286 4573 4298 4576
rect 4240 4567 4298 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 1995 4440 2912 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5368 4477 5396 4644
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5736 4604 5764 4644
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 6104 4644 7144 4672
rect 6104 4604 6132 4644
rect 5736 4576 6132 4604
rect 5629 4567 5687 4573
rect 5644 4536 5672 4567
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6236 4576 6469 4604
rect 6236 4564 6242 4576
rect 6457 4573 6469 4576
rect 6503 4604 6515 4607
rect 6546 4604 6552 4616
rect 6503 4576 6552 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 7116 4613 7144 4644
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7024 4536 7052 4567
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 8772 4604 8800 4703
rect 10060 4672 10088 4768
rect 10060 4644 10548 4672
rect 10520 4613 10548 4644
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 7984 4576 8953 4604
rect 7984 4564 7990 4576
rect 8941 4573 8953 4576
rect 8987 4604 8999 4607
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 8987 4576 9873 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4604 10195 4607
rect 10505 4607 10563 4613
rect 10183 4576 10364 4604
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 7466 4536 7472 4548
rect 5644 4508 6960 4536
rect 7024 4508 7472 4536
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5224 4440 5365 4468
rect 5224 4428 5230 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6604 4440 6837 4468
rect 6604 4428 6610 4440
rect 6825 4437 6837 4440
rect 6871 4437 6883 4471
rect 6932 4468 6960 4508
rect 7466 4496 7472 4508
rect 7524 4496 7530 4548
rect 7644 4539 7702 4545
rect 7644 4505 7656 4539
rect 7690 4536 7702 4539
rect 8662 4536 8668 4548
rect 7690 4508 8668 4536
rect 7690 4505 7702 4508
rect 7644 4499 7702 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 7742 4468 7748 4480
rect 6932 4440 7748 4468
rect 6825 4431 6883 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 10336 4477 10364 4576
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10321 4471 10379 4477
rect 10321 4437 10333 4471
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1581 4267 1639 4273
rect 1581 4233 1593 4267
rect 1627 4264 1639 4267
rect 1854 4264 1860 4276
rect 1627 4236 1860 4264
rect 1627 4233 1639 4236
rect 1581 4227 1639 4233
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 1946 4224 1952 4276
rect 2004 4224 2010 4276
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 2130 4264 2136 4276
rect 2087 4236 2136 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2409 4267 2467 4273
rect 2409 4264 2421 4267
rect 2372 4236 2421 4264
rect 2372 4224 2378 4236
rect 2409 4233 2421 4236
rect 2455 4233 2467 4267
rect 2409 4227 2467 4233
rect 2792 4236 3004 4264
rect 1762 4156 1768 4208
rect 1820 4156 1826 4208
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1780 4128 1808 4156
rect 1964 4137 1992 4224
rect 2792 4196 2820 4236
rect 2240 4168 2820 4196
rect 2976 4196 3004 4236
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 5813 4267 5871 4273
rect 5813 4264 5825 4267
rect 5776 4236 5825 4264
rect 5776 4224 5782 4236
rect 5813 4233 5825 4236
rect 5859 4233 5871 4267
rect 5813 4227 5871 4233
rect 8662 4224 8668 4276
rect 8720 4224 8726 4276
rect 10318 4224 10324 4276
rect 10376 4224 10382 4276
rect 10502 4224 10508 4276
rect 10560 4224 10566 4276
rect 3970 4196 3976 4208
rect 2976 4168 3976 4196
rect 2240 4137 2268 4168
rect 1535 4100 1808 4128
rect 1949 4131 2007 4137
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4097 2283 4131
rect 2225 4091 2283 4097
rect 2317 4131 2375 4137
rect 2769 4134 2827 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2608 4131 2827 4134
rect 2608 4128 2781 4131
rect 2363 4106 2781 4128
rect 2363 4100 2636 4106
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2769 4097 2781 4106
rect 2815 4097 2827 4131
rect 2769 4091 2827 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 2976 4128 3004 4168
rect 2915 4100 3004 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 1412 3992 1440 4088
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 2332 4060 2360 4091
rect 3142 4088 3148 4140
rect 3200 4088 3206 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3620 4137 3648 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 9585 4199 9643 4205
rect 9585 4165 9597 4199
rect 9631 4196 9643 4199
rect 9858 4196 9864 4208
rect 9631 4168 9864 4196
rect 9631 4165 9643 4168
rect 9585 4159 9643 4165
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 10336 4196 10364 4224
rect 10060 4168 10364 4196
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 1912 4032 2360 4060
rect 2792 4032 2973 4060
rect 1912 4020 1918 4032
rect 2593 3995 2651 4001
rect 2593 3992 2605 3995
rect 1412 3964 2605 3992
rect 2593 3961 2605 3964
rect 2639 3961 2651 3995
rect 2593 3955 2651 3961
rect 1762 3884 1768 3936
rect 1820 3884 1826 3936
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 2792 3924 2820 4032
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 2961 4023 3019 4029
rect 3160 3992 3188 4088
rect 3421 3995 3479 4001
rect 3421 3992 3433 3995
rect 3160 3964 3433 3992
rect 3421 3961 3433 3964
rect 3467 3961 3479 3995
rect 3712 3992 3740 4091
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 4120 4100 4169 4128
rect 4120 4088 4126 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 4580 4100 5365 4128
rect 4580 4088 4586 4100
rect 5353 4097 5365 4100
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5500 4100 6009 4128
rect 5500 4088 5506 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6135 4100 7205 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 8938 4088 8944 4140
rect 8996 4088 9002 4140
rect 10060 4137 10088 4168
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9263 4100 9321 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4128 10379 4131
rect 10520 4128 10548 4224
rect 10367 4100 10548 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 4430 4020 4436 4072
rect 4488 4020 4494 4072
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4948 4032 5181 4060
rect 4948 4020 4954 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 6362 4020 6368 4072
rect 6420 4020 6426 4072
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 7466 4060 7472 4072
rect 7423 4032 7472 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 9232 4060 9260 4091
rect 8168 4032 9260 4060
rect 8168 4020 8174 4032
rect 3712 3964 5212 3992
rect 3421 3955 3479 3961
rect 2464 3896 2820 3924
rect 2464 3884 2470 3896
rect 3142 3884 3148 3936
rect 3200 3884 3206 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 3881 3927 3939 3933
rect 3881 3924 3893 3927
rect 3752 3896 3893 3924
rect 3752 3884 3758 3896
rect 3881 3893 3893 3896
rect 3927 3893 3939 3927
rect 3881 3887 3939 3893
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5074 3924 5080 3936
rect 4939 3896 5080 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5184 3924 5212 3964
rect 6178 3952 6184 4004
rect 6236 3992 6242 4004
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 6236 3964 9045 3992
rect 6236 3952 6242 3964
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 6638 3924 6644 3936
rect 5184 3896 6644 3924
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6880 3896 7021 3924
rect 6880 3884 6886 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7009 3887 7067 3893
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 8662 3924 8668 3936
rect 7883 3896 8668 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 9398 3884 9404 3936
rect 9456 3884 9462 3936
rect 10134 3884 10140 3936
rect 10192 3884 10198 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10284 3896 10517 3924
rect 10284 3884 10290 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2590 3720 2596 3732
rect 2179 3692 2596 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4430 3720 4436 3732
rect 3927 3692 4436 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 6178 3720 6184 3732
rect 4540 3692 6184 3720
rect 4540 3652 4568 3692
rect 6178 3680 6184 3692
rect 6236 3680 6242 3732
rect 7374 3720 7380 3732
rect 6288 3692 6776 3720
rect 3436 3624 4568 3652
rect 4985 3655 5043 3661
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 2685 3587 2743 3593
rect 2685 3584 2697 3587
rect 2556 3556 2697 3584
rect 2556 3544 2562 3556
rect 2685 3553 2697 3556
rect 2731 3553 2743 3587
rect 2685 3547 2743 3553
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2832 3556 2881 3584
rect 2832 3544 2838 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2314 3516 2320 3528
rect 1903 3488 2320 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 3436 3525 3464 3624
rect 4985 3621 4997 3655
rect 5031 3652 5043 3655
rect 6288 3652 6316 3692
rect 6748 3661 6776 3692
rect 7024 3692 7380 3720
rect 5031 3624 6316 3652
rect 6733 3655 6791 3661
rect 5031 3621 5043 3624
rect 4985 3615 5043 3621
rect 6733 3621 6745 3655
rect 6779 3652 6791 3655
rect 6914 3652 6920 3664
rect 6779 3624 6920 3652
rect 6779 3621 6791 3624
rect 6733 3615 6791 3621
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4433 3587 4491 3593
rect 3752 3556 3832 3584
rect 3752 3544 3758 3556
rect 3804 3525 3832 3556
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 5074 3584 5080 3596
rect 4479 3556 5080 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 7024 3593 7052 3692
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 8168 3692 8401 3720
rect 8168 3680 8174 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 8389 3683 8447 3689
rect 8662 3680 8668 3732
rect 8720 3680 8726 3732
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6512 3556 7021 3584
rect 6512 3544 6518 3556
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 8680 3584 8708 3680
rect 8846 3584 8852 3596
rect 8680 3556 8852 3584
rect 7009 3547 7067 3553
rect 8846 3544 8852 3556
rect 8904 3584 8910 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8904 3556 9045 3584
rect 8904 3544 8910 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9033 3547 9091 3553
rect 9692 3556 10149 3584
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 2424 3448 2452 3479
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 8478 3476 8484 3528
rect 8536 3476 8542 3528
rect 4430 3448 4436 3460
rect 2424 3420 4436 3448
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 4525 3451 4583 3457
rect 4525 3417 4537 3451
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 3602 3340 3608 3392
rect 3660 3340 3666 3392
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4540 3380 4568 3411
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 6273 3451 6331 3457
rect 4672 3420 6040 3448
rect 4672 3408 4678 3420
rect 4203 3352 4568 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 5813 3383 5871 3389
rect 5813 3380 5825 3383
rect 5408 3352 5825 3380
rect 5408 3340 5414 3352
rect 5813 3349 5825 3352
rect 5859 3349 5871 3383
rect 6012 3380 6040 3420
rect 6273 3417 6285 3451
rect 6319 3448 6331 3451
rect 6546 3448 6552 3460
rect 6319 3420 6552 3448
rect 6319 3417 6331 3420
rect 6273 3411 6331 3417
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 7276 3451 7334 3457
rect 7276 3417 7288 3451
rect 7322 3448 7334 3451
rect 7834 3448 7840 3460
rect 7322 3420 7840 3448
rect 7322 3417 7334 3420
rect 7276 3411 7334 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 9125 3451 9183 3457
rect 8496 3420 8800 3448
rect 8496 3380 8524 3420
rect 6012 3352 8524 3380
rect 8573 3383 8631 3389
rect 5813 3343 5871 3349
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8662 3380 8668 3392
rect 8619 3352 8668 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 8772 3380 8800 3420
rect 9125 3417 9137 3451
rect 9171 3448 9183 3451
rect 9398 3448 9404 3460
rect 9171 3420 9404 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 9692 3457 9720 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 9692 3380 9720 3411
rect 9858 3408 9864 3460
rect 9916 3408 9922 3460
rect 9950 3408 9956 3460
rect 10008 3408 10014 3460
rect 8772 3352 9720 3380
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1762 3136 1768 3188
rect 1820 3136 1826 3188
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3844 3148 3893 3176
rect 3844 3136 3850 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 1489 3111 1547 3117
rect 1489 3077 1501 3111
rect 1535 3108 1547 3111
rect 1780 3108 1808 3136
rect 1535 3080 1808 3108
rect 2041 3111 2099 3117
rect 1535 3077 1547 3080
rect 1489 3071 1547 3077
rect 2041 3077 2053 3111
rect 2087 3108 2099 3111
rect 2222 3108 2228 3120
rect 2087 3080 2228 3108
rect 2087 3077 2099 3080
rect 2041 3071 2099 3077
rect 2222 3068 2228 3080
rect 2280 3068 2286 3120
rect 2332 2972 2360 3136
rect 2593 3111 2651 3117
rect 2593 3077 2605 3111
rect 2639 3108 2651 3111
rect 2639 3080 2774 3108
rect 2639 3077 2651 3080
rect 2593 3071 2651 3077
rect 2746 3040 2774 3080
rect 3896 3040 3924 3139
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4120 3148 4844 3176
rect 4120 3136 4126 3148
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 2746 3012 3832 3040
rect 3896 3012 4629 3040
rect 3804 2972 3832 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4816 3040 4844 3148
rect 5350 3136 5356 3188
rect 5408 3136 5414 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6362 3176 6368 3188
rect 6043 3148 6368 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 4884 3111 4942 3117
rect 4884 3077 4896 3111
rect 4930 3108 4942 3111
rect 5368 3108 5396 3136
rect 4930 3080 5396 3108
rect 4930 3077 4942 3080
rect 4884 3071 4942 3077
rect 5810 3040 5816 3052
rect 4816 3012 5816 3040
rect 4617 3003 4675 3009
rect 5810 3000 5816 3012
rect 5868 3040 5874 3052
rect 6012 3040 6040 3139
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 6822 3136 6828 3188
rect 6880 3136 6886 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 7892 3148 8493 3176
rect 7892 3136 7898 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 8481 3139 8539 3145
rect 8662 3136 8668 3188
rect 8720 3136 8726 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 8846 3136 8852 3188
rect 8904 3136 8910 3188
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 8996 3148 9321 3176
rect 8996 3136 9002 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 9309 3139 9367 3145
rect 10134 3136 10140 3188
rect 10192 3136 10198 3188
rect 6632 3111 6690 3117
rect 6632 3077 6644 3111
rect 6678 3108 6690 3111
rect 6840 3108 6868 3136
rect 6678 3080 6868 3108
rect 6678 3077 6690 3080
rect 6632 3071 6690 3077
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 8386 3108 8392 3120
rect 6972 3080 8392 3108
rect 6972 3068 6978 3080
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 5868 3012 6040 3040
rect 6365 3043 6423 3049
rect 5868 3000 5874 3012
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6454 3040 6460 3052
rect 6411 3012 6460 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8680 3040 8708 3136
rect 8772 3049 8800 3136
rect 8864 3108 8892 3136
rect 9217 3111 9275 3117
rect 9217 3108 9229 3111
rect 8864 3080 9229 3108
rect 9217 3077 9229 3080
rect 9263 3077 9275 3111
rect 9217 3071 9275 3077
rect 8619 3012 8708 3040
rect 8757 3043 8815 3049
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10042 3040 10048 3052
rect 9815 3012 10048 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 4338 2972 4344 2984
rect 2332 2944 2774 2972
rect 3804 2944 4344 2972
rect 1302 2864 1308 2916
rect 1360 2904 1366 2916
rect 1360 2876 2176 2904
rect 1360 2864 1366 2876
rect 382 2796 388 2848
rect 440 2836 446 2848
rect 2148 2845 2176 2876
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 440 2808 1593 2836
rect 440 2796 446 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2805 2191 2839
rect 2746 2836 2774 2944
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 9508 2972 9536 3003
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10152 3049 10180 3136
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 7975 2944 9536 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 5552 2876 6132 2904
rect 5552 2836 5580 2876
rect 2746 2808 5580 2836
rect 6104 2836 6132 2876
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 7944 2904 7972 2935
rect 7800 2876 7972 2904
rect 7800 2864 7806 2876
rect 8202 2864 8208 2916
rect 8260 2864 8266 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8352 2876 9628 2904
rect 8352 2864 8358 2876
rect 8220 2836 8248 2864
rect 9600 2845 9628 2876
rect 6104 2808 8248 2836
rect 9585 2839 9643 2845
rect 2133 2799 2191 2805
rect 9585 2805 9597 2839
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2590 2632 2596 2644
rect 1627 2604 2596 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 4985 2635 5043 2641
rect 3476 2604 4384 2632
rect 3476 2592 3482 2604
rect 3786 2564 3792 2576
rect 2976 2536 3792 2564
rect 2976 2505 3004 2536
rect 3786 2524 3792 2536
rect 3844 2524 3850 2576
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4356 2505 4384 2604
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5074 2632 5080 2644
rect 5031 2604 5080 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6454 2632 6460 2644
rect 5951 2604 6460 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7432 2604 7573 2632
rect 7432 2592 7438 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 7892 2604 9674 2632
rect 7892 2592 7898 2604
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 3108 2468 3157 2496
rect 3108 2456 3114 2468
rect 3145 2465 3157 2468
rect 3191 2465 3203 2499
rect 4341 2499 4399 2505
rect 3145 2459 3203 2465
rect 3252 2468 4292 2496
rect 3252 2440 3280 2468
rect 1394 2388 1400 2440
rect 1452 2388 1458 2440
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 1854 2428 1860 2440
rect 1811 2400 1860 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2096 2400 2513 2428
rect 2096 2388 2102 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 4264 2428 4292 2468
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4982 2496 4988 2508
rect 4571 2468 4988 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 5184 2496 5212 2592
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 7466 2564 7472 2576
rect 5675 2536 7472 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7650 2496 7656 2508
rect 5184 2468 6132 2496
rect 4264 2400 5304 2428
rect 1412 2360 1440 2388
rect 1949 2363 2007 2369
rect 1949 2360 1961 2363
rect 1412 2332 1961 2360
rect 1949 2329 1961 2332
rect 1995 2329 2007 2363
rect 1949 2323 2007 2329
rect 2869 2363 2927 2369
rect 2869 2329 2881 2363
rect 2915 2360 2927 2363
rect 3050 2360 3056 2372
rect 2915 2332 3056 2360
rect 2915 2329 2927 2332
rect 2869 2323 2927 2329
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 5169 2363 5227 2369
rect 5169 2360 5181 2363
rect 4212 2332 5181 2360
rect 4212 2320 4218 2332
rect 5169 2329 5181 2332
rect 5215 2329 5227 2363
rect 5276 2360 5304 2400
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 6104 2437 6132 2468
rect 7024 2468 7656 2496
rect 7024 2437 7052 2468
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7742 2428 7748 2440
rect 7515 2400 7748 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8294 2428 8300 2440
rect 7975 2400 8300 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 6457 2363 6515 2369
rect 6457 2360 6469 2363
rect 5276 2332 6469 2360
rect 5169 2323 5227 2329
rect 6457 2329 6469 2332
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 9033 2363 9091 2369
rect 9033 2360 9045 2363
rect 8527 2332 9045 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 9033 2329 9045 2332
rect 9079 2329 9091 2363
rect 9646 2360 9674 2604
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2428 10287 2431
rect 10410 2428 10416 2440
rect 10275 2400 10416 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 9769 2363 9827 2369
rect 9769 2360 9781 2363
rect 9646 2332 9781 2360
rect 9033 2323 9091 2329
rect 9769 2329 9781 2332
rect 9815 2329 9827 2363
rect 9769 2323 9827 2329
rect 2222 2252 2228 2304
rect 2280 2252 2286 2304
rect 3970 2252 3976 2304
rect 4028 2252 4034 2304
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 5261 2295 5319 2301
rect 5261 2292 5273 2295
rect 5040 2264 5273 2292
rect 5040 2252 5046 2264
rect 5261 2261 5273 2264
rect 5307 2261 5319 2295
rect 5261 2255 5319 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6236 2264 6561 2292
rect 6236 2252 6242 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6972 2264 7113 2292
rect 6972 2252 6978 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8720 2264 9137 2292
rect 8720 2252 8726 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9732 2264 9873 2292
rect 9732 2252 9738 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10008 2264 10425 2292
rect 10008 2252 10014 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 1946 1980 1952 2032
rect 2004 2020 2010 2032
rect 9950 2020 9956 2032
rect 2004 1992 9956 2020
rect 2004 1980 2010 1992
rect 9950 1980 9956 1992
rect 10008 1980 10014 2032
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 3884 9664 3936 9716
rect 7932 9664 7984 9716
rect 1860 9596 1912 9648
rect 2872 9596 2924 9648
rect 4896 9596 4948 9648
rect 6184 9596 6236 9648
rect 6920 9596 6972 9648
rect 8944 9596 8996 9648
rect 9956 9596 10008 9648
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 1676 9528 1728 9580
rect 2780 9528 2832 9580
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 848 9392 900 9444
rect 7380 9528 7432 9580
rect 7840 9528 7892 9580
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9036 9460 9088 9512
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 7932 9324 7984 9376
rect 8208 9324 8260 9376
rect 9220 9324 9272 9376
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 1492 9120 1544 9172
rect 4068 9120 4120 9172
rect 5080 9120 5132 9172
rect 6184 9120 6236 9172
rect 9312 9120 9364 9172
rect 11060 9120 11112 9172
rect 940 8916 992 8968
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2964 8916 3016 8968
rect 9220 9052 9272 9104
rect 7932 8984 7984 9036
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 7288 8848 7340 8900
rect 7564 8916 7616 8968
rect 8116 8916 8168 8968
rect 7932 8848 7984 8900
rect 1492 8780 1544 8832
rect 5356 8780 5408 8832
rect 7656 8780 7708 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8024 8780 8076 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 8852 8780 8904 8832
rect 9128 8780 9180 8832
rect 10324 8848 10376 8900
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 2688 8576 2740 8628
rect 7564 8576 7616 8628
rect 8116 8576 8168 8628
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 9036 8576 9088 8628
rect 10140 8576 10192 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 6828 8372 6880 8424
rect 7840 8440 7892 8492
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8668 8440 8720 8492
rect 8852 8440 8904 8492
rect 9956 8440 10008 8492
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 7288 8304 7340 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 6920 8236 6972 8288
rect 8852 8304 8904 8356
rect 9036 8372 9088 8424
rect 9864 8372 9916 8424
rect 10416 8304 10468 8356
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 1952 8032 2004 8084
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 2504 8032 2556 8041
rect 2688 7964 2740 8016
rect 6460 8032 6512 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 9036 7896 9088 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 6920 7828 6972 7880
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 10232 7828 10284 7880
rect 1860 7692 1912 7744
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2504 7692 2556 7744
rect 6184 7692 6236 7744
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 8116 7692 8168 7744
rect 9864 7692 9916 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 1400 7488 1452 7540
rect 1952 7488 2004 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 3056 7488 3108 7540
rect 7380 7488 7432 7540
rect 9128 7488 9180 7540
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 8116 7420 8168 7472
rect 10232 7531 10284 7540
rect 10232 7497 10241 7531
rect 10241 7497 10275 7531
rect 10275 7497 10284 7531
rect 10232 7488 10284 7497
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 4344 7352 4396 7404
rect 5540 7352 5592 7404
rect 2596 7284 2648 7336
rect 2872 7216 2924 7268
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 4160 7216 4212 7268
rect 2412 7148 2464 7200
rect 2504 7148 2556 7200
rect 4988 7148 5040 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 5816 7148 5868 7200
rect 6460 7352 6512 7404
rect 7380 7352 7432 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 8300 7352 8352 7404
rect 6828 7148 6880 7200
rect 6920 7148 6972 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 10232 7352 10284 7404
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 10048 7284 10100 7336
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 2596 6944 2648 6996
rect 8668 6944 8720 6996
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 2780 6876 2832 6928
rect 3332 6876 3384 6928
rect 3792 6919 3844 6928
rect 3792 6885 3801 6919
rect 3801 6885 3835 6919
rect 3835 6885 3844 6919
rect 3792 6876 3844 6885
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5724 6808 5776 6860
rect 7564 6808 7616 6860
rect 9220 6876 9272 6928
rect 8852 6808 8904 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3332 6740 3384 6792
rect 2136 6672 2188 6724
rect 3056 6672 3108 6724
rect 3792 6672 3844 6724
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5816 6740 5868 6792
rect 6184 6740 6236 6792
rect 6920 6740 6972 6792
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 4252 6604 4304 6656
rect 4344 6604 4396 6656
rect 5632 6604 5684 6656
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 9220 6672 9272 6724
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 10232 6740 10284 6792
rect 10600 6808 10652 6860
rect 10416 6604 10468 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 940 6264 992 6316
rect 1492 6264 1544 6316
rect 1952 6400 2004 6452
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 5172 6400 5224 6452
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2136 6264 2188 6316
rect 2320 6264 2372 6316
rect 4160 6264 4212 6316
rect 1860 6196 1912 6248
rect 3792 6196 3844 6248
rect 3976 6196 4028 6248
rect 3608 6171 3660 6180
rect 3608 6137 3617 6171
rect 3617 6137 3651 6171
rect 3651 6137 3660 6171
rect 3608 6128 3660 6137
rect 3884 6060 3936 6112
rect 5264 6060 5316 6112
rect 6184 6060 6236 6112
rect 9864 6400 9916 6452
rect 10140 6400 10192 6452
rect 6920 6196 6972 6248
rect 7472 6196 7524 6248
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 8300 6239 8352 6248
rect 8300 6205 8309 6239
rect 8309 6205 8343 6239
rect 8343 6205 8352 6239
rect 8300 6196 8352 6205
rect 7380 6060 7432 6112
rect 7840 6060 7892 6112
rect 8944 6264 8996 6316
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10324 6264 10376 6316
rect 10416 6264 10468 6316
rect 11060 6264 11112 6316
rect 8760 6196 8812 6248
rect 9404 6196 9456 6248
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1492 5856 1544 5908
rect 1584 5856 1636 5908
rect 2412 5856 2464 5908
rect 2596 5856 2648 5908
rect 3056 5856 3108 5908
rect 2504 5788 2556 5840
rect 2780 5788 2832 5840
rect 3976 5856 4028 5908
rect 4712 5856 4764 5908
rect 5080 5856 5132 5908
rect 6460 5856 6512 5908
rect 6828 5856 6880 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 10048 5856 10100 5908
rect 8300 5788 8352 5840
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2412 5652 2464 5704
rect 2780 5652 2832 5704
rect 3608 5720 3660 5772
rect 4068 5720 4120 5772
rect 7564 5720 7616 5772
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3976 5584 4028 5636
rect 4344 5584 4396 5636
rect 5264 5627 5316 5636
rect 5264 5593 5273 5627
rect 5273 5593 5307 5627
rect 5307 5593 5316 5627
rect 5264 5584 5316 5593
rect 7472 5652 7524 5704
rect 7932 5652 7984 5704
rect 8116 5652 8168 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 4988 5516 5040 5568
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 7748 5584 7800 5636
rect 10232 5516 10284 5568
rect 10324 5559 10376 5568
rect 10324 5525 10333 5559
rect 10333 5525 10367 5559
rect 10367 5525 10376 5559
rect 10324 5516 10376 5525
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 1676 5312 1728 5364
rect 1768 5312 1820 5364
rect 3792 5312 3844 5364
rect 3976 5312 4028 5364
rect 8116 5312 8168 5364
rect 9956 5312 10008 5364
rect 10324 5312 10376 5364
rect 10508 5312 10560 5364
rect 2044 5244 2096 5296
rect 940 5176 992 5228
rect 1584 5176 1636 5228
rect 2412 5176 2464 5228
rect 4712 5244 4764 5296
rect 6920 5244 6972 5296
rect 7380 5244 7432 5296
rect 3240 5176 3292 5228
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 6184 5176 6236 5228
rect 7932 5176 7984 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 1860 5108 1912 5160
rect 5632 5108 5684 5160
rect 3056 4972 3108 5024
rect 5724 4972 5776 5024
rect 6920 5108 6972 5160
rect 6460 5040 6512 5092
rect 7840 5108 7892 5160
rect 8944 5176 8996 5228
rect 9128 5108 9180 5160
rect 6552 4972 6604 5024
rect 9404 5176 9456 5228
rect 9956 5108 10008 5160
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 1676 4768 1728 4820
rect 1952 4768 2004 4820
rect 2780 4768 2832 4820
rect 3240 4768 3292 4820
rect 4252 4768 4304 4820
rect 5540 4768 5592 4820
rect 3056 4632 3108 4684
rect 3792 4632 3844 4684
rect 6460 4768 6512 4820
rect 6920 4768 6972 4820
rect 8024 4768 8076 4820
rect 8944 4768 8996 4820
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 10048 4768 10100 4820
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 1860 4564 1912 4616
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 2320 4564 2372 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 2504 4496 2556 4548
rect 5172 4564 5224 4616
rect 5172 4428 5224 4480
rect 6184 4564 6236 4616
rect 6552 4564 6604 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 7932 4564 7984 4616
rect 6552 4428 6604 4480
rect 7472 4496 7524 4548
rect 8668 4496 8720 4548
rect 7748 4428 7800 4480
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1860 4224 1912 4276
rect 1952 4224 2004 4276
rect 2136 4224 2188 4276
rect 2320 4224 2372 4276
rect 1768 4156 1820 4208
rect 1400 4088 1452 4140
rect 5724 4224 5776 4276
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 10324 4224 10376 4276
rect 10508 4224 10560 4276
rect 1860 4020 1912 4072
rect 3148 4088 3200 4140
rect 3240 4088 3292 4140
rect 3976 4156 4028 4208
rect 9864 4156 9916 4208
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 2412 3884 2464 3936
rect 4068 4088 4120 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4528 4088 4580 4140
rect 5448 4088 5500 4140
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 4436 4063 4488 4072
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 4896 4020 4948 4072
rect 6368 4063 6420 4072
rect 6368 4029 6377 4063
rect 6377 4029 6411 4063
rect 6411 4029 6420 4063
rect 6368 4020 6420 4029
rect 7472 4020 7524 4072
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 3700 3884 3752 3936
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 5080 3884 5132 3936
rect 6184 3952 6236 4004
rect 6644 3884 6696 3936
rect 6828 3884 6880 3936
rect 8668 3884 8720 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 10232 3884 10284 3936
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 2596 3680 2648 3732
rect 4436 3680 4488 3732
rect 6184 3680 6236 3732
rect 2504 3544 2556 3596
rect 2780 3544 2832 3596
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 6920 3612 6972 3664
rect 3700 3544 3752 3596
rect 5080 3544 5132 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 6460 3544 6512 3596
rect 7380 3680 7432 3732
rect 8116 3680 8168 3732
rect 8668 3680 8720 3732
rect 8852 3544 8904 3596
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 4436 3408 4488 3460
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 4620 3408 4672 3460
rect 5356 3340 5408 3392
rect 6552 3408 6604 3460
rect 7840 3408 7892 3460
rect 8668 3340 8720 3392
rect 9404 3408 9456 3460
rect 9864 3451 9916 3460
rect 9864 3417 9873 3451
rect 9873 3417 9907 3451
rect 9907 3417 9916 3451
rect 9864 3408 9916 3417
rect 9956 3451 10008 3460
rect 9956 3417 9965 3451
rect 9965 3417 9999 3451
rect 9999 3417 10008 3451
rect 9956 3408 10008 3417
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 1768 3136 1820 3188
rect 2320 3136 2372 3188
rect 3792 3136 3844 3188
rect 2228 3068 2280 3120
rect 4068 3136 4120 3188
rect 5356 3136 5408 3188
rect 5816 3000 5868 3052
rect 6368 3136 6420 3188
rect 6828 3136 6880 3188
rect 7840 3136 7892 3188
rect 8668 3136 8720 3188
rect 8760 3136 8812 3188
rect 8852 3136 8904 3188
rect 8944 3136 8996 3188
rect 10140 3136 10192 3188
rect 6920 3068 6972 3120
rect 8392 3068 8444 3120
rect 6460 3000 6512 3052
rect 1308 2864 1360 2916
rect 388 2796 440 2848
rect 4344 2932 4396 2984
rect 10048 3000 10100 3052
rect 7748 2907 7800 2916
rect 7748 2873 7757 2907
rect 7757 2873 7791 2907
rect 7791 2873 7800 2907
rect 7748 2864 7800 2873
rect 8208 2864 8260 2916
rect 8300 2864 8352 2916
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 2596 2592 2648 2644
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 3792 2524 3844 2576
rect 3056 2456 3108 2508
rect 5080 2592 5132 2644
rect 5172 2592 5224 2644
rect 6460 2592 6512 2644
rect 7380 2592 7432 2644
rect 7840 2592 7892 2644
rect 1400 2388 1452 2440
rect 1860 2388 1912 2440
rect 2044 2388 2096 2440
rect 3240 2388 3292 2440
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 4988 2456 5040 2508
rect 7472 2524 7524 2576
rect 3056 2320 3108 2372
rect 4160 2320 4212 2372
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 7656 2456 7708 2508
rect 7748 2388 7800 2440
rect 8300 2388 8352 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 10416 2388 10468 2440
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 4988 2252 5040 2304
rect 6184 2252 6236 2304
rect 6920 2252 6972 2304
rect 7748 2252 7800 2304
rect 8668 2252 8720 2304
rect 9680 2252 9732 2304
rect 9956 2252 10008 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 1952 1980 2004 2032
rect 9956 1980 10008 2032
<< metal2 >>
rect 846 11200 902 12000
rect 1858 11200 1914 12000
rect 2870 11200 2926 12000
rect 3882 11200 3938 12000
rect 4894 11200 4950 12000
rect 5906 11200 5962 12000
rect 6012 11206 6224 11234
rect 860 9450 888 11200
rect 1872 9654 1900 11200
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 2792 9586 2820 10911
rect 2884 9654 2912 11200
rect 2962 10160 3018 10169
rect 2962 10095 3018 10104
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 848 9444 900 9450
rect 848 9386 900 9392
rect 1504 9178 1532 9522
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 952 8974 980 9007
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7546 1440 8230
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 1398 6896 1454 6905
rect 1504 6882 1532 8774
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8265 1624 8434
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1504 6854 1624 6882
rect 1398 6831 1454 6840
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 952 5817 980 6258
rect 1504 5914 1532 6258
rect 1596 5914 1624 6854
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 938 5808 994 5817
rect 1688 5794 1716 9522
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8090 1992 8910
rect 2700 8634 2728 9318
rect 2976 8974 3004 10095
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3896 9722 3924 11200
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 4908 9654 4936 11200
rect 5920 11098 5948 11200
rect 6012 11098 6040 11206
rect 5920 11070 6040 11098
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6196 9654 6224 11206
rect 6918 11200 6974 12000
rect 7930 11200 7986 12000
rect 8942 11200 8998 12000
rect 9310 11248 9366 11257
rect 6932 9654 6960 11200
rect 7944 9722 7972 11200
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8956 9654 8984 11200
rect 9954 11200 10010 12000
rect 10966 11200 11022 12000
rect 9310 11183 9366 11192
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 938 5743 994 5752
rect 1412 5766 1716 5794
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4729 980 5170
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1412 4146 1440 5766
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1308 2916 1360 2922
rect 1308 2858 1360 2864
rect 388 2848 440 2854
rect 388 2790 440 2796
rect 400 800 428 2790
rect 1320 800 1348 2858
rect 1504 2774 1532 5510
rect 1688 5370 1716 5646
rect 1780 5370 1808 7822
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1872 6254 1900 7686
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1964 6458 1992 7482
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5817 1900 6190
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4049 1624 5170
rect 1688 4826 1716 5306
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1412 2746 1532 2774
rect 1412 2446 1440 2746
rect 1688 2689 1716 4558
rect 1780 4214 1808 5306
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1872 4622 1900 5102
rect 1964 4826 1992 6258
rect 2056 5658 2084 7686
rect 2332 7313 2360 7822
rect 2516 7750 2544 8026
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2596 7336 2648 7342
rect 2318 7304 2374 7313
rect 2502 7304 2558 7313
rect 2318 7239 2374 7248
rect 2424 7262 2502 7290
rect 2424 7206 2452 7262
rect 2596 7278 2648 7284
rect 2700 7290 2728 7958
rect 3068 7546 3096 9522
rect 4080 9178 4108 9522
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 5092 9178 5120 9522
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9178 6224 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 2502 7239 2558 7248
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2148 6322 2176 6666
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2320 6316 2372 6322
rect 2516 6304 2544 7142
rect 2608 7002 2636 7278
rect 2700 7262 2774 7290
rect 2746 7018 2774 7262
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2700 6990 2774 7018
rect 2372 6276 2544 6304
rect 2320 6258 2372 6264
rect 2148 6225 2176 6258
rect 2134 6216 2190 6225
rect 2134 6151 2190 6160
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2608 5914 2636 6938
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2424 5710 2452 5850
rect 2504 5840 2556 5846
rect 2556 5788 2636 5794
rect 2504 5782 2636 5788
rect 2516 5766 2636 5782
rect 2412 5704 2464 5710
rect 2056 5630 2176 5658
rect 2412 5646 2464 5652
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5302 2084 5510
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2148 5148 2176 5630
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5234 2452 5510
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2056 5120 2176 5148
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1872 4282 1900 4558
rect 1964 4282 1992 4762
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1768 4208 1820 4214
rect 1768 4150 1820 4156
rect 1860 4072 1912 4078
rect 1912 4032 1992 4060
rect 1860 4014 1912 4020
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3194 1808 3878
rect 1858 3632 1914 3641
rect 1858 3567 1914 3576
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1674 2680 1730 2689
rect 1674 2615 1730 2624
rect 1872 2446 1900 3567
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1964 2038 1992 4032
rect 2056 2446 2084 5120
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2148 4282 2176 4558
rect 2332 4282 2360 4558
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2424 3942 2452 4558
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2516 3602 2544 4490
rect 2608 3738 2636 5766
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2320 3528 2372 3534
rect 2700 3482 2728 6990
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2792 5846 2820 6870
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 4826 2820 5646
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2884 4536 2912 7210
rect 3252 7041 3280 7346
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3344 6934 3372 7346
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3344 6798 3372 6870
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2792 4508 2912 4536
rect 2792 3602 2820 4508
rect 2976 4434 3004 6598
rect 3068 5914 3096 6666
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4690 3096 4966
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2884 4406 3004 4434
rect 2884 4196 2912 4406
rect 2884 4168 3004 4196
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2320 3470 2372 3476
rect 2332 3194 2360 3470
rect 2424 3454 2728 3482
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2228 3120 2280 3126
rect 2424 3074 2452 3454
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2280 3068 2452 3074
rect 2228 3062 2452 3068
rect 2240 3046 2452 3062
rect 2516 2961 2544 3334
rect 2502 2952 2558 2961
rect 2502 2887 2558 2896
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2594 2680 2650 2689
rect 2594 2615 2596 2624
rect 2648 2615 2650 2624
rect 2596 2586 2648 2592
rect 2976 2496 3004 4168
rect 3160 4146 3188 6734
rect 3804 6730 3832 6870
rect 4080 6866 4108 7278
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 4172 6474 4200 7210
rect 4356 6662 4384 7346
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4080 6446 4200 6474
rect 3792 6248 3844 6254
rect 3330 6216 3386 6225
rect 3252 6174 3330 6202
rect 3252 5234 3280 6174
rect 3792 6190 3844 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3330 6151 3386 6160
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3620 5778 3648 6122
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3804 5370 3832 6190
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3252 4146 3280 4762
rect 3804 4690 3832 5170
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3712 3942 3740 3975
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3160 2632 3188 3878
rect 3698 3632 3754 3641
rect 3698 3567 3700 3576
rect 3752 3567 3754 3576
rect 3700 3538 3752 3544
rect 3606 3496 3662 3505
rect 3606 3431 3662 3440
rect 3620 3398 3648 3431
rect 3332 3392 3384 3398
rect 3252 3352 3332 3380
rect 3252 2774 3280 3352
rect 3332 3334 3384 3340
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3804 3194 3832 4626
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3896 2774 3924 6054
rect 3988 5914 4016 6190
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5778 4108 6446
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 3988 5370 4016 5578
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3988 4214 4016 5306
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4080 4146 4108 5714
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3252 2746 3464 2774
rect 3436 2650 3464 2746
rect 3804 2746 3924 2774
rect 3424 2644 3476 2650
rect 3160 2604 3280 2632
rect 3056 2508 3108 2514
rect 2976 2468 3056 2496
rect 3056 2450 3108 2456
rect 3252 2446 3280 2604
rect 3424 2586 3476 2592
rect 3804 2582 3832 2746
rect 3792 2576 3844 2582
rect 3988 2564 4016 3878
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3194 4108 3470
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4172 2774 4200 6258
rect 4264 5794 4292 6598
rect 4356 6458 4384 6598
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4264 5766 4568 5794
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4264 4146 4292 4762
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4356 2990 4384 5578
rect 4540 4146 4568 5766
rect 4724 5302 4752 5850
rect 5000 5658 5028 7142
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5092 5914 5120 6734
rect 5184 6458 5212 6734
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5000 5630 5120 5658
rect 5276 5642 5304 6054
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 5000 4706 5028 5510
rect 4908 4678 5028 4706
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4908 4078 4936 4678
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4896 4072 4948 4078
rect 5092 4026 5120 5630
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 4622 5212 5510
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4896 4014 4948 4020
rect 4448 3738 4476 4014
rect 5000 3998 5120 4026
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4436 3460 4488 3466
rect 4620 3460 4672 3466
rect 4488 3420 4620 3448
rect 4436 3402 4488 3408
rect 4620 3402 4672 3408
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 3792 2518 3844 2524
rect 3896 2536 4016 2564
rect 4080 2746 4200 2774
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 3896 2446 3924 2536
rect 2044 2440 2096 2446
rect 3240 2440 3292 2446
rect 2044 2382 2096 2388
rect 3068 2378 3188 2394
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3056 2372 3188 2378
rect 3108 2366 3188 2372
rect 3056 2314 3108 2320
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 2240 800 2268 2246
rect 3160 800 3188 2366
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3988 1170 4016 2246
rect 4080 1465 4108 2746
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 4158 2544 4214 2553
rect 5000 2514 5028 3998
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3602 5120 3878
rect 5184 3641 5212 4422
rect 5368 4049 5396 8774
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 6472 8090 6500 8910
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5446 5808 5502 5817
rect 5446 5743 5502 5752
rect 5460 4146 5488 5743
rect 5552 4826 5580 7346
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5736 6866 5764 7142
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5828 6798 5856 7142
rect 6196 6798 6224 7686
rect 6472 7410 6500 8026
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 5166 5672 6598
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6196 5234 6224 6054
rect 6472 5914 6500 7346
rect 6840 7206 6868 8366
rect 7300 8362 7328 8842
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7886 6960 8230
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7392 7546 7420 9522
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7576 8634 7604 8910
rect 7852 8838 7880 9522
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7944 9042 7972 9318
rect 8220 9081 8248 9318
rect 8206 9072 8262 9081
rect 7932 9036 7984 9042
rect 8206 9007 8262 9016
rect 7932 8978 7984 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7484 7410 7512 7686
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6840 6610 6868 7142
rect 6932 6798 6960 7142
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6840 6582 6960 6610
rect 6932 6254 6960 6582
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7392 6118 7420 7346
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6866 7604 7142
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6840 5386 6868 5850
rect 7484 5710 7512 6190
rect 7576 5778 7604 6190
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 6840 5358 6960 5386
rect 6932 5302 6960 5358
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5736 4282 5764 4966
rect 6472 4826 6500 5034
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6564 4622 6592 4966
rect 6932 4826 6960 5102
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7392 4690 7420 5238
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 6196 4162 6224 4558
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 6104 4134 6224 4162
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 5170 3632 5226 3641
rect 5080 3596 5132 3602
rect 5170 3567 5172 3576
rect 5080 3538 5132 3544
rect 5224 3567 5226 3576
rect 6104 3584 6132 4134
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6196 3738 6224 3946
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6184 3596 6236 3602
rect 6104 3556 6184 3584
rect 5172 3538 5224 3544
rect 6184 3538 6236 3544
rect 5092 2650 5120 3538
rect 5184 2650 5212 3538
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3194 5396 3334
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 6380 3194 6408 4014
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6472 3058 6500 3538
rect 6564 3466 6592 4422
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3641 6684 3878
rect 6642 3632 6698 3641
rect 6642 3567 6698 3576
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 4158 2479 4214 2488
rect 4988 2508 5040 2514
rect 4172 2378 4200 2479
rect 4988 2450 5040 2456
rect 5828 2446 5856 2994
rect 6748 2774 6776 4558
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3194 6868 3878
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7392 3738 7420 4626
rect 7472 4548 7524 4554
rect 7524 4508 7604 4536
rect 7472 4490 7524 4496
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6932 3126 6960 3606
rect 7484 3380 7512 4014
rect 7392 3352 7512 3380
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6472 2746 6776 2774
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 6472 2650 6500 2746
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7392 2650 7420 3352
rect 7576 2774 7604 4508
rect 7484 2746 7604 2774
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2582 7512 2746
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7668 2514 7696 8774
rect 7852 8498 7880 8774
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5914 7788 6190
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7760 4486 7788 5578
rect 7852 5166 7880 6054
rect 7944 5710 7972 8842
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8498 8064 8774
rect 8128 8634 8156 8910
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8680 8634 8708 8774
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8680 8498 8708 8570
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7478 8156 7686
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 6798 8340 7346
rect 8680 7002 8708 7822
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8772 6254 8800 9522
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8498 8892 8774
rect 9048 8634 9076 9454
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9110 9260 9318
rect 9324 9178 9352 11183
rect 9968 9654 9996 11200
rect 10598 10160 10654 10169
rect 10598 10095 10654 10104
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8864 6866 8892 8298
rect 9048 7954 9076 8366
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9140 7546 9168 8774
rect 10152 8634 10180 9522
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 8090 9444 8230
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9876 7750 9904 8366
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7546 9904 7686
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9968 7426 9996 8434
rect 9876 7398 9996 7426
rect 10060 7426 10088 8434
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 7546 10272 7822
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10060 7398 10180 7426
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6934 9260 7278
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9876 6984 9904 7398
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10060 7002 10088 7278
rect 9784 6956 9904 6984
rect 10048 6996 10100 7002
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8956 6322 8984 6802
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6322 9260 6666
rect 9784 6338 9812 6956
rect 10048 6938 10100 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6458 9904 6734
rect 10152 6458 10180 7398
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 6798 10272 7346
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9220 6316 9272 6322
rect 9784 6310 9904 6338
rect 10336 6322 10364 8842
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 6662 10456 8298
rect 10506 6896 10562 6905
rect 10612 6866 10640 10095
rect 10980 10010 11008 11200
rect 10980 9982 11100 10010
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 11072 9178 11100 9982
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 11058 7984 11114 7993
rect 11058 7919 11114 7928
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10506 6831 10562 6840
rect 10600 6860 10652 6866
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 9220 6258 9272 6264
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 8312 5846 8340 6190
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8128 5370 8156 5646
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7944 4622 7972 5170
rect 8036 4826 8064 5170
rect 8956 4826 8984 5170
rect 9140 5166 9168 5646
rect 9416 5234 9444 6190
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9876 4706 9904 6310
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 9968 5370 9996 6258
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5914 10088 6054
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10428 5817 10456 6258
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9968 5250 9996 5306
rect 9968 5222 10088 5250
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4826 9996 5102
rect 10060 4826 10088 5222
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9876 4678 10088 4706
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8680 4282 8708 4490
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8482 4040 8538 4049
rect 8128 3738 8156 4014
rect 8482 3975 8538 3984
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8496 3534 8524 3975
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8680 3738 8708 3878
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 3194 7880 3402
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8680 3194 8708 3334
rect 8772 3194 8800 3878
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8864 3194 8892 3538
rect 8956 3194 8984 4082
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3466 9444 3878
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9876 3466 9904 4150
rect 9954 3496 10010 3505
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9864 3460 9916 3466
rect 9954 3431 9956 3440
rect 9864 3402 9916 3408
rect 10008 3431 10010 3440
rect 9956 3402 10008 3408
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 7838 2952 7894 2961
rect 7748 2916 7800 2922
rect 7838 2887 7894 2896
rect 8208 2916 8260 2922
rect 7748 2858 7800 2864
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7760 2446 7788 2858
rect 7852 2650 7880 2887
rect 8208 2858 8260 2864
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8220 2553 8248 2858
rect 8206 2544 8262 2553
rect 8206 2479 8262 2488
rect 8312 2446 8340 2858
rect 8404 2446 8432 3062
rect 10060 3058 10088 4678
rect 10244 3942 10272 5510
rect 10336 5370 10364 5510
rect 10520 5370 10548 6831
rect 10600 6802 10652 6808
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 11072 6322 11100 7919
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10336 4282 10364 5306
rect 10506 4720 10562 4729
rect 10506 4655 10562 4664
rect 10520 4282 10548 4655
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10152 3194 10180 3878
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 10428 2530 10456 2790
rect 10428 2502 10548 2530
rect 5816 2440 5868 2446
rect 7748 2440 7800 2446
rect 5816 2382 5868 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 6840 2366 6960 2394
rect 7748 2382 7800 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8392 2440 8444 2446
rect 10416 2440 10468 2446
rect 8392 2382 8444 2388
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 3988 1142 4108 1170
rect 4080 800 4108 1142
rect 5000 800 5028 2246
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 5920 870 6040 898
rect 5920 800 5948 870
rect 386 0 442 800
rect 1306 0 1362 800
rect 2226 0 2282 800
rect 3146 0 3202 800
rect 4066 0 4122 800
rect 4986 0 5042 800
rect 5906 0 5962 800
rect 6012 762 6040 870
rect 6196 762 6224 2246
rect 6840 800 6868 2366
rect 6932 2310 6960 2366
rect 9600 2366 9720 2394
rect 10416 2382 10468 2388
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 7760 800 7788 2246
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8680 800 8708 2246
rect 9600 800 9628 2366
rect 9692 2310 9720 2366
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 2038 9996 2246
rect 9956 2032 10008 2038
rect 9956 1974 10008 1980
rect 10428 1465 10456 2382
rect 10414 1456 10470 1465
rect 10414 1391 10470 1400
rect 10520 800 10548 2502
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 6012 734 6224 762
rect 6826 0 6882 800
rect 7746 0 7802 800
rect 8666 0 8722 800
rect 9586 0 9642 800
rect 10506 0 10562 800
<< via2 >>
rect 2778 10920 2834 10976
rect 2962 10104 3018 10160
rect 938 9016 994 9072
rect 1398 6840 1454 6896
rect 1582 8200 1638 8256
rect 938 5752 994 5808
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 9310 11192 9366 11248
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 938 4664 994 4720
rect 1858 5752 1914 5808
rect 1582 3984 1638 4040
rect 2318 7248 2374 7304
rect 2502 7248 2558 7304
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2134 6160 2190 6216
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 1858 3576 1914 3632
rect 1674 2624 1730 2680
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 3238 6976 3294 7032
rect 2502 2896 2558 2952
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 2594 2644 2650 2680
rect 2594 2624 2596 2644
rect 2596 2624 2648 2644
rect 2648 2624 2650 2644
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 3330 6160 3386 6216
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3698 3984 3754 4040
rect 3698 3596 3754 3632
rect 3698 3576 3700 3596
rect 3700 3576 3752 3596
rect 3752 3576 3754 3596
rect 3606 3440 3662 3496
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 4158 2488 4214 2544
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5446 5752 5502 5808
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 8206 9016 8262 9072
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 5354 3984 5410 4040
rect 5170 3596 5226 3632
rect 5170 3576 5172 3596
rect 5172 3576 5224 3596
rect 5224 3576 5226 3596
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 6642 3576 6698 3632
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 10598 10104 10654 10160
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10506 6840 10562 6896
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 11058 7928 11114 7984
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 10414 5752 10470 5808
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 8482 3984 8538 4040
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9954 3460 10010 3496
rect 9954 3440 9956 3460
rect 9956 3440 10008 3460
rect 10008 3440 10010 3460
rect 7838 2896 7894 2952
rect 8206 2488 8262 2544
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10506 4664 10562 4720
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 4066 1400 4122 1456
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10414 1400 10470 1456
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
<< metal3 >>
rect 0 11250 800 11280
rect 9305 11250 9371 11253
rect 11200 11250 12000 11280
rect 0 11190 1410 11250
rect 0 11160 800 11190
rect 1350 10978 1410 11190
rect 9305 11248 12000 11250
rect 9305 11192 9310 11248
rect 9366 11192 12000 11248
rect 9305 11190 12000 11192
rect 9305 11187 9371 11190
rect 11200 11160 12000 11190
rect 2773 10978 2839 10981
rect 1350 10976 2839 10978
rect 1350 10920 2778 10976
rect 2834 10920 2839 10976
rect 1350 10918 2839 10920
rect 2773 10915 2839 10918
rect 0 10162 800 10192
rect 2957 10162 3023 10165
rect 0 10160 3023 10162
rect 0 10104 2962 10160
rect 3018 10104 3023 10160
rect 0 10102 3023 10104
rect 0 10072 800 10102
rect 2957 10099 3023 10102
rect 10593 10162 10659 10165
rect 11200 10162 12000 10192
rect 10593 10160 12000 10162
rect 10593 10104 10598 10160
rect 10654 10104 12000 10160
rect 10593 10102 12000 10104
rect 10593 10099 10659 10102
rect 11200 10072 12000 10102
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 8201 9074 8267 9077
rect 11200 9074 12000 9104
rect 8201 9072 12000 9074
rect 8201 9016 8206 9072
rect 8262 9016 12000 9072
rect 8201 9014 12000 9016
rect 8201 9011 8267 9014
rect 11200 8984 12000 9014
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 1577 8258 1643 8261
rect 798 8256 1643 8258
rect 798 8200 1582 8256
rect 1638 8200 1643 8256
rect 798 8198 1643 8200
rect 798 8016 858 8198
rect 1577 8195 1643 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7926 858 8016
rect 11053 7986 11119 7989
rect 11200 7986 12000 8016
rect 11053 7984 12000 7986
rect 11053 7928 11058 7984
rect 11114 7928 12000 7984
rect 11053 7926 12000 7928
rect 0 7896 800 7926
rect 11053 7923 11119 7926
rect 11200 7896 12000 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 1894 7244 1900 7308
rect 1964 7306 1970 7308
rect 2313 7306 2379 7309
rect 1964 7304 2379 7306
rect 1964 7248 2318 7304
rect 2374 7248 2379 7304
rect 1964 7246 2379 7248
rect 1964 7244 1970 7246
rect 2313 7243 2379 7246
rect 2497 7306 2563 7309
rect 2630 7306 2636 7308
rect 2497 7304 2636 7306
rect 2497 7248 2502 7304
rect 2558 7248 2636 7304
rect 2497 7246 2636 7248
rect 2497 7243 2563 7246
rect 2630 7244 2636 7246
rect 2700 7244 2706 7308
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 2814 6972 2820 7036
rect 2884 7034 2890 7036
rect 3233 7034 3299 7037
rect 2884 7032 3299 7034
rect 2884 6976 3238 7032
rect 3294 6976 3299 7032
rect 2884 6974 3299 6976
rect 2884 6972 2890 6974
rect 3233 6971 3299 6974
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 10501 6898 10567 6901
rect 11200 6898 12000 6928
rect 10501 6896 12000 6898
rect 10501 6840 10506 6896
rect 10562 6840 12000 6896
rect 10501 6838 12000 6840
rect 10501 6835 10567 6838
rect 11200 6808 12000 6838
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2129 6218 2195 6221
rect 3325 6218 3391 6221
rect 2129 6216 3391 6218
rect 2129 6160 2134 6216
rect 2190 6160 3330 6216
rect 3386 6160 3391 6216
rect 2129 6158 3391 6160
rect 2129 6155 2195 6158
rect 3325 6155 3391 6158
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 1853 5810 1919 5813
rect 5441 5810 5507 5813
rect 1853 5808 5507 5810
rect 1853 5752 1858 5808
rect 1914 5752 5446 5808
rect 5502 5752 5507 5808
rect 1853 5750 5507 5752
rect 1853 5747 1919 5750
rect 5441 5747 5507 5750
rect 10409 5810 10475 5813
rect 11200 5810 12000 5840
rect 10409 5808 12000 5810
rect 10409 5752 10414 5808
rect 10470 5752 12000 5808
rect 10409 5750 12000 5752
rect 10409 5747 10475 5750
rect 11200 5720 12000 5750
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 10501 4722 10567 4725
rect 11200 4722 12000 4752
rect 10501 4720 12000 4722
rect 10501 4664 10506 4720
rect 10562 4664 12000 4720
rect 10501 4662 12000 4664
rect 10501 4659 10567 4662
rect 11200 4632 12000 4662
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 1577 4042 1643 4045
rect 982 4040 1643 4042
rect 982 3984 1582 4040
rect 1638 3984 1643 4040
rect 982 3982 1643 3984
rect 0 3634 800 3664
rect 982 3634 1042 3982
rect 1577 3979 1643 3982
rect 3693 4042 3759 4045
rect 5349 4042 5415 4045
rect 8477 4042 8543 4045
rect 3693 4040 8543 4042
rect 3693 3984 3698 4040
rect 3754 3984 5354 4040
rect 5410 3984 8482 4040
rect 8538 3984 8543 4040
rect 3693 3982 8543 3984
rect 3693 3979 3759 3982
rect 5349 3979 5415 3982
rect 8477 3979 8543 3982
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 0 3574 1042 3634
rect 1853 3634 1919 3637
rect 3693 3634 3759 3637
rect 5165 3634 5231 3637
rect 1853 3632 5231 3634
rect 1853 3576 1858 3632
rect 1914 3576 3698 3632
rect 3754 3576 5170 3632
rect 5226 3576 5231 3632
rect 1853 3574 5231 3576
rect 0 3544 800 3574
rect 1853 3571 1919 3574
rect 3693 3571 3759 3574
rect 5165 3571 5231 3574
rect 6637 3634 6703 3637
rect 11200 3634 12000 3664
rect 6637 3632 12000 3634
rect 6637 3576 6642 3632
rect 6698 3576 12000 3632
rect 6637 3574 12000 3576
rect 6637 3571 6703 3574
rect 11200 3544 12000 3574
rect 3601 3498 3667 3501
rect 9949 3498 10015 3501
rect 3601 3496 10015 3498
rect 3601 3440 3606 3496
rect 3662 3440 9954 3496
rect 10010 3440 10015 3496
rect 3601 3438 10015 3440
rect 3601 3435 3667 3438
rect 9949 3435 10015 3438
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 2497 2954 2563 2957
rect 7833 2954 7899 2957
rect 2497 2952 7899 2954
rect 2497 2896 2502 2952
rect 2558 2896 7838 2952
rect 7894 2896 7899 2952
rect 2497 2894 7899 2896
rect 2497 2891 2563 2894
rect 7833 2891 7899 2894
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 1669 2682 1735 2685
rect 798 2680 1735 2682
rect 798 2624 1674 2680
rect 1730 2624 1735 2680
rect 798 2622 1735 2624
rect 798 2576 858 2622
rect 1669 2619 1735 2622
rect 2589 2682 2655 2685
rect 2814 2682 2820 2684
rect 2589 2680 2820 2682
rect 2589 2624 2594 2680
rect 2650 2624 2820 2680
rect 2589 2622 2820 2624
rect 2589 2619 2655 2622
rect 2814 2620 2820 2622
rect 2884 2620 2890 2684
rect 0 2486 858 2576
rect 0 2456 800 2486
rect 2630 2484 2636 2548
rect 2700 2546 2706 2548
rect 4153 2546 4219 2549
rect 2700 2544 4219 2546
rect 2700 2488 4158 2544
rect 4214 2488 4219 2544
rect 2700 2486 4219 2488
rect 2700 2484 2706 2486
rect 4153 2483 4219 2486
rect 8201 2546 8267 2549
rect 11200 2546 12000 2576
rect 8201 2544 12000 2546
rect 8201 2488 8206 2544
rect 8262 2488 12000 2544
rect 8201 2486 12000 2488
rect 8201 2483 8267 2486
rect 11200 2456 12000 2486
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 10409 1458 10475 1461
rect 11200 1458 12000 1488
rect 10409 1456 12000 1458
rect 10409 1400 10414 1456
rect 10470 1400 12000 1456
rect 10409 1398 12000 1400
rect 10409 1395 10475 1398
rect 11200 1368 12000 1398
rect 1894 308 1900 372
rect 1964 370 1970 372
rect 11200 370 12000 400
rect 1964 310 12000 370
rect 1964 308 1970 310
rect 11200 280 12000 310
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 1900 7244 1964 7308
rect 2636 7244 2700 7308
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 2820 6972 2884 7036
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 2820 2620 2884 2684
rect 2636 2484 2700 2548
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
rect 1900 308 1964 372
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 1899 7308 1965 7309
rect 1899 7244 1900 7308
rect 1964 7244 1965 7308
rect 1899 7243 1965 7244
rect 1902 373 1962 7243
rect 2163 7104 2483 8128
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 2635 7308 2701 7309
rect 2635 7244 2636 7308
rect 2700 7244 2701 7308
rect 2635 7243 2701 7244
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 2638 2549 2698 7243
rect 2819 7036 2885 7037
rect 2819 6972 2820 7036
rect 2884 6972 2885 7036
rect 2819 6971 2885 6972
rect 2822 2685 2882 6971
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 2819 2684 2885 2685
rect 2819 2620 2820 2684
rect 2884 2620 2885 2684
rect 2819 2619 2885 2620
rect 2635 2548 2701 2549
rect 2635 2484 2636 2548
rect 2700 2484 2701 2548
rect 2635 2483 2701 2484
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
rect 1899 372 1965 373
rect 1899 308 1900 372
rect 1964 308 1965 372
rect 1899 307 1965 308
use sky130_fd_sc_hd__inv_2  _059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1688980957
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1688980957
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1688980957
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1688980957
transform 1 0 1472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1688980957
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1688980957
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130_
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _132_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _133_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 1688980957
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 1688980957
transform 1 0 3956 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _137_
timestamp 1688980957
transform 1 0 3772 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 1688980957
transform 1 0 2208 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 1688980957
transform 1 0 1472 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp 1688980957
transform 1 0 8096 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _143_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1688980957
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform 1 0 1472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _167__44 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _167_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _168_
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _169_
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _170_
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _171_
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _172_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _173_
timestamp 1688980957
transform 1 0 5152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _174_
timestamp 1688980957
transform 1 0 7544 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _175_
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _176_
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _177_
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _178_
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _179_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _180__45
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _180_
timestamp 1688980957
transform 1 0 5796 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _181_
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _182_
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _183_
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _184_
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _185_
timestamp 1688980957
transform 1 0 4324 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _186_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _187_
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _188_
timestamp 1688980957
transform 1 0 5152 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _189_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _190_
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _191__46
timestamp 1688980957
transform 1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _191_
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _192_
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _193_
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _194_
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _195__47
timestamp 1688980957
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _195_
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _196_
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _197_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _198_
timestamp 1688980957
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _199__48
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _199_
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _200_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _201_
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _202_
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_91
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_102
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_36
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_95
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_52
timestamp 1688980957
transform 1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_63
timestamp 1688980957
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_42
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_52
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_74
timestamp 1688980957
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_95
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_50
timestamp 1688980957
transform 1 0 5704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_99
timestamp 1688980957
transform 1 0 10212 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_46
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_68
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_74
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_101
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_89
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_99
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_40
timestamp 1688980957
transform 1 0 4784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_6
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_31
timestamp 1688980957
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_41
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_49
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_68
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_8
timestamp 1688980957
transform 1 0 1840 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_66
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_94
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_48
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_57
timestamp 1688980957
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_18
timestamp 1688980957
transform 1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 3956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 6992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 8004 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 5060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal3 s 11200 10072 12000 10192 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 11200 11160 12000 11280 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 5 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 6 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 7 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 8 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 9 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 10 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 11 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 12 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 13 nsew signal input
flabel metal2 s 846 11200 902 12000 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 14 nsew signal tristate
flabel metal2 s 1858 11200 1914 12000 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 15 nsew signal tristate
flabel metal2 s 2870 11200 2926 12000 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 16 nsew signal tristate
flabel metal2 s 3882 11200 3938 12000 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 17 nsew signal tristate
flabel metal2 s 4894 11200 4950 12000 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 18 nsew signal tristate
flabel metal2 s 5906 11200 5962 12000 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 19 nsew signal tristate
flabel metal2 s 6918 11200 6974 12000 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 20 nsew signal tristate
flabel metal2 s 7930 11200 7986 12000 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 21 nsew signal tristate
flabel metal2 s 8942 11200 8998 12000 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 22 nsew signal tristate
flabel metal3 s 11200 280 12000 400 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 23 nsew signal input
flabel metal3 s 11200 1368 12000 1488 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 24 nsew signal input
flabel metal3 s 11200 2456 12000 2576 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 25 nsew signal input
flabel metal3 s 11200 3544 12000 3664 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 26 nsew signal input
flabel metal3 s 11200 4632 12000 4752 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 27 nsew signal input
flabel metal3 s 11200 5720 12000 5840 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 28 nsew signal input
flabel metal3 s 11200 6808 12000 6928 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 29 nsew signal input
flabel metal3 s 11200 7896 12000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 30 nsew signal input
flabel metal3 s 11200 8984 12000 9104 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 31 nsew signal input
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 32 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 33 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 34 nsew signal tristate
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 35 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 36 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 37 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 38 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 39 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 40 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 41 nsew signal input
flabel metal2 s 9954 11200 10010 12000 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 42 nsew signal tristate
flabel metal2 s 10966 11200 11022 12000 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 43 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 44 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 45 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 2254 5644 2254 5644 0 _000_
rlabel metal1 3128 5882 3128 5882 0 _001_
rlabel metal1 2116 4250 2116 4250 0 _002_
rlabel metal1 2116 2618 2116 2618 0 _003_
rlabel metal1 3312 3978 3312 3978 0 _004_
rlabel metal1 6578 2550 6578 2550 0 _005_
rlabel metal1 3082 5814 3082 5814 0 _006_
rlabel metal1 6210 2618 6210 2618 0 _007_
rlabel metal1 9476 6426 9476 6426 0 _008_
rlabel metal1 7084 6290 7084 6290 0 _009_
rlabel metal1 10442 7412 10442 7412 0 _010_
rlabel metal1 9154 8976 9154 8976 0 _011_
rlabel metal1 5520 4794 5520 4794 0 _012_
rlabel metal1 8648 6970 8648 6970 0 _013_
rlabel metal1 9292 4726 9292 4726 0 _014_
rlabel metal1 10258 4590 10258 4590 0 _015_
rlabel metal1 9154 3162 9154 3162 0 _016_
rlabel metal1 3450 3570 3450 3570 0 _017_
rlabel metal1 9154 7956 9154 7956 0 _018_
rlabel metal1 5934 6834 5934 6834 0 _019_
rlabel metal2 10258 7684 10258 7684 0 _020_
rlabel metal1 8510 6188 8510 6188 0 _021_
rlabel metal1 8556 8398 8556 8398 0 _022_
rlabel metal1 9430 6766 9430 6766 0 _023_
rlabel metal1 5612 6766 5612 6766 0 _024_
rlabel metal2 7774 6052 7774 6052 0 _025_
rlabel metal1 7912 8602 7912 8602 0 _026_
rlabel metal1 7636 6834 7636 6834 0 _027_
rlabel metal1 8648 6834 8648 6834 0 _028_
rlabel metal2 10074 7140 10074 7140 0 _029_
rlabel metal1 6440 3434 6440 3434 0 _030_
rlabel metal1 6026 4692 6026 4692 0 _031_
rlabel metal1 4784 2482 4784 2482 0 _032_
rlabel metal1 5704 5134 5704 5134 0 _033_
rlabel metal1 3128 2482 3128 2482 0 _034_
rlabel viali 3174 4587 3174 4587 0 _035_
rlabel metal1 4554 3400 4554 3400 0 _036_
rlabel metal1 7084 4794 7084 4794 0 _037_
rlabel metal1 4186 3706 4186 3706 0 _038_
rlabel metal1 4968 4114 4968 4114 0 _039_
rlabel metal1 2852 3570 2852 3570 0 _040_
rlabel metal1 2898 4046 2898 4046 0 _041_
rlabel metal1 4278 6732 4278 6732 0 _042_
rlabel metal2 2070 5406 2070 5406 0 _043_
rlabel metal1 3772 5882 3772 5882 0 _044_
rlabel metal1 2392 5202 2392 5202 0 _045_
rlabel via2 9982 3451 9982 3451 0 _046_
rlabel metal1 8786 3094 8786 3094 0 _047_
rlabel metal1 9292 3434 9292 3434 0 _048_
rlabel metal1 7498 2618 7498 2618 0 _049_
rlabel metal2 9982 4964 9982 4964 0 _050_
rlabel metal1 8510 4998 8510 4998 0 _051_
rlabel metal1 9982 5746 9982 5746 0 _052_
rlabel metal1 7912 5338 7912 5338 0 _053_
rlabel metal2 8694 1520 8694 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal2 9614 1571 9614 1571 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal2 10534 1639 10534 1639 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal1 10442 6800 10442 6800 0 ccff_head
rlabel metal1 9798 9146 9798 9146 0 ccff_tail
rlabel metal3 751 2516 751 2516 0 chanx_left_in[0]
rlabel metal3 843 3604 843 3604 0 chanx_left_in[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_in[2]
rlabel metal3 820 5780 820 5780 0 chanx_left_in[3]
rlabel metal3 1050 6868 1050 6868 0 chanx_left_in[4]
rlabel metal3 751 7956 751 7956 0 chanx_left_in[5]
rlabel metal3 820 9044 820 9044 0 chanx_left_in[6]
rlabel metal2 2990 9537 2990 9537 0 chanx_left_in[7]
rlabel metal3 1027 11220 1027 11220 0 chanx_left_in[8]
rlabel metal1 1288 9418 1288 9418 0 chanx_left_out[0]
rlabel metal1 2162 9622 2162 9622 0 chanx_left_out[1]
rlabel metal1 3174 9622 3174 9622 0 chanx_left_out[2]
rlabel metal1 4048 9690 4048 9690 0 chanx_left_out[3]
rlabel metal1 5198 9622 5198 9622 0 chanx_left_out[4]
rlabel metal1 6532 9622 6532 9622 0 chanx_left_out[5]
rlabel metal1 7222 9622 7222 9622 0 chanx_left_out[6]
rlabel metal1 8096 9690 8096 9690 0 chanx_left_out[7]
rlabel metal1 9246 9622 9246 9622 0 chanx_left_out[8]
rlabel metal3 2139 7276 2139 7276 0 chanx_right_in[0]
rlabel metal1 10350 2414 10350 2414 0 chanx_right_in[1]
rlabel metal1 2116 3502 2116 3502 0 chanx_right_in[2]
rlabel metal1 3726 4046 3726 4046 0 chanx_right_in[3]
rlabel metal1 10442 4114 10442 4114 0 chanx_right_in[4]
rlabel metal1 9614 6324 9614 6324 0 chanx_right_in[5]
rlabel metal1 10442 5202 10442 5202 0 chanx_right_in[6]
rlabel metal1 10810 6290 10810 6290 0 chanx_right_in[7]
rlabel metal1 6026 9486 6026 9486 0 chanx_right_in[8]
rlabel metal1 1012 2822 1012 2822 0 chanx_right_out[0]
rlabel metal1 1748 2890 1748 2890 0 chanx_right_out[1]
rlabel metal2 2254 1520 2254 1520 0 chanx_right_out[2]
rlabel metal2 3174 1571 3174 1571 0 chanx_right_out[3]
rlabel metal2 4094 959 4094 959 0 chanx_right_out[4]
rlabel metal2 5014 1520 5014 1520 0 chanx_right_out[5]
rlabel metal2 5934 823 5934 823 0 chanx_right_out[6]
rlabel metal2 6854 1571 6854 1571 0 chanx_right_out[7]
rlabel metal2 7774 1520 7774 1520 0 chanx_right_out[8]
rlabel metal1 2691 3094 2691 3094 0 clknet_0_prog_clk
rlabel metal1 2208 6290 2208 6290 0 clknet_1_0__leaf_prog_clk
rlabel metal1 6118 7990 6118 7990 0 clknet_1_1__leaf_prog_clk
rlabel metal1 7728 5678 7728 5678 0 mem_bottom_ipin_0.DFF_0_.Q
rlabel metal1 8924 6766 8924 6766 0 mem_bottom_ipin_0.DFF_1_.Q
rlabel metal1 8464 7174 8464 7174 0 mem_bottom_ipin_0.DFF_2_.Q
rlabel metal2 2622 7140 2622 7140 0 mem_bottom_ipin_1.DFF_0_.Q
rlabel metal1 3726 5746 3726 5746 0 mem_bottom_ipin_1.DFF_1_.Q
rlabel metal1 3634 4148 3634 4148 0 mem_top_ipin_0.DFF_0_.Q
rlabel metal1 3818 3536 3818 3536 0 mem_top_ipin_0.DFF_1_.Q
rlabel metal1 6026 3094 6026 3094 0 mem_top_ipin_0.DFF_2_.Q
rlabel metal1 7636 2414 7636 2414 0 mem_top_ipin_1.DFF_0_.Q
rlabel metal1 8280 3706 8280 3706 0 mem_top_ipin_1.DFF_1_.Q
rlabel metal1 8464 4590 8464 4590 0 mem_top_ipin_2.DFF_0_.Q
rlabel metal1 3542 6392 3542 6392 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 5934 6732 5934 6732 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 7636 5746 7636 5746 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 8786 5746 8786 5746 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 7498 8602 7498 8602 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal2 8050 8636 8050 8636 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 6210 6630 6210 6630 0 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 8464 6086 8464 6086 0 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 8694 8704 8694 8704 0 mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 8832 6902 8832 6902 0 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 9430 8160 9430 8160 0 mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 10120 7718 10120 7718 0 mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 2070 4658 2070 4658 0 mux_bottom_ipin_1.INVTX1_0_.out
rlabel metal1 2668 4658 2668 4658 0 mux_bottom_ipin_1.INVTX1_1_.out
rlabel metal1 3680 5338 3680 5338 0 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4554 6630 4554 6630 0 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2622 3570 2622 3570 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 2254 6120 2254 6120 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal1 3174 5576 3174 5576 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal1 5888 5202 5888 5202 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal1 3128 4726 3128 4726 0 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4370 2550 4370 2550 0 mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 5842 4998 5842 4998 0 mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 5060 2618 5060 2618 0 mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 6532 4590 6532 4590 0 mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 6762 3672 6762 3672 0 mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 6670 4114 6670 4114 0 mux_top_ipin_1.INVTX1_0_.out
rlabel metal1 8648 3026 8648 3026 0 mux_top_ipin_1.INVTX1_1_.out
rlabel via1 8878 3570 8878 3570 0 mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9706 3400 9706 3400 0 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9016 5814 9016 5814 0 mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 10304 5338 10304 5338 0 mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 10350 6630 10350 6630 0 net1
rlabel metal2 2714 8976 2714 8976 0 net10
rlabel metal1 2254 8058 2254 8058 0 net11
rlabel metal1 10212 2278 10212 2278 0 net12
rlabel metal1 1610 6290 1610 6290 0 net13
rlabel metal1 3818 3910 3818 3910 0 net14
rlabel metal1 7406 5644 7406 5644 0 net15
rlabel metal1 9108 6086 9108 6086 0 net16
rlabel metal1 6578 6290 6578 6290 0 net17
rlabel metal1 10258 6426 10258 6426 0 net18
rlabel metal1 9246 9010 9246 9010 0 net19
rlabel metal1 1932 4794 1932 4794 0 net2
rlabel metal1 8786 2346 8786 2346 0 net20
rlabel metal1 9729 2346 9729 2346 0 net21
rlabel metal1 10166 3094 10166 3094 0 net22
rlabel metal1 10166 6290 10166 6290 0 net23
rlabel metal1 1656 9146 1656 9146 0 net24
rlabel metal1 2024 3978 2024 3978 0 net25
rlabel metal1 2944 7514 2944 7514 0 net26
rlabel metal1 4186 9146 4186 9146 0 net27
rlabel metal1 5198 9146 5198 9146 0 net28
rlabel metal1 6486 9520 6486 9520 0 net29
rlabel metal1 1840 5338 1840 5338 0 net3
rlabel metal1 7268 7514 7268 7514 0 net30
rlabel metal1 9476 8602 9476 8602 0 net31
rlabel metal1 9384 9554 9384 9554 0 net32
rlabel metal1 1656 3094 1656 3094 0 net33
rlabel metal2 2714 5236 2714 5236 0 net34
rlabel metal1 1702 2346 1702 2346 0 net35
rlabel metal1 2300 2414 2300 2414 0 net36
rlabel metal2 3956 2550 3956 2550 0 net37
rlabel metal3 2599 7276 2599 7276 0 net38
rlabel metal1 5888 2346 5888 2346 0 net39
rlabel metal1 1656 5338 1656 5338 0 net4
rlabel metal1 7360 2482 7360 2482 0 net40
rlabel metal1 8142 2414 8142 2414 0 net41
rlabel metal1 10212 8602 10212 8602 0 net42
rlabel metal1 6302 7446 6302 7446 0 net43
rlabel metal1 9016 7922 9016 7922 0 net44
rlabel metal1 5842 4726 5842 4726 0 net45
rlabel metal2 4094 7072 4094 7072 0 net46
rlabel metal2 9890 3808 9890 3808 0 net47
rlabel metal1 9522 5202 9522 5202 0 net48
rlabel metal1 6757 3094 6757 3094 0 net49
rlabel metal1 1610 6188 1610 6188 0 net5
rlabel metal1 4411 5270 4411 5270 0 net50
rlabel metal1 9292 4794 9292 4794 0 net51
rlabel viali 2510 6289 2510 6289 0 net52
rlabel metal2 8694 4386 8694 4386 0 net53
rlabel metal1 8188 3162 8188 3162 0 net54
rlabel metal1 2272 6766 2272 6766 0 net55
rlabel metal1 4733 4590 4733 4590 0 net56
rlabel metal1 8091 7446 8091 7446 0 net57
rlabel metal1 5147 3094 5147 3094 0 net58
rlabel metal1 6665 7854 6665 7854 0 net59
rlabel metal1 2185 7242 2185 7242 0 net6
rlabel metal1 1978 7412 1978 7412 0 net7
rlabel metal2 2438 5780 2438 5780 0 net8
rlabel metal1 6302 9010 6302 9010 0 net9
rlabel metal3 2384 1428 2384 1428 0 prog_clk
rlabel metal1 10258 9622 10258 9622 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal1 10488 9078 10488 9078 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
