magic
tech sky130A
magscale 1 2
timestamp 1708041115
<< obsli1 >>
rect 1104 2159 12880 11441
<< obsm1 >>
rect 750 2128 13040 11620
<< metal2 >>
rect 938 13200 994 14000
rect 2134 13200 2190 14000
rect 3330 13200 3386 14000
rect 4526 13200 4582 14000
rect 5722 13200 5778 14000
rect 6918 13200 6974 14000
rect 8114 13200 8170 14000
rect 9310 13200 9366 14000
rect 10506 13200 10562 14000
rect 11702 13200 11758 14000
rect 12898 13200 12954 14000
rect 754 0 810 800
rect 2134 0 2190 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 6274 0 6330 800
rect 7654 0 7710 800
rect 9034 0 9090 800
rect 10414 0 10470 800
rect 11794 0 11850 800
<< obsm2 >>
rect 756 13144 882 13433
rect 1050 13144 2078 13433
rect 2246 13144 3274 13433
rect 3442 13144 4470 13433
rect 4638 13144 5666 13433
rect 5834 13144 6862 13433
rect 7030 13144 8058 13433
rect 8226 13144 9254 13433
rect 9422 13144 10450 13433
rect 10618 13144 11646 13433
rect 11814 13144 12842 13433
rect 13010 13144 13034 13433
rect 756 856 13034 13144
rect 866 303 2078 856
rect 2246 303 3458 856
rect 3626 303 4838 856
rect 5006 303 6218 856
rect 6386 303 7598 856
rect 7766 303 8978 856
rect 9146 303 10358 856
rect 10526 303 11738 856
rect 11906 303 13034 856
<< metal3 >>
rect 13200 13336 14000 13456
rect 0 12248 800 12368
rect 13200 12248 14000 12368
rect 0 11160 800 11280
rect 13200 11160 14000 11280
rect 0 10072 800 10192
rect 13200 10072 14000 10192
rect 0 8984 800 9104
rect 13200 8984 14000 9104
rect 0 7896 800 8016
rect 13200 7896 14000 8016
rect 0 6808 800 6928
rect 13200 6808 14000 6928
rect 0 5720 800 5840
rect 13200 5720 14000 5840
rect 0 4632 800 4752
rect 13200 4632 14000 4752
rect 0 3544 800 3664
rect 13200 3544 14000 3664
rect 0 2456 800 2576
rect 13200 2456 14000 2576
rect 13200 1368 14000 1488
rect 13200 280 14000 400
<< obsm3 >>
rect 798 13256 13120 13429
rect 798 12448 13200 13256
rect 880 12168 13120 12448
rect 798 11360 13200 12168
rect 880 11080 13120 11360
rect 798 10272 13200 11080
rect 880 9992 13120 10272
rect 798 9184 13200 9992
rect 880 8904 13120 9184
rect 798 8096 13200 8904
rect 880 7816 13120 8096
rect 798 7008 13200 7816
rect 880 6728 13120 7008
rect 798 5920 13200 6728
rect 880 5640 13120 5920
rect 798 4832 13200 5640
rect 880 4552 13120 4832
rect 798 3744 13200 4552
rect 880 3464 13120 3744
rect 798 2656 13200 3464
rect 880 2376 13120 2656
rect 798 1568 13200 2376
rect 798 1288 13120 1568
rect 798 480 13200 1288
rect 798 307 13120 480
<< metal4 >>
rect 2416 2128 2736 11472
rect 3888 2128 4208 11472
rect 5360 2128 5680 11472
rect 6832 2128 7152 11472
rect 8304 2128 8624 11472
rect 9776 2128 10096 11472
rect 11248 2128 11568 11472
rect 12720 2128 13040 11472
<< labels >>
rlabel metal3 s 13200 11160 14000 11280 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 13200 12248 14000 12368 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 chanx_right_in[0]
port 3 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 chanx_right_in[1]
port 4 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_right_in[2]
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_right_in[3]
port 6 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 chanx_right_in[4]
port 7 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_right_in[5]
port 8 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_right_in[6]
port 9 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_right_in[7]
port 10 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_right_in[8]
port 11 nsew signal input
rlabel metal2 s 754 0 810 800 6 chanx_right_out[0]
port 12 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 chanx_right_out[1]
port 13 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 chanx_right_out[2]
port 14 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 chanx_right_out[3]
port 15 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 chanx_right_out[4]
port 16 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 chanx_right_out[5]
port 17 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 chanx_right_out[6]
port 18 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 chanx_right_out[7]
port 19 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 chanx_right_out[8]
port 20 nsew signal output
rlabel metal2 s 2134 13200 2190 14000 6 chany_top_in[0]
port 21 nsew signal input
rlabel metal2 s 3330 13200 3386 14000 6 chany_top_in[1]
port 22 nsew signal input
rlabel metal2 s 4526 13200 4582 14000 6 chany_top_in[2]
port 23 nsew signal input
rlabel metal2 s 5722 13200 5778 14000 6 chany_top_in[3]
port 24 nsew signal input
rlabel metal2 s 6918 13200 6974 14000 6 chany_top_in[4]
port 25 nsew signal input
rlabel metal2 s 8114 13200 8170 14000 6 chany_top_in[5]
port 26 nsew signal input
rlabel metal2 s 9310 13200 9366 14000 6 chany_top_in[6]
port 27 nsew signal input
rlabel metal2 s 10506 13200 10562 14000 6 chany_top_in[7]
port 28 nsew signal input
rlabel metal2 s 11702 13200 11758 14000 6 chany_top_in[8]
port 29 nsew signal input
rlabel metal3 s 13200 1368 14000 1488 6 chany_top_out[0]
port 30 nsew signal output
rlabel metal3 s 13200 2456 14000 2576 6 chany_top_out[1]
port 31 nsew signal output
rlabel metal3 s 13200 3544 14000 3664 6 chany_top_out[2]
port 32 nsew signal output
rlabel metal3 s 13200 4632 14000 4752 6 chany_top_out[3]
port 33 nsew signal output
rlabel metal3 s 13200 5720 14000 5840 6 chany_top_out[4]
port 34 nsew signal output
rlabel metal3 s 13200 6808 14000 6928 6 chany_top_out[5]
port 35 nsew signal output
rlabel metal3 s 13200 7896 14000 8016 6 chany_top_out[6]
port 36 nsew signal output
rlabel metal3 s 13200 8984 14000 9104 6 chany_top_out[7]
port 37 nsew signal output
rlabel metal3 s 13200 10072 14000 10192 6 chany_top_out[8]
port 38 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 prog_clk
port 39 nsew signal input
rlabel metal3 s 13200 13336 14000 13456 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 40 nsew signal input
rlabel metal3 s 13200 280 14000 400 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_
port 41 nsew signal input
rlabel metal2 s 12898 13200 12954 14000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 42 nsew signal input
rlabel metal2 s 938 13200 994 14000 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 43 nsew signal input
rlabel metal4 s 2416 2128 2736 11472 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 5360 2128 5680 11472 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 8304 2128 8624 11472 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 11248 2128 11568 11472 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 3888 2128 4208 11472 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 6832 2128 7152 11472 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 9776 2128 10096 11472 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 12720 2128 13040 11472 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 14000 14000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 360690
string GDS_FILE /home/baungarten2/Desktop/Caravel_FPGA/openlane/sb_0__0_/runs/24_02_15_17_51/results/signoff/sb_0__0_.magic.gds
string GDS_START 89992
<< end >>

